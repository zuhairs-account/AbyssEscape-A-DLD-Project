module distortBG_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		14'b00000001000001: color_data = 12'b001000000000;
		14'b00000001011001: color_data = 12'b001000000000;
		14'b00000001011010: color_data = 12'b010000000000;
		14'b00000001011011: color_data = 12'b010000000000;
		14'b00000001011100: color_data = 12'b010000000000;
		14'b00000001011101: color_data = 12'b010000000000;
		14'b00000001011110: color_data = 12'b010000000000;
		14'b00000001011111: color_data = 12'b010000000000;
		14'b00000001100000: color_data = 12'b010000000000;
		14'b00000001100001: color_data = 12'b010000000000;
		14'b00000001100010: color_data = 12'b010000000000;
		14'b00000001100011: color_data = 12'b010000000000;
		14'b00000001100100: color_data = 12'b010000000000;
		14'b00000001100101: color_data = 12'b010000000000;
		14'b00000001100110: color_data = 12'b010000000000;
		14'b00000001100111: color_data = 12'b001000000000;
		14'b00000011000101: color_data = 12'b001000000000;
		14'b00000011000110: color_data = 12'b001000000000;
		14'b00000011000111: color_data = 12'b001000000000;
		14'b00000011001000: color_data = 12'b001000000000;
		14'b00000011001001: color_data = 12'b001000000000;
		14'b00000011001011: color_data = 12'b001000000000;
		14'b00000011011010: color_data = 12'b001000000000;
		14'b00000011011011: color_data = 12'b010000000000;
		14'b00000011011100: color_data = 12'b010000000000;
		14'b00000011011101: color_data = 12'b010000000000;
		14'b00000011011110: color_data = 12'b010000000000;
		14'b00000011011111: color_data = 12'b010000000000;
		14'b00000011100000: color_data = 12'b010000000000;
		14'b00000011100001: color_data = 12'b010000000000;
		14'b00000011100010: color_data = 12'b010000000000;
		14'b00000011100011: color_data = 12'b010000000000;
		14'b00000011100100: color_data = 12'b010000000000;
		14'b00000011100101: color_data = 12'b010000000000;
		14'b00000011100110: color_data = 12'b010000000000;
		14'b00000011100111: color_data = 12'b010000000000;
		14'b00000011101000: color_data = 12'b001000000000;
		14'b00000100010101: color_data = 12'b001000000000;
		14'b00000100011100: color_data = 12'b001000000000;
		14'b00000100011101: color_data = 12'b001000000000;
		14'b00000100011110: color_data = 12'b001000000000;
		14'b00000100011111: color_data = 12'b001000000000;
		14'b00000100100000: color_data = 12'b001000000000;
		14'b00000101000110: color_data = 12'b001000000000;
		14'b00000101000111: color_data = 12'b001000000000;
		14'b00000101001000: color_data = 12'b001000000000;
		14'b00000101001001: color_data = 12'b001000000000;
		14'b00000101001010: color_data = 12'b001000000000;
		14'b00000101001011: color_data = 12'b001000000000;
		14'b00000101001100: color_data = 12'b001000000000;
		14'b00000101001101: color_data = 12'b001000000000;
		14'b00000101011011: color_data = 12'b001000000000;
		14'b00000101011100: color_data = 12'b001000000000;
		14'b00000101011101: color_data = 12'b010000000000;
		14'b00000101011110: color_data = 12'b010000000000;
		14'b00000101011111: color_data = 12'b010000000000;
		14'b00000101100000: color_data = 12'b010000000000;
		14'b00000101100001: color_data = 12'b010000000000;
		14'b00000101100010: color_data = 12'b010000000000;
		14'b00000101100011: color_data = 12'b010000000000;
		14'b00000101100100: color_data = 12'b010000000000;
		14'b00000101100101: color_data = 12'b010000000000;
		14'b00000101100110: color_data = 12'b010000000000;
		14'b00000101100111: color_data = 12'b001000000000;
		14'b00000101101000: color_data = 12'b001000000000;
		14'b00000110000011: color_data = 12'b001000000000;
		14'b00000110000100: color_data = 12'b001000000000;
		14'b00000110000101: color_data = 12'b001000000000;
		14'b00000110000110: color_data = 12'b001000000000;
		14'b00000110000111: color_data = 12'b001000000000;
		14'b00000110001000: color_data = 12'b001000000000;
		14'b00000110001001: color_data = 12'b001000000000;
		14'b00000110001010: color_data = 12'b001000000000;
		14'b00000110001011: color_data = 12'b001000000000;
		14'b00000110001101: color_data = 12'b001000000000;
		14'b00000110001110: color_data = 12'b001000000000;
		14'b00000110010011: color_data = 12'b001000000000;
		14'b00000110010101: color_data = 12'b010000000000;
		14'b00000110011100: color_data = 12'b001000000000;
		14'b00000110011101: color_data = 12'b001000000000;
		14'b00000110011110: color_data = 12'b001000000000;
		14'b00000110011111: color_data = 12'b001000000000;
		14'b00000110100000: color_data = 12'b001000000000;
		14'b00000110100001: color_data = 12'b001000000000;
		14'b00000110100010: color_data = 12'b001000000000;
		14'b00000111001101: color_data = 12'b001000000000;
		14'b00000111011101: color_data = 12'b001000000000;
		14'b00000111011110: color_data = 12'b010000000000;
		14'b00000111011111: color_data = 12'b010000000000;
		14'b00000111100000: color_data = 12'b010000000000;
		14'b00000111100001: color_data = 12'b010000000000;
		14'b00000111100010: color_data = 12'b010000000000;
		14'b00000111100011: color_data = 12'b010000000000;
		14'b00000111100100: color_data = 12'b010000000000;
		14'b00000111100101: color_data = 12'b010000000000;
		14'b00000111100110: color_data = 12'b010000000000;
		14'b00000111100111: color_data = 12'b001000000000;
		14'b00000111110000: color_data = 12'b001000000000;
		14'b00001000001001: color_data = 12'b001000000000;
		14'b00001000001010: color_data = 12'b001000000000;
		14'b00001000001011: color_data = 12'b001000000000;
		14'b00001000001101: color_data = 12'b001000000000;
		14'b00001000001110: color_data = 12'b001000000000;
		14'b00001000001111: color_data = 12'b010000000000;
		14'b00001000010000: color_data = 12'b010000000000;
		14'b00001000010011: color_data = 12'b001000000000;
		14'b00001000010100: color_data = 12'b010000000000;
		14'b00001000010101: color_data = 12'b010000000000;
		14'b00001000010110: color_data = 12'b010000000000;
		14'b00001000010111: color_data = 12'b010000000000;
		14'b00001000011000: color_data = 12'b010000000000;
		14'b00001000011001: color_data = 12'b010000000000;
		14'b00001000011010: color_data = 12'b010000000000;
		14'b00001000011011: color_data = 12'b010000000000;
		14'b00001000011100: color_data = 12'b010000000000;
		14'b00001000011101: color_data = 12'b001000000000;
		14'b00001000011110: color_data = 12'b001000000000;
		14'b00001000011111: color_data = 12'b001000000000;
		14'b00001000100000: color_data = 12'b001000000000;
		14'b00001000100001: color_data = 12'b001000000000;
		14'b00001000100010: color_data = 12'b001000000000;
		14'b00001001011101: color_data = 12'b001000000000;
		14'b00001001011110: color_data = 12'b010000000000;
		14'b00001001011111: color_data = 12'b010000000000;
		14'b00001001100000: color_data = 12'b010000000000;
		14'b00001001100001: color_data = 12'b010000000000;
		14'b00001001100010: color_data = 12'b010000000000;
		14'b00001001100011: color_data = 12'b010000000000;
		14'b00001001100100: color_data = 12'b010000000000;
		14'b00001001100101: color_data = 12'b010000000000;
		14'b00001001100110: color_data = 12'b001000000000;
		14'b00001001101110: color_data = 12'b010000000000;
		14'b00001001101111: color_data = 12'b010000000000;
		14'b00001010001010: color_data = 12'b001000000000;
		14'b00001010001011: color_data = 12'b001000000000;
		14'b00001010001100: color_data = 12'b001000000000;
		14'b00001010001101: color_data = 12'b010000000000;
		14'b00001010001110: color_data = 12'b010000000000;
		14'b00001010001111: color_data = 12'b010000000000;
		14'b00001010010000: color_data = 12'b010000000000;
		14'b00001010010001: color_data = 12'b001000000000;
		14'b00001010010010: color_data = 12'b001000000000;
		14'b00001010010011: color_data = 12'b001000000000;
		14'b00001010010100: color_data = 12'b010000000000;
		14'b00001010010101: color_data = 12'b010000000000;
		14'b00001010010110: color_data = 12'b010000000000;
		14'b00001010010111: color_data = 12'b010000000000;
		14'b00001010011000: color_data = 12'b010000000000;
		14'b00001010011001: color_data = 12'b010000000000;
		14'b00001010011010: color_data = 12'b010000000000;
		14'b00001010011011: color_data = 12'b010000000000;
		14'b00001010011100: color_data = 12'b010000000000;
		14'b00001010011101: color_data = 12'b010000000000;
		14'b00001010011110: color_data = 12'b010000000000;
		14'b00001010011111: color_data = 12'b010000000000;
		14'b00001010100000: color_data = 12'b001000000000;
		14'b00001010100001: color_data = 12'b001000000000;
		14'b00001010100010: color_data = 12'b001000000000;
		14'b00001010100011: color_data = 12'b001000000000;
		14'b00001011011100: color_data = 12'b001000000000;
		14'b00001011011101: color_data = 12'b010000000000;
		14'b00001011011110: color_data = 12'b010000000000;
		14'b00001011011111: color_data = 12'b010000000000;
		14'b00001011100000: color_data = 12'b010000000000;
		14'b00001011100001: color_data = 12'b010000000000;
		14'b00001011100010: color_data = 12'b010000000000;
		14'b00001011100011: color_data = 12'b010000000000;
		14'b00001011100100: color_data = 12'b010000000000;
		14'b00001011100101: color_data = 12'b010000000000;
		14'b00001011100110: color_data = 12'b001000000000;
		14'b00001011101100: color_data = 12'b001000000000;
		14'b00001011101101: color_data = 12'b010000000000;
		14'b00001011101110: color_data = 12'b010000000000;
		14'b00001011101111: color_data = 12'b001000000000;
		14'b00001100001010: color_data = 12'b001000000000;
		14'b00001100001011: color_data = 12'b001000000000;
		14'b00001100001100: color_data = 12'b010000000000;
		14'b00001100001101: color_data = 12'b010000000000;
		14'b00001100001110: color_data = 12'b010000000000;
		14'b00001100001111: color_data = 12'b010000000000;
		14'b00001100010000: color_data = 12'b010000000000;
		14'b00001100010001: color_data = 12'b010000000000;
		14'b00001100010010: color_data = 12'b010000000000;
		14'b00001100010011: color_data = 12'b010000000000;
		14'b00001100010100: color_data = 12'b010000000000;
		14'b00001100010101: color_data = 12'b010000000000;
		14'b00001100010110: color_data = 12'b010000000000;
		14'b00001100010111: color_data = 12'b010000000000;
		14'b00001100011000: color_data = 12'b010000000000;
		14'b00001100011001: color_data = 12'b010000000000;
		14'b00001100011010: color_data = 12'b010000000000;
		14'b00001100011011: color_data = 12'b010000000000;
		14'b00001100011100: color_data = 12'b010000000000;
		14'b00001100011101: color_data = 12'b010000000000;
		14'b00001100011110: color_data = 12'b010000000000;
		14'b00001100011111: color_data = 12'b010000000000;
		14'b00001100100000: color_data = 12'b010000000000;
		14'b00001100100001: color_data = 12'b010000000000;
		14'b00001100100010: color_data = 12'b010000000000;
		14'b00001100100011: color_data = 12'b010000000000;
		14'b00001100100100: color_data = 12'b010000000000;
		14'b00001100100101: color_data = 12'b001000000000;
		14'b00001101011011: color_data = 12'b010000000000;
		14'b00001101011100: color_data = 12'b010000000000;
		14'b00001101011101: color_data = 12'b010000000000;
		14'b00001101011110: color_data = 12'b010000000000;
		14'b00001101011111: color_data = 12'b010000000000;
		14'b00001101100000: color_data = 12'b010000000000;
		14'b00001101100001: color_data = 12'b010000000000;
		14'b00001101100010: color_data = 12'b010000000000;
		14'b00001101100011: color_data = 12'b010000000000;
		14'b00001101100100: color_data = 12'b010000000000;
		14'b00001101100101: color_data = 12'b001000000000;
		14'b00001101101011: color_data = 12'b010000000000;
		14'b00001101101100: color_data = 12'b010000000000;
		14'b00001101101101: color_data = 12'b010000000000;
		14'b00001110001000: color_data = 12'b001000000000;
		14'b00001110001001: color_data = 12'b010000000000;
		14'b00001110001010: color_data = 12'b010000000000;
		14'b00001110001011: color_data = 12'b010000000000;
		14'b00001110001100: color_data = 12'b010000000000;
		14'b00001110001101: color_data = 12'b010000000000;
		14'b00001110001110: color_data = 12'b010000000000;
		14'b00001110001111: color_data = 12'b010000000000;
		14'b00001110010000: color_data = 12'b010000000000;
		14'b00001110010001: color_data = 12'b010000000000;
		14'b00001110010010: color_data = 12'b010000000000;
		14'b00001110010011: color_data = 12'b010000000000;
		14'b00001110010100: color_data = 12'b010000000000;
		14'b00001110010101: color_data = 12'b010000000000;
		14'b00001110010110: color_data = 12'b010000000000;
		14'b00001110010111: color_data = 12'b010000000000;
		14'b00001110011000: color_data = 12'b010000000000;
		14'b00001110011001: color_data = 12'b010000000000;
		14'b00001110011010: color_data = 12'b010000000000;
		14'b00001110011011: color_data = 12'b010000000000;
		14'b00001110011100: color_data = 12'b010000000000;
		14'b00001110011101: color_data = 12'b001000000000;
		14'b00001110011110: color_data = 12'b001000000000;
		14'b00001110011111: color_data = 12'b010000000000;
		14'b00001110100000: color_data = 12'b010000000000;
		14'b00001110100001: color_data = 12'b010000000000;
		14'b00001110100010: color_data = 12'b010000000000;
		14'b00001110100011: color_data = 12'b010000000000;
		14'b00001110100100: color_data = 12'b010000000000;
		14'b00001110100101: color_data = 12'b010000000000;
		14'b00001110100110: color_data = 12'b010000000000;
		14'b00001111011010: color_data = 12'b001000000000;
		14'b00001111011011: color_data = 12'b010000000000;
		14'b00001111011100: color_data = 12'b010000000000;
		14'b00001111011101: color_data = 12'b010000000000;
		14'b00001111011110: color_data = 12'b010000000000;
		14'b00001111011111: color_data = 12'b010000000000;
		14'b00001111100000: color_data = 12'b010000000000;
		14'b00001111100001: color_data = 12'b010000000000;
		14'b00001111100010: color_data = 12'b010000000000;
		14'b00001111100011: color_data = 12'b010000000000;
		14'b00001111100100: color_data = 12'b010000000000;
		14'b00001111100101: color_data = 12'b001000000000;
		14'b00001111101010: color_data = 12'b010000000000;
		14'b00001111101011: color_data = 12'b010000000000;
		14'b00001111101100: color_data = 12'b010000000000;
		14'b00010000000111: color_data = 12'b001000000000;
		14'b00010000001000: color_data = 12'b010000000000;
		14'b00010000001001: color_data = 12'b010000000000;
		14'b00010000001010: color_data = 12'b010000000000;
		14'b00010000001011: color_data = 12'b010000000000;
		14'b00010000001100: color_data = 12'b010000000000;
		14'b00010000001101: color_data = 12'b010000000000;
		14'b00010000001110: color_data = 12'b010000000000;
		14'b00010000001111: color_data = 12'b010000000000;
		14'b00010000010000: color_data = 12'b010000000000;
		14'b00010000010001: color_data = 12'b010000000000;
		14'b00010000010010: color_data = 12'b010000000000;
		14'b00010000010011: color_data = 12'b010000000000;
		14'b00010000010100: color_data = 12'b010000000000;
		14'b00010000010101: color_data = 12'b010000000000;
		14'b00010000010110: color_data = 12'b010000000000;
		14'b00010000010111: color_data = 12'b010000000000;
		14'b00010000011000: color_data = 12'b010000000000;
		14'b00010000011001: color_data = 12'b010000000000;
		14'b00010000011010: color_data = 12'b010000000000;
		14'b00010000011011: color_data = 12'b010000000000;
		14'b00010000011100: color_data = 12'b010000000000;
		14'b00010000011101: color_data = 12'b001000000000;
		14'b00010000011110: color_data = 12'b001000000000;
		14'b00010000100000: color_data = 12'b001000000000;
		14'b00010000100001: color_data = 12'b010000000000;
		14'b00010000100010: color_data = 12'b010000000000;
		14'b00010000100011: color_data = 12'b010000000000;
		14'b00010000100100: color_data = 12'b010000000000;
		14'b00010000100101: color_data = 12'b010000000000;
		14'b00010000100110: color_data = 12'b010000000000;
		14'b00010000100111: color_data = 12'b010000000000;
		14'b00010000101000: color_data = 12'b010000000000;
		14'b00010001011010: color_data = 12'b001000000000;
		14'b00010001011011: color_data = 12'b010000000000;
		14'b00010001011100: color_data = 12'b010000000000;
		14'b00010001011101: color_data = 12'b010000000000;
		14'b00010001011110: color_data = 12'b010000000000;
		14'b00010001011111: color_data = 12'b010000000000;
		14'b00010001100000: color_data = 12'b010000000000;
		14'b00010001100001: color_data = 12'b010000000000;
		14'b00010001100010: color_data = 12'b010000000000;
		14'b00010001100011: color_data = 12'b010000000000;
		14'b00010001100100: color_data = 12'b010000000000;
		14'b00010001100101: color_data = 12'b010000000000;
		14'b00010001100110: color_data = 12'b001000000000;
		14'b00010001101000: color_data = 12'b001000000000;
		14'b00010001101001: color_data = 12'b010000000000;
		14'b00010001101010: color_data = 12'b010000000000;
		14'b00010001101011: color_data = 12'b010000000000;
		14'b00010010000110: color_data = 12'b001000000000;
		14'b00010010000111: color_data = 12'b001000000000;
		14'b00010010001000: color_data = 12'b010000000000;
		14'b00010010001001: color_data = 12'b010000000000;
		14'b00010010001010: color_data = 12'b001000000000;
		14'b00010010001011: color_data = 12'b001000000000;
		14'b00010010001100: color_data = 12'b001000000000;
		14'b00010010001101: color_data = 12'b001000000000;
		14'b00010010001110: color_data = 12'b010000000000;
		14'b00010010001111: color_data = 12'b010000000000;
		14'b00010010010000: color_data = 12'b010000000000;
		14'b00010010010001: color_data = 12'b010000000000;
		14'b00010010010010: color_data = 12'b010000000000;
		14'b00010010010011: color_data = 12'b010000000000;
		14'b00010010011010: color_data = 12'b001000000000;
		14'b00010010011011: color_data = 12'b010000000000;
		14'b00010010011100: color_data = 12'b010000000000;
		14'b00010010011101: color_data = 12'b010000000000;
		14'b00010010011110: color_data = 12'b001000000000;
		14'b00010010100011: color_data = 12'b001000000000;
		14'b00010010100100: color_data = 12'b001000000000;
		14'b00010010100101: color_data = 12'b010000000000;
		14'b00010010100110: color_data = 12'b010000000000;
		14'b00010010100111: color_data = 12'b010000000000;
		14'b00010010101000: color_data = 12'b010000000000;
		14'b00010010101001: color_data = 12'b001000000000;
		14'b00010010101010: color_data = 12'b001000000000;
		14'b00010011011010: color_data = 12'b001000000000;
		14'b00010011011011: color_data = 12'b010000000000;
		14'b00010011011100: color_data = 12'b010000000000;
		14'b00010011011101: color_data = 12'b010000000000;
		14'b00010011011110: color_data = 12'b010000000000;
		14'b00010011011111: color_data = 12'b010000000000;
		14'b00010011100000: color_data = 12'b010000000000;
		14'b00010011100001: color_data = 12'b010000000000;
		14'b00010011100010: color_data = 12'b010000000000;
		14'b00010011100011: color_data = 12'b010000000000;
		14'b00010011100100: color_data = 12'b010000000000;
		14'b00010011100101: color_data = 12'b010000000000;
		14'b00010011100110: color_data = 12'b001000000000;
		14'b00010011100111: color_data = 12'b001000000000;
		14'b00010011101000: color_data = 12'b001000000000;
		14'b00010011101001: color_data = 12'b010000000000;
		14'b00010011101010: color_data = 12'b010000000000;
		14'b00010100000110: color_data = 12'b001000000000;
		14'b00010100000111: color_data = 12'b001000000000;
		14'b00010100001011: color_data = 12'b001000000000;
		14'b00010100001100: color_data = 12'b001000000000;
		14'b00010100001101: color_data = 12'b001000000000;
		14'b00010100001110: color_data = 12'b010000000000;
		14'b00010100001111: color_data = 12'b010000000000;
		14'b00010100010000: color_data = 12'b010000000000;
		14'b00010100010001: color_data = 12'b010000000000;
		14'b00010100011011: color_data = 12'b001000000000;
		14'b00010100011100: color_data = 12'b010000000000;
		14'b00010100011101: color_data = 12'b010000000000;
		14'b00010100011110: color_data = 12'b010000000000;
		14'b00010100011111: color_data = 12'b001000000000;
		14'b00010100100111: color_data = 12'b001000000000;
		14'b00010100101000: color_data = 12'b010000000000;
		14'b00010100101001: color_data = 12'b010000000000;
		14'b00010100101010: color_data = 12'b010000000000;
		14'b00010100101011: color_data = 12'b001000000000;
		14'b00010100101100: color_data = 12'b001000000000;
		14'b00010101011010: color_data = 12'b001000000000;
		14'b00010101011011: color_data = 12'b010000000000;
		14'b00010101011100: color_data = 12'b010000000000;
		14'b00010101011101: color_data = 12'b010000000000;
		14'b00010101011110: color_data = 12'b010000000000;
		14'b00010101011111: color_data = 12'b010000000000;
		14'b00010101100000: color_data = 12'b010000000000;
		14'b00010101100001: color_data = 12'b010000000000;
		14'b00010101100010: color_data = 12'b010000000000;
		14'b00010101100011: color_data = 12'b010000000000;
		14'b00010101100100: color_data = 12'b010000000000;
		14'b00010101100101: color_data = 12'b010000000000;
		14'b00010101100110: color_data = 12'b001000000000;
		14'b00010101100111: color_data = 12'b001000000000;
		14'b00010101101000: color_data = 12'b001000000000;
		14'b00010101101001: color_data = 12'b010000000000;
		14'b00010101101010: color_data = 12'b010000000000;
		14'b00010110000101: color_data = 12'b001000000000;
		14'b00010110000110: color_data = 12'b001000000000;
		14'b00010110001011: color_data = 12'b001000000000;
		14'b00010110001100: color_data = 12'b001000000000;
		14'b00010110001101: color_data = 12'b001000000000;
		14'b00010110001110: color_data = 12'b010000000000;
		14'b00010110001111: color_data = 12'b010000000000;
		14'b00010110010000: color_data = 12'b010000000000;
		14'b00010110011011: color_data = 12'b001000000000;
		14'b00010110011100: color_data = 12'b010000000000;
		14'b00010110011101: color_data = 12'b010000000000;
		14'b00010110011110: color_data = 12'b010000000000;
		14'b00010110011111: color_data = 12'b010000000000;
		14'b00010110100000: color_data = 12'b010000000000;
		14'b00010110100001: color_data = 12'b001000000000;
		14'b00010110100010: color_data = 12'b001000000000;
		14'b00010110101001: color_data = 12'b001000000000;
		14'b00010110101010: color_data = 12'b010000000000;
		14'b00010110101011: color_data = 12'b010000000000;
		14'b00010110101100: color_data = 12'b010000000000;
		14'b00010110101101: color_data = 12'b001000000000;
		14'b00010110101110: color_data = 12'b001000000000;
		14'b00010111010001: color_data = 12'b001000000000;
		14'b00010111010010: color_data = 12'b001000000000;
		14'b00010111011010: color_data = 12'b001000000000;
		14'b00010111011011: color_data = 12'b010000000000;
		14'b00010111011100: color_data = 12'b010000000000;
		14'b00010111011101: color_data = 12'b010000000000;
		14'b00010111011110: color_data = 12'b010000000000;
		14'b00010111011111: color_data = 12'b010000000000;
		14'b00010111100000: color_data = 12'b010000000000;
		14'b00010111100001: color_data = 12'b010000000000;
		14'b00010111100010: color_data = 12'b010000000000;
		14'b00010111100011: color_data = 12'b010000000000;
		14'b00010111100100: color_data = 12'b010000000000;
		14'b00010111100101: color_data = 12'b010000000000;
		14'b00010111100110: color_data = 12'b001000000000;
		14'b00010111100111: color_data = 12'b001000000000;
		14'b00010111101000: color_data = 12'b010000000000;
		14'b00010111101001: color_data = 12'b010000000000;
		14'b00011000000101: color_data = 12'b001000000000;
		14'b00011000000110: color_data = 12'b001000000000;
		14'b00011000001011: color_data = 12'b001000000000;
		14'b00011000001100: color_data = 12'b001000000000;
		14'b00011000001101: color_data = 12'b010000000000;
		14'b00011000001110: color_data = 12'b010000000000;
		14'b00011000001111: color_data = 12'b010000000000;
		14'b00011000010000: color_data = 12'b001000000000;
		14'b00011000010111: color_data = 12'b001000000000;
		14'b00011000011000: color_data = 12'b001000000000;
		14'b00011000011001: color_data = 12'b001000000000;
		14'b00011000011010: color_data = 12'b001000000000;
		14'b00011000011011: color_data = 12'b010000000000;
		14'b00011000011100: color_data = 12'b010000000000;
		14'b00011000011101: color_data = 12'b010000000000;
		14'b00011000011110: color_data = 12'b010000000000;
		14'b00011000011111: color_data = 12'b010000000000;
		14'b00011000100000: color_data = 12'b010000000000;
		14'b00011000100001: color_data = 12'b010000000000;
		14'b00011000100010: color_data = 12'b010000000000;
		14'b00011000100011: color_data = 12'b010000000000;
		14'b00011000100100: color_data = 12'b001000000000;
		14'b00011000100101: color_data = 12'b001000000000;
		14'b00011000101011: color_data = 12'b010000000000;
		14'b00011000101100: color_data = 12'b010000000000;
		14'b00011000101101: color_data = 12'b001000000000;
		14'b00011000101110: color_data = 12'b001000000000;
		14'b00011000101111: color_data = 12'b001000000000;
		14'b00011001011010: color_data = 12'b001000000000;
		14'b00011001011011: color_data = 12'b010000000000;
		14'b00011001011100: color_data = 12'b010000000000;
		14'b00011001011101: color_data = 12'b010000000000;
		14'b00011001011110: color_data = 12'b010000000000;
		14'b00011001011111: color_data = 12'b010000000000;
		14'b00011001100000: color_data = 12'b010000000000;
		14'b00011001100001: color_data = 12'b010000000000;
		14'b00011001100010: color_data = 12'b010000000000;
		14'b00011001100011: color_data = 12'b010000000000;
		14'b00011001100100: color_data = 12'b010000000000;
		14'b00011001100101: color_data = 12'b001000000000;
		14'b00011001100110: color_data = 12'b001000000000;
		14'b00011001100111: color_data = 12'b001000000000;
		14'b00011001101000: color_data = 12'b010000000000;
		14'b00011001101001: color_data = 12'b010000000000;
		14'b00011010001010: color_data = 12'b001000000000;
		14'b00011010001011: color_data = 12'b001000000000;
		14'b00011010001100: color_data = 12'b001000000000;
		14'b00011010001101: color_data = 12'b001000000000;
		14'b00011010001110: color_data = 12'b001000000000;
		14'b00011010001111: color_data = 12'b001000000000;
		14'b00011010010000: color_data = 12'b001000000000;
		14'b00011010010001: color_data = 12'b001000000000;
		14'b00011010010010: color_data = 12'b001000000000;
		14'b00011010010011: color_data = 12'b001000000000;
		14'b00011010010100: color_data = 12'b010000000000;
		14'b00011010010101: color_data = 12'b010000000000;
		14'b00011010010110: color_data = 12'b010000000000;
		14'b00011010010111: color_data = 12'b010000000000;
		14'b00011010011000: color_data = 12'b010000000000;
		14'b00011010011001: color_data = 12'b010000000000;
		14'b00011010011010: color_data = 12'b010000000000;
		14'b00011010011011: color_data = 12'b010000000000;
		14'b00011010011100: color_data = 12'b010000000000;
		14'b00011010011101: color_data = 12'b010000000000;
		14'b00011010011110: color_data = 12'b010000000000;
		14'b00011010011111: color_data = 12'b010000000000;
		14'b00011010100000: color_data = 12'b010000000000;
		14'b00011010100001: color_data = 12'b010000000000;
		14'b00011010100010: color_data = 12'b010000000000;
		14'b00011010100011: color_data = 12'b010000000000;
		14'b00011010100100: color_data = 12'b010000000000;
		14'b00011010100101: color_data = 12'b010000000000;
		14'b00011010100110: color_data = 12'b001000000000;
		14'b00011010100111: color_data = 12'b001000000000;
		14'b00011010101100: color_data = 12'b001000000000;
		14'b00011010101101: color_data = 12'b001000000000;
		14'b00011010101110: color_data = 12'b001000000000;
		14'b00011010101111: color_data = 12'b001000000000;
		14'b00011010110000: color_data = 12'b001000000000;
		14'b00011010110001: color_data = 12'b001000000000;
		14'b00011011011010: color_data = 12'b001000000000;
		14'b00011011011011: color_data = 12'b010000000000;
		14'b00011011011100: color_data = 12'b010000000000;
		14'b00011011011101: color_data = 12'b010000000000;
		14'b00011011011110: color_data = 12'b010000000000;
		14'b00011011011111: color_data = 12'b010000000000;
		14'b00011011100000: color_data = 12'b010000000000;
		14'b00011011100001: color_data = 12'b010000000000;
		14'b00011011100010: color_data = 12'b010000000000;
		14'b00011011100011: color_data = 12'b010000000000;
		14'b00011011100100: color_data = 12'b010000000000;
		14'b00011011100101: color_data = 12'b001000000000;
		14'b00011011100110: color_data = 12'b001000000000;
		14'b00011011100111: color_data = 12'b010000000000;
		14'b00011011101000: color_data = 12'b010000000000;
		14'b00011011101001: color_data = 12'b001000000000;
		14'b00011100001001: color_data = 12'b001000000000;
		14'b00011100001010: color_data = 12'b001000000000;
		14'b00011100001110: color_data = 12'b001000000000;
		14'b00011100001111: color_data = 12'b001000000000;
		14'b00011100010000: color_data = 12'b001000000000;
		14'b00011100010001: color_data = 12'b010000000000;
		14'b00011100010010: color_data = 12'b010000000000;
		14'b00011100010011: color_data = 12'b010000000000;
		14'b00011100010100: color_data = 12'b010000000000;
		14'b00011100010101: color_data = 12'b010000000000;
		14'b00011100010110: color_data = 12'b010000000000;
		14'b00011100010111: color_data = 12'b010000000000;
		14'b00011100011000: color_data = 12'b010000000000;
		14'b00011100011001: color_data = 12'b010000000000;
		14'b00011100011010: color_data = 12'b010000000000;
		14'b00011100011011: color_data = 12'b010000000000;
		14'b00011100011100: color_data = 12'b010000000000;
		14'b00011100011101: color_data = 12'b010000000000;
		14'b00011100011110: color_data = 12'b010000000000;
		14'b00011100011111: color_data = 12'b010000000000;
		14'b00011100100000: color_data = 12'b010000000000;
		14'b00011100100001: color_data = 12'b010000000000;
		14'b00011100100010: color_data = 12'b010000000000;
		14'b00011100100011: color_data = 12'b010000000000;
		14'b00011100100100: color_data = 12'b010000000000;
		14'b00011100100101: color_data = 12'b010000000000;
		14'b00011100100110: color_data = 12'b010000000000;
		14'b00011100100111: color_data = 12'b010000000000;
		14'b00011100101000: color_data = 12'b010000000000;
		14'b00011100101001: color_data = 12'b001000000000;
		14'b00011100101010: color_data = 12'b001000000000;
		14'b00011100101110: color_data = 12'b001000000000;
		14'b00011100101111: color_data = 12'b001000000000;
		14'b00011100110000: color_data = 12'b001000000000;
		14'b00011101011010: color_data = 12'b010000000000;
		14'b00011101011011: color_data = 12'b010000000000;
		14'b00011101011100: color_data = 12'b010000000000;
		14'b00011101011101: color_data = 12'b010000000000;
		14'b00011101011110: color_data = 12'b010000000000;
		14'b00011101011111: color_data = 12'b010000000000;
		14'b00011101100000: color_data = 12'b010000000000;
		14'b00011101100001: color_data = 12'b010000000000;
		14'b00011101100010: color_data = 12'b010000000000;
		14'b00011101100011: color_data = 12'b010000000000;
		14'b00011101100100: color_data = 12'b010000000000;
		14'b00011101100101: color_data = 12'b001000000000;
		14'b00011101100110: color_data = 12'b001000000000;
		14'b00011101100111: color_data = 12'b010000000000;
		14'b00011101101000: color_data = 12'b010000000000;
		14'b00011110001111: color_data = 12'b001000000000;
		14'b00011110010000: color_data = 12'b010000000000;
		14'b00011110010001: color_data = 12'b010000000000;
		14'b00011110010010: color_data = 12'b010000000000;
		14'b00011110010011: color_data = 12'b010000000000;
		14'b00011110010100: color_data = 12'b010000000000;
		14'b00011110010101: color_data = 12'b001000000000;
		14'b00011110010110: color_data = 12'b001000000000;
		14'b00011110010111: color_data = 12'b001000000000;
		14'b00011110011000: color_data = 12'b001000000000;
		14'b00011110011001: color_data = 12'b001000000000;
		14'b00011110011010: color_data = 12'b010000000000;
		14'b00011110011011: color_data = 12'b010000000000;
		14'b00011110011100: color_data = 12'b010000000000;
		14'b00011110011101: color_data = 12'b010000000000;
		14'b00011110011110: color_data = 12'b010000000000;
		14'b00011110011111: color_data = 12'b010000000000;
		14'b00011110100000: color_data = 12'b010000000000;
		14'b00011110100001: color_data = 12'b010000000000;
		14'b00011110100010: color_data = 12'b010000000000;
		14'b00011110100011: color_data = 12'b010000000000;
		14'b00011110100100: color_data = 12'b010000000000;
		14'b00011110100101: color_data = 12'b010000000000;
		14'b00011110100110: color_data = 12'b010000000000;
		14'b00011110100111: color_data = 12'b010000000000;
		14'b00011110101000: color_data = 12'b010000000000;
		14'b00011110101001: color_data = 12'b010000000000;
		14'b00011110101010: color_data = 12'b010000000000;
		14'b00011110101011: color_data = 12'b010000000000;
		14'b00011110101100: color_data = 12'b001000000000;
		14'b00011110101111: color_data = 12'b001000000000;
		14'b00011110110000: color_data = 12'b001000000000;
		14'b00011110110001: color_data = 12'b001000000000;
		14'b00011111011001: color_data = 12'b001000000000;
		14'b00011111011010: color_data = 12'b010000000000;
		14'b00011111011011: color_data = 12'b010000000000;
		14'b00011111011100: color_data = 12'b010000000000;
		14'b00011111011101: color_data = 12'b010000000000;
		14'b00011111011110: color_data = 12'b010000000000;
		14'b00011111011111: color_data = 12'b010000000000;
		14'b00011111100000: color_data = 12'b010000000000;
		14'b00011111100001: color_data = 12'b010000000000;
		14'b00011111100010: color_data = 12'b010000000000;
		14'b00011111100011: color_data = 12'b010000000000;
		14'b00011111100100: color_data = 12'b001000000000;
		14'b00011111100101: color_data = 12'b001000000000;
		14'b00011111100110: color_data = 12'b010000000000;
		14'b00011111100111: color_data = 12'b010000000000;
		14'b00011111101000: color_data = 12'b001000000000;
		14'b00100000001110: color_data = 12'b001000000000;
		14'b00100000001111: color_data = 12'b001000000000;
		14'b00100000010000: color_data = 12'b001000000000;
		14'b00100000010001: color_data = 12'b001000000000;
		14'b00100000010010: color_data = 12'b001000000000;
		14'b00100000010011: color_data = 12'b001000000000;
		14'b00100000010100: color_data = 12'b001000000000;
		14'b00100000010111: color_data = 12'b001000000000;
		14'b00100000011000: color_data = 12'b001000000000;
		14'b00100000011001: color_data = 12'b010000000000;
		14'b00100000011010: color_data = 12'b010000000000;
		14'b00100000011011: color_data = 12'b010000000000;
		14'b00100000011100: color_data = 12'b010000000000;
		14'b00100000011101: color_data = 12'b010000000000;
		14'b00100000011110: color_data = 12'b010000000000;
		14'b00100000011111: color_data = 12'b001000000000;
		14'b00100000100000: color_data = 12'b001000000000;
		14'b00100000100100: color_data = 12'b001000000000;
		14'b00100000100101: color_data = 12'b010000000000;
		14'b00100000100110: color_data = 12'b010000000000;
		14'b00100000100111: color_data = 12'b001000000000;
		14'b00100000101000: color_data = 12'b010000000000;
		14'b00100000101001: color_data = 12'b010000000000;
		14'b00100000101010: color_data = 12'b010000000000;
		14'b00100000101011: color_data = 12'b010000000000;
		14'b00100000101100: color_data = 12'b010000000000;
		14'b00100000101101: color_data = 12'b010000000000;
		14'b00100000101110: color_data = 12'b001000000000;
		14'b00100000101111: color_data = 12'b001000000000;
		14'b00100000110000: color_data = 12'b001000000000;
		14'b00100000110001: color_data = 12'b010000000000;
		14'b00100000110010: color_data = 12'b010000000000;
		14'b00100000110011: color_data = 12'b001000000000;
		14'b00100001011001: color_data = 12'b010000000000;
		14'b00100001011010: color_data = 12'b010000000000;
		14'b00100001011011: color_data = 12'b010000000000;
		14'b00100001011100: color_data = 12'b010000000000;
		14'b00100001011101: color_data = 12'b010000000000;
		14'b00100001011110: color_data = 12'b010000000000;
		14'b00100001011111: color_data = 12'b010000000000;
		14'b00100001100000: color_data = 12'b010000000000;
		14'b00100001100001: color_data = 12'b010000000000;
		14'b00100001100010: color_data = 12'b010000000000;
		14'b00100001100011: color_data = 12'b010000000000;
		14'b00100001100100: color_data = 12'b001000000000;
		14'b00100001100101: color_data = 12'b001000000000;
		14'b00100001100110: color_data = 12'b010000000000;
		14'b00100001100111: color_data = 12'b010000000000;
		14'b00100010001101: color_data = 12'b001000000000;
		14'b00100010001110: color_data = 12'b001000000000;
		14'b00100010010110: color_data = 12'b001000000000;
		14'b00100010010111: color_data = 12'b001000000000;
		14'b00100010011000: color_data = 12'b010000000000;
		14'b00100010011001: color_data = 12'b010000000000;
		14'b00100010011010: color_data = 12'b010000000000;
		14'b00100010011011: color_data = 12'b010000000000;
		14'b00100010011100: color_data = 12'b010000000000;
		14'b00100010011101: color_data = 12'b001000000000;
		14'b00100010100100: color_data = 12'b001000000000;
		14'b00100010100101: color_data = 12'b010000000000;
		14'b00100010100110: color_data = 12'b010000000000;
		14'b00100010100111: color_data = 12'b001000000000;
		14'b00100010101001: color_data = 12'b001000000000;
		14'b00100010101010: color_data = 12'b001000000000;
		14'b00100010101011: color_data = 12'b010000000000;
		14'b00100010101100: color_data = 12'b010000000000;
		14'b00100010101101: color_data = 12'b010000000000;
		14'b00100010101110: color_data = 12'b010000000000;
		14'b00100010101111: color_data = 12'b010000000000;
		14'b00100010110000: color_data = 12'b001000000000;
		14'b00100010110001: color_data = 12'b001000000000;
		14'b00100010110010: color_data = 12'b001000000000;
		14'b00100010110011: color_data = 12'b010000000000;
		14'b00100010110100: color_data = 12'b001000000000;
		14'b00100011011001: color_data = 12'b001000000000;
		14'b00100011011010: color_data = 12'b010000000000;
		14'b00100011011011: color_data = 12'b010000000000;
		14'b00100011011100: color_data = 12'b010000000000;
		14'b00100011011101: color_data = 12'b010000000000;
		14'b00100011011110: color_data = 12'b010000000000;
		14'b00100011011111: color_data = 12'b010000000000;
		14'b00100011100000: color_data = 12'b010000000000;
		14'b00100011100001: color_data = 12'b010000000000;
		14'b00100011100010: color_data = 12'b010000000000;
		14'b00100011100011: color_data = 12'b001000000000;
		14'b00100011100100: color_data = 12'b001000000000;
		14'b00100011100101: color_data = 12'b010000000000;
		14'b00100011100110: color_data = 12'b010000000000;
		14'b00100011100111: color_data = 12'b001000000000;
		14'b00100100010100: color_data = 12'b001000000000;
		14'b00100100010101: color_data = 12'b001000000000;
		14'b00100100010110: color_data = 12'b010000000000;
		14'b00100100010111: color_data = 12'b010000000000;
		14'b00100100011000: color_data = 12'b010000000000;
		14'b00100100011001: color_data = 12'b010000000000;
		14'b00100100011010: color_data = 12'b010000000000;
		14'b00100100011011: color_data = 12'b010000000000;
		14'b00100100011100: color_data = 12'b001000000000;
		14'b00100100011101: color_data = 12'b001000000000;
		14'b00100100100000: color_data = 12'b001000000000;
		14'b00100100100001: color_data = 12'b001000000000;
		14'b00100100100010: color_data = 12'b001000000000;
		14'b00100100100011: color_data = 12'b010000000000;
		14'b00100100100100: color_data = 12'b010000000000;
		14'b00100100100101: color_data = 12'b010000000000;
		14'b00100100100110: color_data = 12'b010000000000;
		14'b00100100100111: color_data = 12'b010000000000;
		14'b00100100101011: color_data = 12'b001000000000;
		14'b00100100101100: color_data = 12'b010000000000;
		14'b00100100101101: color_data = 12'b010000000000;
		14'b00100100101110: color_data = 12'b010000000000;
		14'b00100100101111: color_data = 12'b010000000000;
		14'b00100100110000: color_data = 12'b010000000000;
		14'b00100100110001: color_data = 12'b001000000000;
		14'b00100100110010: color_data = 12'b001000000000;
		14'b00100100110011: color_data = 12'b001000000000;
		14'b00100100110100: color_data = 12'b001000000000;
		14'b00100100110101: color_data = 12'b001000000000;
		14'b00100101011001: color_data = 12'b001000000000;
		14'b00100101011010: color_data = 12'b010000000000;
		14'b00100101011011: color_data = 12'b010000000000;
		14'b00100101011100: color_data = 12'b010000000000;
		14'b00100101011101: color_data = 12'b010000000000;
		14'b00100101011110: color_data = 12'b010000000000;
		14'b00100101011111: color_data = 12'b010000000000;
		14'b00100101100000: color_data = 12'b010000000000;
		14'b00100101100001: color_data = 12'b010000000000;
		14'b00100101100010: color_data = 12'b001000000000;
		14'b00100101100011: color_data = 12'b001000000000;
		14'b00100101100100: color_data = 12'b010000000000;
		14'b00100101100101: color_data = 12'b010000000000;
		14'b00100101100110: color_data = 12'b001000000000;
		14'b00100110010100: color_data = 12'b010000000000;
		14'b00100110010101: color_data = 12'b010000000000;
		14'b00100110010110: color_data = 12'b010000000000;
		14'b00100110010111: color_data = 12'b010000000000;
		14'b00100110011000: color_data = 12'b010000000000;
		14'b00100110011001: color_data = 12'b010000000000;
		14'b00100110011010: color_data = 12'b010000000000;
		14'b00100110011011: color_data = 12'b010000000000;
		14'b00100110011100: color_data = 12'b010000000000;
		14'b00100110011101: color_data = 12'b010000000000;
		14'b00100110011110: color_data = 12'b010000000000;
		14'b00100110011111: color_data = 12'b010000000000;
		14'b00100110100000: color_data = 12'b010000000000;
		14'b00100110100001: color_data = 12'b010000000000;
		14'b00100110100010: color_data = 12'b001000000000;
		14'b00100110100011: color_data = 12'b001000000000;
		14'b00100110100100: color_data = 12'b010000000000;
		14'b00100110100101: color_data = 12'b010000000000;
		14'b00100110100110: color_data = 12'b010000000000;
		14'b00100110100111: color_data = 12'b010000000000;
		14'b00100110101000: color_data = 12'b010000000000;
		14'b00100110101001: color_data = 12'b010000000000;
		14'b00100110101011: color_data = 12'b001000000000;
		14'b00100110101100: color_data = 12'b010000000000;
		14'b00100110101101: color_data = 12'b010000000000;
		14'b00100110101110: color_data = 12'b010000000000;
		14'b00100110101111: color_data = 12'b010000000000;
		14'b00100110110000: color_data = 12'b010000000000;
		14'b00100110110001: color_data = 12'b010000000000;
		14'b00100110110010: color_data = 12'b010000000000;
		14'b00100110110011: color_data = 12'b001000000000;
		14'b00100110110101: color_data = 12'b001000000000;
		14'b00100111011001: color_data = 12'b001000000000;
		14'b00100111011010: color_data = 12'b010000000000;
		14'b00100111011011: color_data = 12'b010000000000;
		14'b00100111011100: color_data = 12'b010000000000;
		14'b00100111011101: color_data = 12'b010000000000;
		14'b00100111011110: color_data = 12'b010000000000;
		14'b00100111011111: color_data = 12'b010000000000;
		14'b00100111100000: color_data = 12'b010000000000;
		14'b00100111100001: color_data = 12'b010000000000;
		14'b00100111100010: color_data = 12'b001000000000;
		14'b00100111100011: color_data = 12'b001000000000;
		14'b00100111100100: color_data = 12'b010000000000;
		14'b00100111100101: color_data = 12'b010000000000;
		14'b00100111100110: color_data = 12'b001000000000;
		14'b00101000010010: color_data = 12'b010000000000;
		14'b00101000010011: color_data = 12'b010000000000;
		14'b00101000010100: color_data = 12'b010000000000;
		14'b00101000010101: color_data = 12'b010000000000;
		14'b00101000010110: color_data = 12'b010000000000;
		14'b00101000010111: color_data = 12'b010000000000;
		14'b00101000011000: color_data = 12'b010000000000;
		14'b00101000011001: color_data = 12'b010000000000;
		14'b00101000011010: color_data = 12'b010000000000;
		14'b00101000011011: color_data = 12'b010000000000;
		14'b00101000011100: color_data = 12'b010000000000;
		14'b00101000011101: color_data = 12'b010000000000;
		14'b00101000011110: color_data = 12'b010000000000;
		14'b00101000011111: color_data = 12'b010000000000;
		14'b00101000100000: color_data = 12'b001000000000;
		14'b00101000100001: color_data = 12'b001000000000;
		14'b00101000100100: color_data = 12'b001000000000;
		14'b00101000100101: color_data = 12'b010000000000;
		14'b00101000100110: color_data = 12'b010000000000;
		14'b00101000100111: color_data = 12'b010000000000;
		14'b00101000101000: color_data = 12'b010000000000;
		14'b00101000101001: color_data = 12'b010000000000;
		14'b00101000101010: color_data = 12'b010000000000;
		14'b00101000101011: color_data = 12'b010000000000;
		14'b00101000101100: color_data = 12'b010000000000;
		14'b00101000101101: color_data = 12'b010000000000;
		14'b00101000101110: color_data = 12'b010000000000;
		14'b00101000101111: color_data = 12'b010000000000;
		14'b00101000110000: color_data = 12'b010000000000;
		14'b00101000110001: color_data = 12'b001000000000;
		14'b00101000110010: color_data = 12'b010000000000;
		14'b00101000110011: color_data = 12'b010000000000;
		14'b00101001010010: color_data = 12'b001000000000;
		14'b00101001011001: color_data = 12'b001000000000;
		14'b00101001011010: color_data = 12'b010000000000;
		14'b00101001011011: color_data = 12'b010000000000;
		14'b00101001011100: color_data = 12'b010000000000;
		14'b00101001011101: color_data = 12'b010000000000;
		14'b00101001011110: color_data = 12'b010000000000;
		14'b00101001011111: color_data = 12'b010000000000;
		14'b00101001100000: color_data = 12'b010000000000;
		14'b00101001100001: color_data = 12'b001000000000;
		14'b00101001100010: color_data = 12'b001000000000;
		14'b00101001100011: color_data = 12'b010000000000;
		14'b00101001100100: color_data = 12'b010000000000;
		14'b00101001100101: color_data = 12'b010000000000;
		14'b00101010010000: color_data = 12'b001000000000;
		14'b00101010010001: color_data = 12'b010000000000;
		14'b00101010010010: color_data = 12'b010000000000;
		14'b00101010010011: color_data = 12'b010000000000;
		14'b00101010010100: color_data = 12'b010000000000;
		14'b00101010010101: color_data = 12'b010000000000;
		14'b00101010010110: color_data = 12'b010000000000;
		14'b00101010010111: color_data = 12'b010000000000;
		14'b00101010011000: color_data = 12'b010000000000;
		14'b00101010011001: color_data = 12'b010000000000;
		14'b00101010011010: color_data = 12'b001000000000;
		14'b00101010011011: color_data = 12'b001000000000;
		14'b00101010011100: color_data = 12'b001000000000;
		14'b00101010011101: color_data = 12'b001000000000;
		14'b00101010011110: color_data = 12'b001000000000;
		14'b00101010100100: color_data = 12'b001000000000;
		14'b00101010100101: color_data = 12'b001000000000;
		14'b00101010100110: color_data = 12'b010000000000;
		14'b00101010100111: color_data = 12'b010000000000;
		14'b00101010101000: color_data = 12'b010000000000;
		14'b00101010101001: color_data = 12'b010000000000;
		14'b00101010101010: color_data = 12'b010000000000;
		14'b00101010101011: color_data = 12'b010000000000;
		14'b00101010101100: color_data = 12'b010000000000;
		14'b00101010101101: color_data = 12'b010000000000;
		14'b00101010101110: color_data = 12'b010000000000;
		14'b00101010101111: color_data = 12'b010000000000;
		14'b00101010110000: color_data = 12'b010000000000;
		14'b00101010110001: color_data = 12'b001000000000;
		14'b00101010110010: color_data = 12'b001000000000;
		14'b00101010110011: color_data = 12'b010000000000;
		14'b00101010110100: color_data = 12'b010000000000;
		14'b00101011011001: color_data = 12'b001000000000;
		14'b00101011011010: color_data = 12'b010000000000;
		14'b00101011011011: color_data = 12'b010000000000;
		14'b00101011011100: color_data = 12'b010000000000;
		14'b00101011011101: color_data = 12'b010000000000;
		14'b00101011011110: color_data = 12'b010000000000;
		14'b00101011011111: color_data = 12'b010000000000;
		14'b00101011100000: color_data = 12'b001000000000;
		14'b00101011100001: color_data = 12'b001000000000;
		14'b00101011100010: color_data = 12'b001000000000;
		14'b00101011100011: color_data = 12'b010000000000;
		14'b00101011100100: color_data = 12'b010000000000;
		14'b00101011100101: color_data = 12'b001000000000;
		14'b00101100001111: color_data = 12'b001000000000;
		14'b00101100010000: color_data = 12'b010000000000;
		14'b00101100010001: color_data = 12'b010000000000;
		14'b00101100010010: color_data = 12'b010000000000;
		14'b00101100010011: color_data = 12'b010000000000;
		14'b00101100010100: color_data = 12'b010000000000;
		14'b00101100010101: color_data = 12'b010000000000;
		14'b00101100010110: color_data = 12'b001000000000;
		14'b00101100010111: color_data = 12'b001000000000;
		14'b00101100011000: color_data = 12'b001000000000;
		14'b00101100011001: color_data = 12'b001000000000;
		14'b00101100100101: color_data = 12'b001000000000;
		14'b00101100100110: color_data = 12'b001000000000;
		14'b00101100100111: color_data = 12'b001000000000;
		14'b00101100101000: color_data = 12'b010000000000;
		14'b00101100101001: color_data = 12'b010000000000;
		14'b00101100101010: color_data = 12'b010000000000;
		14'b00101100101011: color_data = 12'b010000000000;
		14'b00101100101100: color_data = 12'b010000000000;
		14'b00101100101101: color_data = 12'b010000000000;
		14'b00101100101110: color_data = 12'b010000000000;
		14'b00101100101111: color_data = 12'b010000000000;
		14'b00101100110000: color_data = 12'b010000000000;
		14'b00101100110001: color_data = 12'b001000000000;
		14'b00101100110011: color_data = 12'b001000000000;
		14'b00101100110100: color_data = 12'b010000000000;
		14'b00101100110101: color_data = 12'b010000000000;
		14'b00101101011001: color_data = 12'b010000000000;
		14'b00101101011010: color_data = 12'b010000000000;
		14'b00101101011011: color_data = 12'b010000000000;
		14'b00101101011100: color_data = 12'b010000000000;
		14'b00101101011101: color_data = 12'b010000000000;
		14'b00101101011110: color_data = 12'b010000000000;
		14'b00101101011111: color_data = 12'b010000000000;
		14'b00101101100000: color_data = 12'b001000000000;
		14'b00101101100001: color_data = 12'b001000000000;
		14'b00101101100010: color_data = 12'b010000000000;
		14'b00101101100011: color_data = 12'b010000000000;
		14'b00101101100100: color_data = 12'b010000000000;
		14'b00101101100101: color_data = 12'b001000000000;
		14'b00101110001110: color_data = 12'b001000000000;
		14'b00101110001111: color_data = 12'b010000000000;
		14'b00101110010000: color_data = 12'b010000000000;
		14'b00101110010001: color_data = 12'b010000000000;
		14'b00101110010010: color_data = 12'b010000000000;
		14'b00101110010011: color_data = 12'b010000000000;
		14'b00101110010100: color_data = 12'b010000000000;
		14'b00101110010101: color_data = 12'b001000000000;
		14'b00101110100101: color_data = 12'b001000000000;
		14'b00101110100110: color_data = 12'b001000000000;
		14'b00101110100111: color_data = 12'b001000000000;
		14'b00101110101000: color_data = 12'b001000000000;
		14'b00101110101001: color_data = 12'b010000000000;
		14'b00101110101010: color_data = 12'b010000000000;
		14'b00101110101011: color_data = 12'b001000000000;
		14'b00101110101100: color_data = 12'b001000000000;
		14'b00101110101101: color_data = 12'b010000000000;
		14'b00101110101110: color_data = 12'b010000000000;
		14'b00101110101111: color_data = 12'b001000000000;
		14'b00101110110000: color_data = 12'b010000000000;
		14'b00101110110001: color_data = 12'b010000000000;
		14'b00101110110100: color_data = 12'b001000000000;
		14'b00101110110101: color_data = 12'b010000000000;
		14'b00101110110110: color_data = 12'b001000000000;
		14'b00101111011001: color_data = 12'b010000000000;
		14'b00101111011010: color_data = 12'b010000000000;
		14'b00101111011011: color_data = 12'b010000000000;
		14'b00101111011100: color_data = 12'b010000000000;
		14'b00101111011101: color_data = 12'b010000000000;
		14'b00101111011110: color_data = 12'b010000000000;
		14'b00101111011111: color_data = 12'b001000000000;
		14'b00101111100000: color_data = 12'b001000000000;
		14'b00101111100001: color_data = 12'b010000000000;
		14'b00101111100010: color_data = 12'b010000000000;
		14'b00101111100011: color_data = 12'b010000000000;
		14'b00101111100100: color_data = 12'b010000000000;
		14'b00110000001101: color_data = 12'b001000000000;
		14'b00110000001110: color_data = 12'b001000000000;
		14'b00110000001111: color_data = 12'b010000000000;
		14'b00110000010000: color_data = 12'b010000000000;
		14'b00110000010001: color_data = 12'b010000000000;
		14'b00110000011111: color_data = 12'b001000000000;
		14'b00110000100111: color_data = 12'b001000000000;
		14'b00110000101000: color_data = 12'b001000000000;
		14'b00110000101001: color_data = 12'b010000000000;
		14'b00110000101010: color_data = 12'b010000000000;
		14'b00110000101011: color_data = 12'b001000000000;
		14'b00110000101100: color_data = 12'b001000000000;
		14'b00110000101111: color_data = 12'b001000000000;
		14'b00110000110000: color_data = 12'b001000000000;
		14'b00110000110001: color_data = 12'b010000000000;
		14'b00110000110010: color_data = 12'b001000000000;
		14'b00110000110110: color_data = 12'b001000000000;
		14'b00110001011000: color_data = 12'b001000000000;
		14'b00110001011001: color_data = 12'b010000000000;
		14'b00110001011010: color_data = 12'b010000000000;
		14'b00110001011011: color_data = 12'b010000000000;
		14'b00110001011100: color_data = 12'b010000000000;
		14'b00110001011101: color_data = 12'b010000000000;
		14'b00110001011110: color_data = 12'b010000000000;
		14'b00110001011111: color_data = 12'b001000000000;
		14'b00110001100000: color_data = 12'b001000000000;
		14'b00110001100001: color_data = 12'b010000000000;
		14'b00110001100010: color_data = 12'b010000000000;
		14'b00110001100011: color_data = 12'b010000000000;
		14'b00110010001010: color_data = 12'b001000000000;
		14'b00110010001011: color_data = 12'b001000000000;
		14'b00110010001100: color_data = 12'b001000000000;
		14'b00110010001101: color_data = 12'b001000000000;
		14'b00110010001110: color_data = 12'b010000000000;
		14'b00110010001111: color_data = 12'b010000000000;
		14'b00110010010000: color_data = 12'b010000000000;
		14'b00110010100010: color_data = 12'b001000000000;
		14'b00110010100011: color_data = 12'b001000000000;
		14'b00110010101000: color_data = 12'b001000000000;
		14'b00110010101001: color_data = 12'b001000000000;
		14'b00110010101010: color_data = 12'b001000000000;
		14'b00110010101111: color_data = 12'b001000000000;
		14'b00110010110000: color_data = 12'b001000000000;
		14'b00110010110001: color_data = 12'b010000000000;
		14'b00110010110010: color_data = 12'b001000000000;
		14'b00110010110110: color_data = 12'b001000000000;
		14'b00110010110111: color_data = 12'b001000000000;
		14'b00110011011000: color_data = 12'b001000000000;
		14'b00110011011001: color_data = 12'b010000000000;
		14'b00110011011010: color_data = 12'b010000000000;
		14'b00110011011011: color_data = 12'b010000000000;
		14'b00110011011100: color_data = 12'b010000000000;
		14'b00110011011101: color_data = 12'b010000000000;
		14'b00110011011110: color_data = 12'b001000000000;
		14'b00110011011111: color_data = 12'b001000000000;
		14'b00110011100000: color_data = 12'b001000000000;
		14'b00110011100001: color_data = 12'b010000000000;
		14'b00110011100010: color_data = 12'b010000000000;
		14'b00110011100011: color_data = 12'b010000000000;
		14'b00110011100110: color_data = 12'b001000000000;
		14'b00110011111011: color_data = 12'b001000000000;
		14'b00110100001010: color_data = 12'b001000000000;
		14'b00110100001011: color_data = 12'b001000000000;
		14'b00110100001100: color_data = 12'b001000000000;
		14'b00110100001101: color_data = 12'b010000000000;
		14'b00110100001110: color_data = 12'b010000000000;
		14'b00110100001111: color_data = 12'b010000000000;
		14'b00110100010000: color_data = 12'b001000000000;
		14'b00110100101111: color_data = 12'b001000000000;
		14'b00110100110000: color_data = 12'b010000000000;
		14'b00110100110001: color_data = 12'b010000000000;
		14'b00110100110010: color_data = 12'b010000000000;
		14'b00110100110011: color_data = 12'b001000000000;
		14'b00110100110111: color_data = 12'b001000000000;
		14'b00110101010111: color_data = 12'b001000000000;
		14'b00110101011000: color_data = 12'b010000000000;
		14'b00110101011001: color_data = 12'b010000000000;
		14'b00110101011010: color_data = 12'b010000000000;
		14'b00110101011011: color_data = 12'b010000000000;
		14'b00110101011100: color_data = 12'b010000000000;
		14'b00110101011101: color_data = 12'b010000000000;
		14'b00110101011110: color_data = 12'b001000000000;
		14'b00110101011111: color_data = 12'b001000000000;
		14'b00110101100000: color_data = 12'b010000000000;
		14'b00110101100001: color_data = 12'b010000000000;
		14'b00110101100010: color_data = 12'b010000000000;
		14'b00110101100011: color_data = 12'b010000000000;
		14'b00110101100100: color_data = 12'b001000000000;
		14'b00110101100101: color_data = 12'b001000000000;
		14'b00110101100110: color_data = 12'b001000000000;
		14'b00110101111010: color_data = 12'b001000000000;
		14'b00110101111011: color_data = 12'b001000000000;
		14'b00110110001001: color_data = 12'b001000000000;
		14'b00110110001010: color_data = 12'b001000000000;
		14'b00110110001011: color_data = 12'b001000000000;
		14'b00110110001100: color_data = 12'b010000000000;
		14'b00110110001101: color_data = 12'b010000000000;
		14'b00110110001110: color_data = 12'b010000000000;
		14'b00110110001111: color_data = 12'b001000000000;
		14'b00110110010000: color_data = 12'b001000000000;
		14'b00110110100101: color_data = 12'b001000000000;
		14'b00110110100110: color_data = 12'b001000000000;
		14'b00110110101110: color_data = 12'b001000000000;
		14'b00110110101111: color_data = 12'b010000000000;
		14'b00110110110000: color_data = 12'b010000000000;
		14'b00110110110001: color_data = 12'b010000000000;
		14'b00110110110010: color_data = 12'b010000000000;
		14'b00110110110011: color_data = 12'b001000000000;
		14'b00110110110111: color_data = 12'b001000000000;
		14'b00110111010111: color_data = 12'b001000000000;
		14'b00110111011000: color_data = 12'b010000000000;
		14'b00110111011001: color_data = 12'b010000000000;
		14'b00110111011010: color_data = 12'b010000000000;
		14'b00110111011011: color_data = 12'b010000000000;
		14'b00110111011100: color_data = 12'b010000000000;
		14'b00110111011101: color_data = 12'b001000000000;
		14'b00110111011110: color_data = 12'b001000000000;
		14'b00110111011111: color_data = 12'b001000000000;
		14'b00110111100000: color_data = 12'b010000000000;
		14'b00110111100001: color_data = 12'b010000000000;
		14'b00110111100010: color_data = 12'b010000000000;
		14'b00110111100011: color_data = 12'b010000000000;
		14'b00110111100100: color_data = 12'b001000000000;
		14'b00110111100101: color_data = 12'b001000000000;
		14'b00110111100110: color_data = 12'b001000000000;
		14'b00110111111001: color_data = 12'b001000000000;
		14'b00110111111010: color_data = 12'b001000000000;
		14'b00110111111011: color_data = 12'b001000000000;
		14'b00111000001001: color_data = 12'b001000000000;
		14'b00111000001010: color_data = 12'b001000000000;
		14'b00111000001011: color_data = 12'b010000000000;
		14'b00111000001100: color_data = 12'b010000000000;
		14'b00111000001101: color_data = 12'b001000000000;
		14'b00111000001111: color_data = 12'b001000000000;
		14'b00111000010000: color_data = 12'b001000000000;
		14'b00111000100101: color_data = 12'b001000000000;
		14'b00111000100110: color_data = 12'b010000000000;
		14'b00111000100111: color_data = 12'b001000000000;
		14'b00111000101101: color_data = 12'b001000000000;
		14'b00111000101110: color_data = 12'b001000000000;
		14'b00111000101111: color_data = 12'b010000000000;
		14'b00111000110000: color_data = 12'b010000000000;
		14'b00111000110001: color_data = 12'b010000000000;
		14'b00111000110010: color_data = 12'b010000000000;
		14'b00111000110011: color_data = 12'b001000000000;
		14'b00111000110111: color_data = 12'b001000000000;
		14'b00111001010110: color_data = 12'b001000000000;
		14'b00111001010111: color_data = 12'b010000000000;
		14'b00111001011000: color_data = 12'b010000000000;
		14'b00111001011001: color_data = 12'b010000000000;
		14'b00111001011010: color_data = 12'b010000000000;
		14'b00111001011011: color_data = 12'b010000000000;
		14'b00111001011100: color_data = 12'b001000000000;
		14'b00111001011101: color_data = 12'b001000000000;
		14'b00111001011110: color_data = 12'b001000000000;
		14'b00111001011111: color_data = 12'b010000000000;
		14'b00111001100000: color_data = 12'b010000000000;
		14'b00111001100001: color_data = 12'b010000000000;
		14'b00111001100010: color_data = 12'b010000000000;
		14'b00111001100011: color_data = 12'b010000000000;
		14'b00111001100100: color_data = 12'b001000000000;
		14'b00111001100101: color_data = 12'b001000000000;
		14'b00111001100110: color_data = 12'b001000000000;
		14'b00111001111000: color_data = 12'b001000000000;
		14'b00111001111001: color_data = 12'b001000000000;
		14'b00111001111010: color_data = 12'b001000000000;
		14'b00111001111011: color_data = 12'b001000000000;
		14'b00111010001001: color_data = 12'b001000000000;
		14'b00111010001010: color_data = 12'b001000000000;
		14'b00111010001011: color_data = 12'b001000000000;
		14'b00111010001100: color_data = 12'b001000000000;
		14'b00111010001101: color_data = 12'b001000000000;
		14'b00111010001111: color_data = 12'b001000000000;
		14'b00111010010000: color_data = 12'b001000000000;
		14'b00111010101100: color_data = 12'b001000000000;
		14'b00111010101101: color_data = 12'b001000000000;
		14'b00111010101110: color_data = 12'b010000000000;
		14'b00111010101111: color_data = 12'b010000000000;
		14'b00111010110000: color_data = 12'b010000000000;
		14'b00111010110001: color_data = 12'b010000000000;
		14'b00111010110010: color_data = 12'b010000000000;
		14'b00111010110011: color_data = 12'b001000000000;
		14'b00111011010101: color_data = 12'b001000000000;
		14'b00111011010110: color_data = 12'b010000000000;
		14'b00111011010111: color_data = 12'b010000000000;
		14'b00111011011000: color_data = 12'b010000000000;
		14'b00111011011001: color_data = 12'b010000000000;
		14'b00111011011010: color_data = 12'b010000000000;
		14'b00111011011011: color_data = 12'b010000000000;
		14'b00111011011100: color_data = 12'b001000000000;
		14'b00111011011101: color_data = 12'b001000000000;
		14'b00111011011110: color_data = 12'b001000000000;
		14'b00111011011111: color_data = 12'b010000000000;
		14'b00111011100000: color_data = 12'b010000000000;
		14'b00111011100001: color_data = 12'b010000000000;
		14'b00111011100010: color_data = 12'b010000000000;
		14'b00111011100011: color_data = 12'b010000000000;
		14'b00111011100100: color_data = 12'b001000000000;
		14'b00111011100101: color_data = 12'b001000000000;
		14'b00111011100110: color_data = 12'b001000000000;
		14'b00111011110111: color_data = 12'b001000000000;
		14'b00111011111000: color_data = 12'b001000000000;
		14'b00111011111001: color_data = 12'b001000000000;
		14'b00111011111010: color_data = 12'b001000000000;
		14'b00111011111011: color_data = 12'b001000000000;
		14'b00111100001001: color_data = 12'b001000000000;
		14'b00111100001010: color_data = 12'b001000000000;
		14'b00111100001011: color_data = 12'b001000000000;
		14'b00111100001100: color_data = 12'b001000000000;
		14'b00111100001101: color_data = 12'b001000000000;
		14'b00111100010000: color_data = 12'b001000000000;
		14'b00111100010001: color_data = 12'b001000000000;
		14'b00111100101011: color_data = 12'b001000000000;
		14'b00111100101100: color_data = 12'b001000000000;
		14'b00111100101101: color_data = 12'b010000000000;
		14'b00111100101110: color_data = 12'b010000000000;
		14'b00111100101111: color_data = 12'b010000000000;
		14'b00111100110000: color_data = 12'b010000000000;
		14'b00111100110001: color_data = 12'b010000000000;
		14'b00111100110010: color_data = 12'b001000000000;
		14'b00111100110011: color_data = 12'b001000000000;
		14'b00111101010100: color_data = 12'b001000000000;
		14'b00111101010101: color_data = 12'b010000000000;
		14'b00111101010110: color_data = 12'b010000000000;
		14'b00111101010111: color_data = 12'b010000000000;
		14'b00111101011000: color_data = 12'b010000000000;
		14'b00111101011001: color_data = 12'b010000000000;
		14'b00111101011010: color_data = 12'b010000000000;
		14'b00111101011011: color_data = 12'b010000000000;
		14'b00111101011100: color_data = 12'b001000000000;
		14'b00111101011101: color_data = 12'b001000000000;
		14'b00111101011110: color_data = 12'b001000000000;
		14'b00111101011111: color_data = 12'b010000000000;
		14'b00111101100000: color_data = 12'b010000000000;
		14'b00111101100001: color_data = 12'b010000000000;
		14'b00111101100010: color_data = 12'b010000000000;
		14'b00111101100011: color_data = 12'b010000000000;
		14'b00111101100100: color_data = 12'b001000000000;
		14'b00111101100101: color_data = 12'b001000000000;
		14'b00111101100110: color_data = 12'b001000000000;
		14'b00111101100111: color_data = 12'b001000000000;
		14'b00111101111000: color_data = 12'b001000000000;
		14'b00111101111001: color_data = 12'b001000000000;
		14'b00111101111010: color_data = 12'b001000000000;
		14'b00111101111011: color_data = 12'b001000000000;
		14'b00111110001001: color_data = 12'b001000000000;
		14'b00111110001010: color_data = 12'b001000000000;
		14'b00111110001011: color_data = 12'b001000000000;
		14'b00111110001100: color_data = 12'b001000000000;
		14'b00111110001101: color_data = 12'b001000000000;
		14'b00111110010001: color_data = 12'b001000000000;
		14'b00111110010010: color_data = 12'b001000000000;
		14'b00111110101001: color_data = 12'b001000000000;
		14'b00111110101010: color_data = 12'b001000000000;
		14'b00111110101011: color_data = 12'b001000000000;
		14'b00111110101100: color_data = 12'b010000000000;
		14'b00111110101101: color_data = 12'b010000000000;
		14'b00111110101110: color_data = 12'b010000000000;
		14'b00111110101111: color_data = 12'b010000000000;
		14'b00111110110000: color_data = 12'b010000000000;
		14'b00111110110001: color_data = 12'b010000000000;
		14'b00111110110010: color_data = 12'b001000000000;
		14'b00111111010011: color_data = 12'b001000000000;
		14'b00111111010100: color_data = 12'b010000000000;
		14'b00111111010101: color_data = 12'b001000000000;
		14'b00111111010110: color_data = 12'b001000000000;
		14'b00111111010111: color_data = 12'b001000000000;
		14'b00111111011000: color_data = 12'b001000000000;
		14'b00111111011001: color_data = 12'b010000000000;
		14'b00111111011010: color_data = 12'b010000000000;
		14'b00111111011011: color_data = 12'b010000000000;
		14'b00111111011100: color_data = 12'b001000000000;
		14'b00111111011101: color_data = 12'b001000000000;
		14'b00111111011110: color_data = 12'b001000000000;
		14'b00111111011111: color_data = 12'b010000000000;
		14'b00111111100000: color_data = 12'b010000000000;
		14'b00111111100001: color_data = 12'b010000000000;
		14'b00111111100010: color_data = 12'b010000000000;
		14'b00111111100011: color_data = 12'b010000000000;
		14'b00111111100100: color_data = 12'b001000000000;
		14'b00111111100101: color_data = 12'b001000000000;
		14'b00111111100110: color_data = 12'b001000000000;
		14'b00111111100111: color_data = 12'b001000000000;
		14'b00111111111000: color_data = 12'b001000000000;
		14'b00111111111001: color_data = 12'b001000000000;
		14'b00111111111010: color_data = 12'b001000000000;
		14'b00111111111011: color_data = 12'b001000000000;
		14'b01000000001010: color_data = 12'b001000000000;
		14'b01000000001011: color_data = 12'b001000000000;
		14'b01000000001100: color_data = 12'b001000000000;
		14'b01000000001101: color_data = 12'b001000000000;
		14'b01000000010010: color_data = 12'b001000000000;
		14'b01000000010011: color_data = 12'b001000000000;
		14'b01000000010100: color_data = 12'b001000000000;
		14'b01000000010101: color_data = 12'b001000000000;
		14'b01000000100111: color_data = 12'b001000000000;
		14'b01000000101000: color_data = 12'b001000000000;
		14'b01000000101001: color_data = 12'b001000000000;
		14'b01000000101010: color_data = 12'b010000000000;
		14'b01000000101011: color_data = 12'b010000000000;
		14'b01000000101100: color_data = 12'b010000000000;
		14'b01000000101101: color_data = 12'b010000000000;
		14'b01000000101110: color_data = 12'b010000000000;
		14'b01000000101111: color_data = 12'b010000000000;
		14'b01000000110000: color_data = 12'b010000000000;
		14'b01000000110001: color_data = 12'b001000000000;
		14'b01000001010010: color_data = 12'b001000000000;
		14'b01000001010011: color_data = 12'b001000000000;
		14'b01000001010100: color_data = 12'b001000000000;
		14'b01000001010101: color_data = 12'b001000000000;
		14'b01000001010110: color_data = 12'b001000000000;
		14'b01000001010111: color_data = 12'b001000000000;
		14'b01000001011000: color_data = 12'b010000000000;
		14'b01000001011001: color_data = 12'b010000000000;
		14'b01000001011010: color_data = 12'b010000000000;
		14'b01000001011011: color_data = 12'b010000000000;
		14'b01000001011100: color_data = 12'b001000000000;
		14'b01000001011101: color_data = 12'b001000000000;
		14'b01000001011110: color_data = 12'b001000000000;
		14'b01000001011111: color_data = 12'b010000000000;
		14'b01000001100000: color_data = 12'b010000000000;
		14'b01000001100001: color_data = 12'b010000000000;
		14'b01000001100010: color_data = 12'b010000000000;
		14'b01000001100011: color_data = 12'b010000000000;
		14'b01000001100100: color_data = 12'b001000000000;
		14'b01000001100101: color_data = 12'b001000000000;
		14'b01000001100110: color_data = 12'b001000000000;
		14'b01000001100111: color_data = 12'b001000000000;
		14'b01000001111000: color_data = 12'b001000000000;
		14'b01000001111001: color_data = 12'b001000000000;
		14'b01000001111010: color_data = 12'b001000000000;
		14'b01000001111011: color_data = 12'b001000000000;
		14'b01000010001010: color_data = 12'b001000000000;
		14'b01000010001011: color_data = 12'b001000000000;
		14'b01000010001100: color_data = 12'b001000000000;
		14'b01000010100110: color_data = 12'b001000000000;
		14'b01000010100111: color_data = 12'b001000000000;
		14'b01000010101000: color_data = 12'b010000000000;
		14'b01000010101001: color_data = 12'b010000000000;
		14'b01000010101010: color_data = 12'b010000000000;
		14'b01000010101011: color_data = 12'b010000000000;
		14'b01000010101100: color_data = 12'b010000000000;
		14'b01000010101101: color_data = 12'b010000000000;
		14'b01000010101110: color_data = 12'b010000000000;
		14'b01000010101111: color_data = 12'b001000000000;
		14'b01000010110000: color_data = 12'b001000000000;
		14'b01000011010001: color_data = 12'b001000000000;
		14'b01000011010010: color_data = 12'b001000000000;
		14'b01000011010011: color_data = 12'b001000000000;
		14'b01000011010100: color_data = 12'b001000000000;
		14'b01000011010101: color_data = 12'b010000000000;
		14'b01000011010110: color_data = 12'b010000000000;
		14'b01000011010111: color_data = 12'b010000000000;
		14'b01000011011000: color_data = 12'b010000000000;
		14'b01000011011001: color_data = 12'b010000000000;
		14'b01000011011010: color_data = 12'b010000000000;
		14'b01000011011011: color_data = 12'b010000000000;
		14'b01000011011100: color_data = 12'b001000000000;
		14'b01000011011101: color_data = 12'b001000000000;
		14'b01000011011110: color_data = 12'b001000000000;
		14'b01000011011111: color_data = 12'b001000000000;
		14'b01000011100000: color_data = 12'b010000000000;
		14'b01000011100001: color_data = 12'b010000000000;
		14'b01000011100010: color_data = 12'b010000000000;
		14'b01000011100011: color_data = 12'b010000000000;
		14'b01000011100100: color_data = 12'b001000000000;
		14'b01000011100101: color_data = 12'b001000000000;
		14'b01000011100110: color_data = 12'b001000000000;
		14'b01000011100111: color_data = 12'b001000000000;
		14'b01000011111000: color_data = 12'b001000000000;
		14'b01000011111001: color_data = 12'b001000000000;
		14'b01000011111010: color_data = 12'b001000000000;
		14'b01000011111011: color_data = 12'b001000000000;
		14'b01000100001011: color_data = 12'b001000000000;
		14'b01000100001100: color_data = 12'b001000000000;
		14'b01000100100101: color_data = 12'b001000000000;
		14'b01000100100110: color_data = 12'b001000000000;
		14'b01000100100111: color_data = 12'b010000000000;
		14'b01000100101000: color_data = 12'b010000000000;
		14'b01000100101001: color_data = 12'b010000000000;
		14'b01000100101010: color_data = 12'b010000000000;
		14'b01000100101011: color_data = 12'b010000000000;
		14'b01000100101100: color_data = 12'b010000000000;
		14'b01000100101101: color_data = 12'b010000000000;
		14'b01000100101110: color_data = 12'b001000000000;
		14'b01000101010000: color_data = 12'b001000000000;
		14'b01000101010001: color_data = 12'b001000000000;
		14'b01000101010010: color_data = 12'b010000000000;
		14'b01000101010011: color_data = 12'b010000000000;
		14'b01000101010100: color_data = 12'b010000000000;
		14'b01000101010101: color_data = 12'b010000000000;
		14'b01000101010110: color_data = 12'b010000000000;
		14'b01000101010111: color_data = 12'b010000000000;
		14'b01000101011000: color_data = 12'b010000000000;
		14'b01000101011001: color_data = 12'b010000000000;
		14'b01000101011010: color_data = 12'b010000000000;
		14'b01000101011011: color_data = 12'b010000000000;
		14'b01000101011100: color_data = 12'b010000000000;
		14'b01000101011101: color_data = 12'b001000000000;
		14'b01000101011110: color_data = 12'b001000000000;
		14'b01000101011111: color_data = 12'b001000000000;
		14'b01000101100000: color_data = 12'b001000000000;
		14'b01000101100001: color_data = 12'b010000000000;
		14'b01000101100010: color_data = 12'b010000000000;
		14'b01000101100011: color_data = 12'b010000000000;
		14'b01000101100100: color_data = 12'b010000000000;
		14'b01000101100101: color_data = 12'b001000000000;
		14'b01000101100110: color_data = 12'b001000000000;
		14'b01000101100111: color_data = 12'b001000000000;
		14'b01000101101000: color_data = 12'b001000000000;
		14'b01000101111010: color_data = 12'b001000000000;
		14'b01000101111011: color_data = 12'b001000000000;
		14'b01000110001011: color_data = 12'b001000000000;
		14'b01000110001100: color_data = 12'b001000000000;
		14'b01000110100011: color_data = 12'b001000000000;
		14'b01000110100100: color_data = 12'b001000000000;
		14'b01000110100101: color_data = 12'b001000000000;
		14'b01000110100110: color_data = 12'b010000000000;
		14'b01000110100111: color_data = 12'b010000000000;
		14'b01000110101000: color_data = 12'b010000000000;
		14'b01000110101001: color_data = 12'b010000000000;
		14'b01000110101010: color_data = 12'b010000000000;
		14'b01000110101011: color_data = 12'b001000000000;
		14'b01000110101100: color_data = 12'b001000000000;
		14'b01000110101101: color_data = 12'b001000000000;
		14'b01000111010000: color_data = 12'b010000000000;
		14'b01000111010001: color_data = 12'b010000000000;
		14'b01000111010010: color_data = 12'b010000000000;
		14'b01000111010011: color_data = 12'b010000000000;
		14'b01000111010100: color_data = 12'b010000000000;
		14'b01000111010101: color_data = 12'b010000000000;
		14'b01000111010110: color_data = 12'b010000000000;
		14'b01000111010111: color_data = 12'b010000000000;
		14'b01000111011000: color_data = 12'b010000000000;
		14'b01000111011001: color_data = 12'b010000000000;
		14'b01000111011010: color_data = 12'b010000000000;
		14'b01000111011011: color_data = 12'b010000000000;
		14'b01000111011100: color_data = 12'b010000000000;
		14'b01000111011101: color_data = 12'b010000000000;
		14'b01000111011110: color_data = 12'b001000000000;
		14'b01000111011111: color_data = 12'b001000000000;
		14'b01000111100000: color_data = 12'b001000000000;
		14'b01000111100001: color_data = 12'b001000000000;
		14'b01000111100010: color_data = 12'b010000000000;
		14'b01000111100011: color_data = 12'b010000000000;
		14'b01000111100100: color_data = 12'b010000000000;
		14'b01000111100101: color_data = 12'b010000000000;
		14'b01000111100110: color_data = 12'b001000000000;
		14'b01000111100111: color_data = 12'b001000000000;
		14'b01000111101000: color_data = 12'b001000000000;
		14'b01000111111010: color_data = 12'b001000000000;
		14'b01000111111011: color_data = 12'b001000000000;
		14'b01000111111100: color_data = 12'b001000000000;
		14'b01001000001100: color_data = 12'b001000000000;
		14'b01001000100011: color_data = 12'b001000000000;
		14'b01001000100100: color_data = 12'b001000000000;
		14'b01001000100101: color_data = 12'b001000000000;
		14'b01001000100110: color_data = 12'b001000000000;
		14'b01001000100111: color_data = 12'b001000000000;
		14'b01001000101000: color_data = 12'b001000000000;
		14'b01001000101001: color_data = 12'b001000000000;
		14'b01001000101010: color_data = 12'b001000000000;
		14'b01001000101011: color_data = 12'b001000000000;
		14'b01001000101100: color_data = 12'b001000000000;
		14'b01001001001110: color_data = 12'b010000000000;
		14'b01001001001111: color_data = 12'b010000000000;
		14'b01001001010000: color_data = 12'b010000000000;
		14'b01001001010001: color_data = 12'b010000000000;
		14'b01001001010010: color_data = 12'b010000000000;
		14'b01001001010011: color_data = 12'b010000000000;
		14'b01001001010100: color_data = 12'b010000000000;
		14'b01001001010101: color_data = 12'b010000000000;
		14'b01001001010110: color_data = 12'b010000000000;
		14'b01001001010111: color_data = 12'b010000000000;
		14'b01001001011000: color_data = 12'b010000000000;
		14'b01001001011001: color_data = 12'b010000000000;
		14'b01001001011010: color_data = 12'b010000000000;
		14'b01001001011011: color_data = 12'b010000000000;
		14'b01001001011100: color_data = 12'b010000000000;
		14'b01001001011101: color_data = 12'b010000000000;
		14'b01001001011110: color_data = 12'b001000000000;
		14'b01001001011111: color_data = 12'b001000000000;
		14'b01001001100000: color_data = 12'b001000000000;
		14'b01001001100001: color_data = 12'b001000000000;
		14'b01001001100010: color_data = 12'b001000000000;
		14'b01001001100011: color_data = 12'b010000000000;
		14'b01001001100100: color_data = 12'b010000000000;
		14'b01001001100101: color_data = 12'b010000000000;
		14'b01001001100110: color_data = 12'b010000000000;
		14'b01001001100111: color_data = 12'b001000000000;
		14'b01001001101000: color_data = 12'b001000000000;
		14'b01001001111011: color_data = 12'b001000000000;
		14'b01001010001101: color_data = 12'b001000000000;
		14'b01001010100010: color_data = 12'b001000000000;
		14'b01001010100011: color_data = 12'b001000000000;
		14'b01001010100100: color_data = 12'b001000000000;
		14'b01001010100101: color_data = 12'b001000000000;
		14'b01001010100110: color_data = 12'b001000000000;
		14'b01001010100111: color_data = 12'b001000000000;
		14'b01001010101000: color_data = 12'b001000000000;
		14'b01001010101001: color_data = 12'b001000000000;
		14'b01001010101010: color_data = 12'b001000000000;
		14'b01001011001101: color_data = 12'b010000000000;
		14'b01001011001110: color_data = 12'b010000000000;
		14'b01001011001111: color_data = 12'b010000000000;
		14'b01001011010000: color_data = 12'b010000000000;
		14'b01001011010001: color_data = 12'b010000000000;
		14'b01001011010010: color_data = 12'b010000000000;
		14'b01001011010011: color_data = 12'b010000000000;
		14'b01001011010100: color_data = 12'b010000000000;
		14'b01001011010101: color_data = 12'b010000000000;
		14'b01001011010110: color_data = 12'b010000000000;
		14'b01001011010111: color_data = 12'b010000000000;
		14'b01001011011000: color_data = 12'b010000000000;
		14'b01001011011001: color_data = 12'b010000000000;
		14'b01001011011010: color_data = 12'b010000000000;
		14'b01001011011011: color_data = 12'b010000000000;
		14'b01001011011100: color_data = 12'b010000000000;
		14'b01001011011101: color_data = 12'b010000000000;
		14'b01001011011110: color_data = 12'b010000000000;
		14'b01001011011111: color_data = 12'b001000000000;
		14'b01001011100000: color_data = 12'b001000000000;
		14'b01001011100001: color_data = 12'b001000000000;
		14'b01001011100010: color_data = 12'b001000000000;
		14'b01001011100011: color_data = 12'b001000000000;
		14'b01001011100100: color_data = 12'b001000000000;
		14'b01001011100101: color_data = 12'b001000000000;
		14'b01001011100110: color_data = 12'b001000000000;
		14'b01001011100111: color_data = 12'b001000000000;
		14'b01001011101000: color_data = 12'b001000000000;
		14'b01001100001110: color_data = 12'b001000000000;
		14'b01001100100001: color_data = 12'b001000000000;
		14'b01001100100010: color_data = 12'b001000000000;
		14'b01001100100011: color_data = 12'b001000000000;
		14'b01001100100100: color_data = 12'b001000000000;
		14'b01001100100101: color_data = 12'b001000000000;
		14'b01001100100110: color_data = 12'b001000000000;
		14'b01001100100111: color_data = 12'b001000000000;
		14'b01001101001011: color_data = 12'b001000000000;
		14'b01001101001100: color_data = 12'b010000000000;
		14'b01001101001101: color_data = 12'b010000000000;
		14'b01001101001110: color_data = 12'b010000000000;
		14'b01001101001111: color_data = 12'b010000000000;
		14'b01001101010000: color_data = 12'b010000000000;
		14'b01001101010001: color_data = 12'b010000000000;
		14'b01001101010010: color_data = 12'b010000000000;
		14'b01001101010011: color_data = 12'b010000000000;
		14'b01001101010100: color_data = 12'b010000000000;
		14'b01001101010101: color_data = 12'b010000000000;
		14'b01001101010110: color_data = 12'b010000000000;
		14'b01001101010111: color_data = 12'b010000000000;
		14'b01001101011000: color_data = 12'b010000000000;
		14'b01001101011001: color_data = 12'b010000000000;
		14'b01001101011010: color_data = 12'b010000000000;
		14'b01001101011011: color_data = 12'b010000000000;
		14'b01001101011100: color_data = 12'b010000000000;
		14'b01001101011101: color_data = 12'b010000000000;
		14'b01001101011110: color_data = 12'b010000000000;
		14'b01001101011111: color_data = 12'b010000000000;
		14'b01001101100000: color_data = 12'b001000000000;
		14'b01001101100011: color_data = 12'b001000000000;
		14'b01001101100100: color_data = 12'b001000000000;
		14'b01001101100101: color_data = 12'b001000000000;
		14'b01001101100110: color_data = 12'b001000000000;
		14'b01001101100111: color_data = 12'b001000000000;
		14'b01001101101000: color_data = 12'b001000000000;
		14'b01001110100001: color_data = 12'b001000000000;
		14'b01001110100010: color_data = 12'b001000000000;
		14'b01001110100011: color_data = 12'b001000000000;
		14'b01001110100100: color_data = 12'b001000000000;
		14'b01001110100101: color_data = 12'b001000000000;
		14'b01001111001010: color_data = 12'b010000000000;
		14'b01001111001011: color_data = 12'b010000000000;
		14'b01001111001100: color_data = 12'b010000000000;
		14'b01001111001101: color_data = 12'b010000000000;
		14'b01001111001110: color_data = 12'b010000000000;
		14'b01001111001111: color_data = 12'b010000000000;
		14'b01001111010000: color_data = 12'b010000000000;
		14'b01001111010001: color_data = 12'b010000000000;
		14'b01001111010010: color_data = 12'b010000000000;
		14'b01001111010011: color_data = 12'b010000000000;
		14'b01001111010100: color_data = 12'b010000000000;
		14'b01001111010101: color_data = 12'b010000000000;
		14'b01001111010110: color_data = 12'b010000000000;
		14'b01001111010111: color_data = 12'b010000000000;
		14'b01001111011000: color_data = 12'b010000000000;
		14'b01001111011001: color_data = 12'b010000000000;
		14'b01001111011010: color_data = 12'b010000000000;
		14'b01001111011011: color_data = 12'b010000000000;
		14'b01001111011100: color_data = 12'b010000000000;
		14'b01001111011101: color_data = 12'b010000000000;
		14'b01001111011110: color_data = 12'b010000000000;
		14'b01001111011111: color_data = 12'b010000000000;
		14'b01001111100000: color_data = 12'b001000000000;
		14'b01001111100101: color_data = 12'b001000000000;
		14'b01001111100110: color_data = 12'b001000000000;
		14'b01001111100111: color_data = 12'b001000000000;
		14'b01001111101000: color_data = 12'b001000000000;
		14'b01001111101001: color_data = 12'b001000000000;
		14'b01010000100001: color_data = 12'b001000000000;
		14'b01010000100010: color_data = 12'b001000000000;
		14'b01010001000111: color_data = 12'b010000000000;
		14'b01010001001000: color_data = 12'b010000000000;
		14'b01010001001001: color_data = 12'b010000000000;
		14'b01010001001010: color_data = 12'b010000000000;
		14'b01010001001011: color_data = 12'b010000000000;
		14'b01010001001100: color_data = 12'b010000000000;
		14'b01010001001101: color_data = 12'b010000000000;
		14'b01010001001110: color_data = 12'b010000000000;
		14'b01010001001111: color_data = 12'b010000000000;
		14'b01010001010000: color_data = 12'b010000000000;
		14'b01010001010001: color_data = 12'b010000000000;
		14'b01010001010010: color_data = 12'b010000000000;
		14'b01010001010011: color_data = 12'b010000000000;
		14'b01010001010100: color_data = 12'b010000000000;
		14'b01010001010101: color_data = 12'b010000000000;
		14'b01010001010110: color_data = 12'b010000000000;
		14'b01010001010111: color_data = 12'b010000000000;
		14'b01010001011000: color_data = 12'b010000000000;
		14'b01010001011001: color_data = 12'b010000000000;
		14'b01010001011010: color_data = 12'b010000000000;
		14'b01010001011011: color_data = 12'b010000000000;
		14'b01010001011100: color_data = 12'b010000000000;
		14'b01010001011101: color_data = 12'b010000000000;
		14'b01010001011110: color_data = 12'b010000000000;
		14'b01010001011111: color_data = 12'b010000000000;
		14'b01010001100000: color_data = 12'b001000000000;
		14'b01010001100111: color_data = 12'b001000000000;
		14'b01010001101000: color_data = 12'b001000000000;
		14'b01010001101001: color_data = 12'b001000000000;
		14'b01010010100010: color_data = 12'b001000000000;
		14'b01010011000101: color_data = 12'b001000000000;
		14'b01010011000110: color_data = 12'b001000000000;
		14'b01010011000111: color_data = 12'b010000000000;
		14'b01010011001000: color_data = 12'b010000000000;
		14'b01010011001001: color_data = 12'b010000000000;
		14'b01010011001010: color_data = 12'b010000000000;
		14'b01010011001011: color_data = 12'b010000000000;
		14'b01010011001100: color_data = 12'b010000000000;
		14'b01010011001101: color_data = 12'b010000000000;
		14'b01010011001110: color_data = 12'b010000000000;
		14'b01010011001111: color_data = 12'b010000000000;
		14'b01010011010000: color_data = 12'b010000000000;
		14'b01010011010001: color_data = 12'b010000000000;
		14'b01010011010010: color_data = 12'b010000000000;
		14'b01010011010011: color_data = 12'b010000000000;
		14'b01010011010100: color_data = 12'b010000000000;
		14'b01010011010101: color_data = 12'b010000000000;
		14'b01010011010110: color_data = 12'b010000000000;
		14'b01010011010111: color_data = 12'b010000000000;
		14'b01010011011000: color_data = 12'b010000000000;
		14'b01010011011001: color_data = 12'b010000000000;
		14'b01010011011010: color_data = 12'b010000000000;
		14'b01010011011011: color_data = 12'b010000000000;
		14'b01010011011100: color_data = 12'b010000000000;
		14'b01010011011101: color_data = 12'b010000000000;
		14'b01010011011110: color_data = 12'b010000000000;
		14'b01010011011111: color_data = 12'b010000000000;
		14'b01010011100000: color_data = 12'b010000000000;
		14'b01010011100001: color_data = 12'b001000000000;
		14'b01010011101001: color_data = 12'b001000000000;
		14'b01010011101010: color_data = 12'b001000000000;
		14'b01010100100011: color_data = 12'b001000000000;
		14'b01010101000011: color_data = 12'b001000000000;
		14'b01010101000100: color_data = 12'b001000000000;
		14'b01010101000101: color_data = 12'b010000000000;
		14'b01010101000110: color_data = 12'b010000000000;
		14'b01010101000111: color_data = 12'b010000000000;
		14'b01010101001000: color_data = 12'b010000000000;
		14'b01010101001001: color_data = 12'b010000000000;
		14'b01010101001010: color_data = 12'b010000000000;
		14'b01010101001011: color_data = 12'b010000000000;
		14'b01010101001100: color_data = 12'b010000000000;
		14'b01010101001101: color_data = 12'b010000000000;
		14'b01010101001110: color_data = 12'b010000000000;
		14'b01010101001111: color_data = 12'b010000000000;
		14'b01010101010000: color_data = 12'b010000000000;
		14'b01010101010001: color_data = 12'b010000000000;
		14'b01010101010010: color_data = 12'b010000000000;
		14'b01010101010011: color_data = 12'b010000000000;
		14'b01010101010100: color_data = 12'b010000000000;
		14'b01010101010101: color_data = 12'b010000000000;
		14'b01010101010110: color_data = 12'b010000000000;
		14'b01010101010111: color_data = 12'b010000000000;
		14'b01010101011000: color_data = 12'b010000000000;
		14'b01010101011001: color_data = 12'b010000000000;
		14'b01010101011010: color_data = 12'b010000000000;
		14'b01010101011011: color_data = 12'b010000000000;
		14'b01010101011100: color_data = 12'b010000000000;
		14'b01010101011101: color_data = 12'b010000000000;
		14'b01010101011110: color_data = 12'b010000000000;
		14'b01010101011111: color_data = 12'b010000000000;
		14'b01010101100000: color_data = 12'b010000000000;
		14'b01010101100001: color_data = 12'b010000000000;
		14'b01010101100010: color_data = 12'b001000000000;
		14'b01010101100011: color_data = 12'b001000000000;
		14'b01010111000001: color_data = 12'b001000000000;
		14'b01010111000010: color_data = 12'b001000000000;
		14'b01010111000011: color_data = 12'b010000000000;
		14'b01010111000100: color_data = 12'b010000000000;
		14'b01010111000101: color_data = 12'b010000000000;
		14'b01010111000110: color_data = 12'b010000000000;
		14'b01010111000111: color_data = 12'b010000000000;
		14'b01010111001000: color_data = 12'b010000000000;
		14'b01010111001001: color_data = 12'b010000000000;
		14'b01010111001010: color_data = 12'b010000000000;
		14'b01010111001011: color_data = 12'b010000000000;
		14'b01010111001100: color_data = 12'b010000000000;
		14'b01010111001101: color_data = 12'b010000000000;
		14'b01010111001110: color_data = 12'b010000000000;
		14'b01010111001111: color_data = 12'b010000000000;
		14'b01010111010000: color_data = 12'b010000000000;
		14'b01010111010001: color_data = 12'b010000000000;
		14'b01010111010010: color_data = 12'b010000000000;
		14'b01010111010011: color_data = 12'b010000000000;
		14'b01010111010100: color_data = 12'b010000000000;
		14'b01010111010101: color_data = 12'b010000000000;
		14'b01010111010110: color_data = 12'b010000000000;
		14'b01010111010111: color_data = 12'b010000000000;
		14'b01010111011000: color_data = 12'b010000000000;
		14'b01010111011001: color_data = 12'b010000000000;
		14'b01010111011010: color_data = 12'b010000000000;
		14'b01010111011011: color_data = 12'b001000000000;
		14'b01010111011100: color_data = 12'b001000000000;
		14'b01010111011101: color_data = 12'b001000000000;
		14'b01010111011110: color_data = 12'b010000000000;
		14'b01010111011111: color_data = 12'b010000000000;
		14'b01010111100000: color_data = 12'b010000000000;
		14'b01010111100001: color_data = 12'b010000000000;
		14'b01010111100010: color_data = 12'b010000000000;
		14'b01010111100011: color_data = 12'b001000000000;
		14'b01010111100100: color_data = 12'b001000000000;
		14'b01011000111110: color_data = 12'b001000000000;
		14'b01011000111111: color_data = 12'b001000000000;
		14'b01011001000000: color_data = 12'b001000000000;
		14'b01011001000001: color_data = 12'b001000000000;
		14'b01011001000010: color_data = 12'b010000000000;
		14'b01011001000011: color_data = 12'b010000000000;
		14'b01011001000100: color_data = 12'b010000000000;
		14'b01011001000101: color_data = 12'b010000000000;
		14'b01011001000110: color_data = 12'b010000000000;
		14'b01011001000111: color_data = 12'b010000000000;
		14'b01011001001000: color_data = 12'b010000000000;
		14'b01011001001001: color_data = 12'b010000000000;
		14'b01011001001010: color_data = 12'b010000000000;
		14'b01011001001011: color_data = 12'b010000000000;
		14'b01011001001100: color_data = 12'b010000000000;
		14'b01011001001101: color_data = 12'b010000000000;
		14'b01011001001110: color_data = 12'b010000000000;
		14'b01011001001111: color_data = 12'b010000000000;
		14'b01011001010000: color_data = 12'b010000000000;
		14'b01011001010001: color_data = 12'b010000000000;
		14'b01011001010010: color_data = 12'b010000000000;
		14'b01011001010011: color_data = 12'b010000000000;
		14'b01011001010100: color_data = 12'b010000000000;
		14'b01011001010101: color_data = 12'b010000000000;
		14'b01011001010110: color_data = 12'b010000000000;
		14'b01011001010111: color_data = 12'b010000000000;
		14'b01011001011000: color_data = 12'b010000000000;
		14'b01011001011001: color_data = 12'b010000000000;
		14'b01011001011010: color_data = 12'b010000000000;
		14'b01011001011011: color_data = 12'b010000000000;
		14'b01011001011100: color_data = 12'b001000000000;
		14'b01011001011101: color_data = 12'b001000000000;
		14'b01011001011110: color_data = 12'b001000000000;
		14'b01011001011111: color_data = 12'b001000000000;
		14'b01011001100000: color_data = 12'b010000000000;
		14'b01011001100001: color_data = 12'b010000000000;
		14'b01011001100010: color_data = 12'b010000000000;
		14'b01011001100011: color_data = 12'b010000000000;
		14'b01011001100100: color_data = 12'b001000000000;
		14'b01011001100101: color_data = 12'b001000000000;
		14'b01011010000000: color_data = 12'b001000000000;
		14'b01011010000001: color_data = 12'b001000000000;
		14'b01011010000010: color_data = 12'b001000000000;
		14'b01011010010101: color_data = 12'b001000000000;
		14'b01011010010110: color_data = 12'b001000000000;
		14'b01011010010111: color_data = 12'b001000000000;
		14'b01011010110010: color_data = 12'b001000000000;
		14'b01011010110011: color_data = 12'b001000000000;
		14'b01011010110100: color_data = 12'b001000000000;
		14'b01011010111010: color_data = 12'b001000000000;
		14'b01011010111011: color_data = 12'b001000000000;
		14'b01011010111100: color_data = 12'b001000000000;
		14'b01011010111101: color_data = 12'b001000000000;
		14'b01011010111110: color_data = 12'b001000000000;
		14'b01011010111111: color_data = 12'b001000000000;
		14'b01011011000000: color_data = 12'b010000000000;
		14'b01011011000001: color_data = 12'b010000000000;
		14'b01011011000010: color_data = 12'b010000000000;
		14'b01011011000011: color_data = 12'b010000000000;
		14'b01011011000100: color_data = 12'b010000000000;
		14'b01011011000101: color_data = 12'b010000000000;
		14'b01011011000110: color_data = 12'b010000000000;
		14'b01011011000111: color_data = 12'b010000000000;
		14'b01011011001000: color_data = 12'b010000000000;
		14'b01011011001001: color_data = 12'b010000000000;
		14'b01011011001010: color_data = 12'b010000000000;
		14'b01011011001011: color_data = 12'b010000000000;
		14'b01011011001100: color_data = 12'b010000000000;
		14'b01011011001101: color_data = 12'b010000000000;
		14'b01011011001110: color_data = 12'b010000000000;
		14'b01011011001111: color_data = 12'b010000000000;
		14'b01011011010000: color_data = 12'b010000000000;
		14'b01011011010001: color_data = 12'b010000000000;
		14'b01011011010010: color_data = 12'b010000000000;
		14'b01011011010011: color_data = 12'b010000000000;
		14'b01011011010100: color_data = 12'b010000000000;
		14'b01011011010101: color_data = 12'b010000000000;
		14'b01011011010110: color_data = 12'b010000000000;
		14'b01011011010111: color_data = 12'b010000000000;
		14'b01011011011000: color_data = 12'b010000000000;
		14'b01011011011001: color_data = 12'b010000000000;
		14'b01011011011010: color_data = 12'b010000000000;
		14'b01011011011011: color_data = 12'b010000000000;
		14'b01011011011100: color_data = 12'b010000000000;
		14'b01011011011101: color_data = 12'b010000000000;
		14'b01011011011110: color_data = 12'b010000000000;
		14'b01011011011111: color_data = 12'b001000000000;
		14'b01011011100000: color_data = 12'b001000000000;
		14'b01011011100001: color_data = 12'b010000000000;
		14'b01011011100010: color_data = 12'b010000000000;
		14'b01011011100011: color_data = 12'b010000000000;
		14'b01011011100100: color_data = 12'b010000000000;
		14'b01011011100101: color_data = 12'b010000000000;
		14'b01011011100110: color_data = 12'b001000000000;
		14'b01011100000000: color_data = 12'b001000000000;
		14'b01011100000001: color_data = 12'b001000000000;
		14'b01011100000010: color_data = 12'b010000000000;
		14'b01011100000011: color_data = 12'b010000000000;
		14'b01011100000100: color_data = 12'b001000000000;
		14'b01011100000101: color_data = 12'b001000000000;
		14'b01011100000110: color_data = 12'b001000000000;
		14'b01011100010101: color_data = 12'b001000000000;
		14'b01011100010110: color_data = 12'b010000000000;
		14'b01011100010111: color_data = 12'b010000000000;
		14'b01011100011000: color_data = 12'b010000000000;
		14'b01011100011001: color_data = 12'b001000000000;
		14'b01011100011010: color_data = 12'b001000000000;
		14'b01011100011011: color_data = 12'b001000000000;
		14'b01011100101101: color_data = 12'b001000000000;
		14'b01011100101110: color_data = 12'b001000000000;
		14'b01011100101111: color_data = 12'b001000000000;
		14'b01011100110000: color_data = 12'b001000000000;
		14'b01011100110001: color_data = 12'b001000000000;
		14'b01011100110010: color_data = 12'b001000000000;
		14'b01011100110011: color_data = 12'b001000000000;
		14'b01011100110100: color_data = 12'b001000000000;
		14'b01011100110101: color_data = 12'b001000000000;
		14'b01011100110110: color_data = 12'b001000000000;
		14'b01011100110111: color_data = 12'b001000000000;
		14'b01011100111000: color_data = 12'b001000000000;
		14'b01011100111001: color_data = 12'b001000000000;
		14'b01011100111010: color_data = 12'b001000000000;
		14'b01011100111011: color_data = 12'b001000000000;
		14'b01011100111100: color_data = 12'b010000000000;
		14'b01011100111101: color_data = 12'b010000000000;
		14'b01011100111110: color_data = 12'b010000000000;
		14'b01011100111111: color_data = 12'b010000000000;
		14'b01011101000000: color_data = 12'b010000000000;
		14'b01011101000001: color_data = 12'b010000000000;
		14'b01011101000010: color_data = 12'b010000000000;
		14'b01011101000011: color_data = 12'b010000000000;
		14'b01011101000100: color_data = 12'b010000000000;
		14'b01011101000101: color_data = 12'b010000000000;
		14'b01011101000110: color_data = 12'b010000000000;
		14'b01011101000111: color_data = 12'b010000000000;
		14'b01011101001000: color_data = 12'b010000000000;
		14'b01011101001001: color_data = 12'b010000000000;
		14'b01011101001010: color_data = 12'b010000000000;
		14'b01011101001011: color_data = 12'b001000000000;
		14'b01011101001100: color_data = 12'b001000000000;
		14'b01011101001101: color_data = 12'b001000000000;
		14'b01011101001110: color_data = 12'b001000000000;
		14'b01011101001111: color_data = 12'b001000000000;
		14'b01011101010000: color_data = 12'b001000000000;
		14'b01011101010001: color_data = 12'b001000000000;
		14'b01011101010010: color_data = 12'b010000000000;
		14'b01011101010011: color_data = 12'b010000000000;
		14'b01011101010100: color_data = 12'b010000000000;
		14'b01011101010101: color_data = 12'b010000000000;
		14'b01011101010110: color_data = 12'b010000000000;
		14'b01011101010111: color_data = 12'b010000000000;
		14'b01011101011000: color_data = 12'b010000000000;
		14'b01011101011001: color_data = 12'b001000000000;
		14'b01011101011010: color_data = 12'b010000000000;
		14'b01011101011011: color_data = 12'b010000000000;
		14'b01011101011100: color_data = 12'b010000000000;
		14'b01011101011101: color_data = 12'b010000000000;
		14'b01011101011110: color_data = 12'b010000000000;
		14'b01011101011111: color_data = 12'b010000000000;
		14'b01011101100000: color_data = 12'b010000000000;
		14'b01011101100001: color_data = 12'b001000000000;
		14'b01011101100010: color_data = 12'b001000000000;
		14'b01011101100011: color_data = 12'b010000000000;
		14'b01011101100100: color_data = 12'b010000000000;
		14'b01011101100101: color_data = 12'b010000000000;
		14'b01011101100110: color_data = 12'b010000000000;
		14'b01011101100111: color_data = 12'b001000000000;
		14'b01011101111111: color_data = 12'b001000000000;
		14'b01011110000011: color_data = 12'b001000000000;
		14'b01011110000100: color_data = 12'b010000000000;
		14'b01011110000101: color_data = 12'b010000000000;
		14'b01011110000110: color_data = 12'b010000000000;
		14'b01011110000111: color_data = 12'b010000000000;
		14'b01011110001000: color_data = 12'b001000000000;
		14'b01011110001001: color_data = 12'b001000000000;
		14'b01011110010000: color_data = 12'b001000000000;
		14'b01011110010110: color_data = 12'b001000000000;
		14'b01011110010111: color_data = 12'b010000000000;
		14'b01011110011000: color_data = 12'b010000000000;
		14'b01011110011001: color_data = 12'b010000000000;
		14'b01011110011010: color_data = 12'b010000000000;
		14'b01011110011011: color_data = 12'b010000000000;
		14'b01011110011100: color_data = 12'b010000000000;
		14'b01011110011101: color_data = 12'b010000000000;
		14'b01011110011110: color_data = 12'b001000000000;
		14'b01011110011111: color_data = 12'b010000000000;
		14'b01011110100000: color_data = 12'b010000000000;
		14'b01011110100001: color_data = 12'b010000000000;
		14'b01011110100010: color_data = 12'b010000000000;
		14'b01011110100011: color_data = 12'b010000000000;
		14'b01011110100100: color_data = 12'b001000000000;
		14'b01011110100101: color_data = 12'b001000000000;
		14'b01011110100110: color_data = 12'b001000000000;
		14'b01011110100111: color_data = 12'b001000000000;
		14'b01011110101000: color_data = 12'b001000000000;
		14'b01011110101001: color_data = 12'b001000000000;
		14'b01011110101010: color_data = 12'b001000000000;
		14'b01011110101011: color_data = 12'b001000000000;
		14'b01011110101100: color_data = 12'b001000000000;
		14'b01011110101101: color_data = 12'b001000000000;
		14'b01011110101110: color_data = 12'b001000000000;
		14'b01011110101111: color_data = 12'b001000000000;
		14'b01011110110000: color_data = 12'b001000000000;
		14'b01011110110001: color_data = 12'b001000000000;
		14'b01011110110010: color_data = 12'b001000000000;
		14'b01011110110011: color_data = 12'b001000000000;
		14'b01011110110100: color_data = 12'b001000000000;
		14'b01011110110101: color_data = 12'b001000000000;
		14'b01011110110110: color_data = 12'b001000000000;
		14'b01011110110111: color_data = 12'b001000000000;
		14'b01011110111000: color_data = 12'b010000000000;
		14'b01011110111001: color_data = 12'b010000000000;
		14'b01011110111010: color_data = 12'b010000000000;
		14'b01011110111011: color_data = 12'b010000000000;
		14'b01011110111100: color_data = 12'b010000000000;
		14'b01011110111101: color_data = 12'b010000000000;
		14'b01011110111110: color_data = 12'b010000000000;
		14'b01011110111111: color_data = 12'b010000000000;
		14'b01011111000000: color_data = 12'b010000000000;
		14'b01011111000001: color_data = 12'b010000000000;
		14'b01011111000010: color_data = 12'b010000000000;
		14'b01011111000011: color_data = 12'b010000000000;
		14'b01011111000100: color_data = 12'b010000000000;
		14'b01011111000101: color_data = 12'b010000000000;
		14'b01011111000110: color_data = 12'b010000000000;
		14'b01011111000111: color_data = 12'b010000000000;
		14'b01011111001000: color_data = 12'b001000000000;
		14'b01011111001001: color_data = 12'b001000000000;
		14'b01011111001010: color_data = 12'b001000000000;
		14'b01011111001011: color_data = 12'b001000000000;
		14'b01011111001100: color_data = 12'b001000000000;
		14'b01011111001101: color_data = 12'b001000000000;
		14'b01011111001110: color_data = 12'b001000000000;
		14'b01011111001111: color_data = 12'b001000000000;
		14'b01011111010000: color_data = 12'b001000000000;
		14'b01011111010001: color_data = 12'b001000000000;
		14'b01011111010010: color_data = 12'b001000000000;
		14'b01011111010011: color_data = 12'b001000000000;
		14'b01011111010100: color_data = 12'b001000000000;
		14'b01011111010101: color_data = 12'b010000000000;
		14'b01011111010110: color_data = 12'b010000000000;
		14'b01011111010111: color_data = 12'b001000000000;
		14'b01011111011000: color_data = 12'b001000000000;
		14'b01011111011001: color_data = 12'b001000000000;
		14'b01011111011010: color_data = 12'b001000000000;
		14'b01011111011011: color_data = 12'b001000000000;
		14'b01011111011100: color_data = 12'b001000000000;
		14'b01011111011101: color_data = 12'b010000000000;
		14'b01011111011110: color_data = 12'b010000000000;
		14'b01011111011111: color_data = 12'b010000000000;
		14'b01011111100000: color_data = 12'b010000000000;
		14'b01011111100001: color_data = 12'b010000000000;
		14'b01011111100010: color_data = 12'b001000000000;
		14'b01011111100011: color_data = 12'b001000000000;
		14'b01011111100100: color_data = 12'b010000000000;
		14'b01011111100101: color_data = 12'b010000000000;
		14'b01011111100110: color_data = 12'b010000000000;
		14'b01011111100111: color_data = 12'b010000000000;
		14'b01011111101000: color_data = 12'b010000000000;
		14'b01011111101001: color_data = 12'b001000000000;
		14'b01100000000101: color_data = 12'b001000000000;
		14'b01100000000110: color_data = 12'b001000000000;
		14'b01100000000111: color_data = 12'b010000000000;
		14'b01100000001000: color_data = 12'b010000000000;
		14'b01100000001001: color_data = 12'b010000000000;
		14'b01100000001010: color_data = 12'b010000000000;
		14'b01100000001011: color_data = 12'b010000000000;
		14'b01100000001100: color_data = 12'b001000000000;
		14'b01100000001101: color_data = 12'b001000000000;
		14'b01100000001110: color_data = 12'b001000000000;
		14'b01100000001111: color_data = 12'b001000000000;
		14'b01100000010000: color_data = 12'b001000000000;
		14'b01100000010001: color_data = 12'b001000000000;
		14'b01100000010010: color_data = 12'b010000000000;
		14'b01100000010011: color_data = 12'b001000000000;
		14'b01100000010111: color_data = 12'b001000000000;
		14'b01100000011000: color_data = 12'b010000000000;
		14'b01100000011001: color_data = 12'b010000000000;
		14'b01100000011010: color_data = 12'b010000000000;
		14'b01100000011011: color_data = 12'b010000000000;
		14'b01100000011100: color_data = 12'b010000000000;
		14'b01100000011101: color_data = 12'b010000000000;
		14'b01100000011110: color_data = 12'b010000000000;
		14'b01100000011111: color_data = 12'b001000000000;
		14'b01100000100000: color_data = 12'b001000000000;
		14'b01100000100001: color_data = 12'b010000000000;
		14'b01100000100010: color_data = 12'b010000000000;
		14'b01100000100011: color_data = 12'b010000000000;
		14'b01100000100100: color_data = 12'b010000000000;
		14'b01100000100101: color_data = 12'b010000000000;
		14'b01100000100110: color_data = 12'b010000000000;
		14'b01100000100111: color_data = 12'b010000000000;
		14'b01100000101000: color_data = 12'b010000000000;
		14'b01100000101001: color_data = 12'b001000000000;
		14'b01100000101010: color_data = 12'b001000000000;
		14'b01100000101011: color_data = 12'b001000000000;
		14'b01100000101100: color_data = 12'b001000000000;
		14'b01100000101101: color_data = 12'b001000000000;
		14'b01100000101110: color_data = 12'b001000000000;
		14'b01100000101111: color_data = 12'b001000000000;
		14'b01100000110000: color_data = 12'b001000000000;
		14'b01100000110001: color_data = 12'b001000000000;
		14'b01100000110010: color_data = 12'b001000000000;
		14'b01100000110011: color_data = 12'b001000000000;
		14'b01100000110100: color_data = 12'b001000000000;
		14'b01100000110101: color_data = 12'b010000000000;
		14'b01100000110110: color_data = 12'b010000000000;
		14'b01100000110111: color_data = 12'b010000000000;
		14'b01100000111000: color_data = 12'b010000000000;
		14'b01100000111001: color_data = 12'b010000000000;
		14'b01100000111010: color_data = 12'b010000000000;
		14'b01100000111011: color_data = 12'b010000000000;
		14'b01100000111100: color_data = 12'b010000000000;
		14'b01100000111101: color_data = 12'b010000000000;
		14'b01100000111110: color_data = 12'b010000000000;
		14'b01100000111111: color_data = 12'b010000000000;
		14'b01100001000000: color_data = 12'b010000000000;
		14'b01100001000001: color_data = 12'b010000000000;
		14'b01100001000010: color_data = 12'b010000000000;
		14'b01100001000011: color_data = 12'b010000000000;
		14'b01100001000100: color_data = 12'b010000000000;
		14'b01100001000101: color_data = 12'b010000000000;
		14'b01100001000110: color_data = 12'b010000000000;
		14'b01100001000111: color_data = 12'b001000000000;
		14'b01100001001000: color_data = 12'b001000000000;
		14'b01100001001001: color_data = 12'b001000000000;
		14'b01100001001010: color_data = 12'b001000000000;
		14'b01100001001011: color_data = 12'b001000000000;
		14'b01100001001100: color_data = 12'b001000000000;
		14'b01100001001101: color_data = 12'b001000000000;
		14'b01100001001110: color_data = 12'b001000000000;
		14'b01100001001111: color_data = 12'b001000000000;
		14'b01100001010000: color_data = 12'b001000000000;
		14'b01100001010001: color_data = 12'b001000000000;
		14'b01100001010010: color_data = 12'b001000000000;
		14'b01100001010011: color_data = 12'b001000000000;
		14'b01100001010100: color_data = 12'b001000000000;
		14'b01100001010101: color_data = 12'b001000000000;
		14'b01100001010110: color_data = 12'b001000000000;
		14'b01100001010111: color_data = 12'b001000000000;
		14'b01100001011000: color_data = 12'b001000000000;
		14'b01100001011001: color_data = 12'b001000000000;
		14'b01100001011010: color_data = 12'b001000000000;
		14'b01100001011011: color_data = 12'b001000000000;
		14'b01100001011100: color_data = 12'b001000000000;
		14'b01100001011101: color_data = 12'b001000000000;
		14'b01100001011110: color_data = 12'b001000000000;
		14'b01100001011111: color_data = 12'b001000000000;
		14'b01100001100000: color_data = 12'b010000000000;
		14'b01100001100001: color_data = 12'b010000000000;
		14'b01100001100010: color_data = 12'b010000000000;
		14'b01100001100011: color_data = 12'b010000000000;
		14'b01100001100100: color_data = 12'b001000000000;
		14'b01100001100101: color_data = 12'b010000000000;
		14'b01100001100110: color_data = 12'b010000000000;
		14'b01100001100111: color_data = 12'b010000000000;
		14'b01100001101000: color_data = 12'b010000000000;
		14'b01100001101001: color_data = 12'b010000000000;
		14'b01100001101010: color_data = 12'b001000000000;
		14'b01100010001000: color_data = 12'b001000000000;
		14'b01100010001001: color_data = 12'b001000000000;
		14'b01100010001010: color_data = 12'b001000000000;
		14'b01100010001011: color_data = 12'b010000000000;
		14'b01100010001100: color_data = 12'b010000000000;
		14'b01100010001101: color_data = 12'b010000000000;
		14'b01100010001110: color_data = 12'b010000000000;
		14'b01100010001111: color_data = 12'b010000000000;
		14'b01100010010000: color_data = 12'b010000000000;
		14'b01100010010001: color_data = 12'b010000000000;
		14'b01100010010010: color_data = 12'b010000000000;
		14'b01100010010011: color_data = 12'b010000000000;
		14'b01100010010100: color_data = 12'b001000000000;
		14'b01100010011001: color_data = 12'b001000000000;
		14'b01100010011010: color_data = 12'b001000000000;
		14'b01100010011011: color_data = 12'b010000000000;
		14'b01100010011100: color_data = 12'b010000000000;
		14'b01100010011101: color_data = 12'b010000000000;
		14'b01100010011110: color_data = 12'b010000000000;
		14'b01100010011111: color_data = 12'b001000000000;
		14'b01100010100000: color_data = 12'b001000000000;
		14'b01100010100001: color_data = 12'b001000000000;
		14'b01100010100011: color_data = 12'b001000000000;
		14'b01100010100100: color_data = 12'b001000000000;
		14'b01100010100101: color_data = 12'b001000000000;
		14'b01100010100110: color_data = 12'b010000000000;
		14'b01100010100111: color_data = 12'b010000000000;
		14'b01100010101000: color_data = 12'b010000000000;
		14'b01100010101001: color_data = 12'b010000000000;
		14'b01100010101010: color_data = 12'b010000000000;
		14'b01100010101011: color_data = 12'b010000000000;
		14'b01100010101100: color_data = 12'b010000000000;
		14'b01100010101101: color_data = 12'b010000000000;
		14'b01100010101110: color_data = 12'b010000000000;
		14'b01100010101111: color_data = 12'b001000000000;
		14'b01100010110000: color_data = 12'b001000000000;
		14'b01100010110001: color_data = 12'b001000000000;
		14'b01100010110010: color_data = 12'b001000000000;
		14'b01100010110011: color_data = 12'b001000000000;
		14'b01100010110100: color_data = 12'b001000000000;
		14'b01100010110101: color_data = 12'b010000000000;
		14'b01100010110110: color_data = 12'b010000000000;
		14'b01100010110111: color_data = 12'b010000000000;
		14'b01100010111000: color_data = 12'b010000000000;
		14'b01100010111001: color_data = 12'b010000000000;
		14'b01100010111010: color_data = 12'b010000000000;
		14'b01100010111011: color_data = 12'b010000000000;
		14'b01100010111100: color_data = 12'b010000000000;
		14'b01100010111101: color_data = 12'b010000000000;
		14'b01100010111110: color_data = 12'b010000000000;
		14'b01100010111111: color_data = 12'b010000000000;
		14'b01100011000000: color_data = 12'b010000000000;
		14'b01100011000001: color_data = 12'b010000000000;
		14'b01100011000010: color_data = 12'b001000000000;
		14'b01100011000011: color_data = 12'b001000000000;
		14'b01100011000100: color_data = 12'b001000000000;
		14'b01100011000101: color_data = 12'b010000000000;
		14'b01100011000110: color_data = 12'b001000000000;
		14'b01100011000111: color_data = 12'b001000000000;
		14'b01100011001000: color_data = 12'b001000000000;
		14'b01100011001001: color_data = 12'b001000000000;
		14'b01100011001010: color_data = 12'b001000000000;
		14'b01100011001011: color_data = 12'b001000000000;
		14'b01100011011001: color_data = 12'b001000000000;
		14'b01100011011010: color_data = 12'b001000000000;
		14'b01100011011011: color_data = 12'b001000000000;
		14'b01100011011100: color_data = 12'b001000000000;
		14'b01100011011101: color_data = 12'b001000000000;
		14'b01100011011110: color_data = 12'b001000000000;
		14'b01100011011111: color_data = 12'b001000000000;
		14'b01100011100000: color_data = 12'b001000000000;
		14'b01100011100001: color_data = 12'b010000000000;
		14'b01100011100010: color_data = 12'b010000000000;
		14'b01100011100011: color_data = 12'b010000000000;
		14'b01100011100100: color_data = 12'b010000000000;
		14'b01100011100101: color_data = 12'b001000000000;
		14'b01100011100110: color_data = 12'b010000000000;
		14'b01100011100111: color_data = 12'b010000000000;
		14'b01100011101000: color_data = 12'b010000000000;
		14'b01100011101001: color_data = 12'b010000000000;
		14'b01100011101010: color_data = 12'b010000000000;
		14'b01100011101011: color_data = 12'b001000000000;
		14'b01100100010000: color_data = 12'b001000000000;
		14'b01100100010001: color_data = 12'b001000000000;
		14'b01100100010010: color_data = 12'b010000000000;
		14'b01100100010011: color_data = 12'b010000000000;
		14'b01100100010100: color_data = 12'b010000000000;
		14'b01100100010101: color_data = 12'b010000000000;
		14'b01100100011011: color_data = 12'b001000000000;
		14'b01100100011100: color_data = 12'b010000000000;
		14'b01100100011101: color_data = 12'b010000000000;
		14'b01100100011110: color_data = 12'b010000000000;
		14'b01100100011111: color_data = 12'b010000000000;
		14'b01100100100000: color_data = 12'b010000000000;
		14'b01100100100001: color_data = 12'b010000000000;
		14'b01100100100011: color_data = 12'b001000000000;
		14'b01100100100111: color_data = 12'b001000000000;
		14'b01100100101000: color_data = 12'b001000000000;
		14'b01100100101001: color_data = 12'b010000000000;
		14'b01100100101010: color_data = 12'b010000000000;
		14'b01100100101011: color_data = 12'b010000000000;
		14'b01100100101100: color_data = 12'b010000000000;
		14'b01100100101101: color_data = 12'b010000000000;
		14'b01100100101110: color_data = 12'b010000000000;
		14'b01100100101111: color_data = 12'b010000000000;
		14'b01100100110000: color_data = 12'b010000000000;
		14'b01100100110001: color_data = 12'b001000000000;
		14'b01100100110010: color_data = 12'b001000000000;
		14'b01100100110011: color_data = 12'b001000000000;
		14'b01100100110100: color_data = 12'b001000000000;
		14'b01100100110101: color_data = 12'b001000000000;
		14'b01100100110110: color_data = 12'b010000000000;
		14'b01100100110111: color_data = 12'b010000000000;
		14'b01100100111000: color_data = 12'b010000000000;
		14'b01100100111001: color_data = 12'b010000000000;
		14'b01100100111010: color_data = 12'b010000000000;
		14'b01100100111011: color_data = 12'b010000000000;
		14'b01100100111100: color_data = 12'b010000000000;
		14'b01100100111101: color_data = 12'b010000000000;
		14'b01100100111110: color_data = 12'b010000000000;
		14'b01100100111111: color_data = 12'b010000000000;
		14'b01100101000000: color_data = 12'b010000000000;
		14'b01100101000001: color_data = 12'b001000000000;
		14'b01100101000010: color_data = 12'b001000000000;
		14'b01100101000011: color_data = 12'b001000000000;
		14'b01100101000100: color_data = 12'b001000000000;
		14'b01100101000101: color_data = 12'b001000000000;
		14'b01100101000110: color_data = 12'b001000000000;
		14'b01100101011111: color_data = 12'b001000000000;
		14'b01100101100000: color_data = 12'b001000000000;
		14'b01100101100001: color_data = 12'b001000000000;
		14'b01100101100010: color_data = 12'b001000000000;
		14'b01100101100011: color_data = 12'b010000000000;
		14'b01100101100100: color_data = 12'b010000000000;
		14'b01100101100101: color_data = 12'b001000000000;
		14'b01100101100110: color_data = 12'b001000000000;
		14'b01100101100111: color_data = 12'b010000000000;
		14'b01100101101000: color_data = 12'b010000000000;
		14'b01100101101001: color_data = 12'b010000000000;
		14'b01100101101010: color_data = 12'b010000000000;
		14'b01100101101011: color_data = 12'b010000000000;
		14'b01100101101100: color_data = 12'b001000000000;
		14'b01100110010011: color_data = 12'b001000000000;
		14'b01100110010100: color_data = 12'b010000000000;
		14'b01100110010101: color_data = 12'b010000000000;
		14'b01100110010110: color_data = 12'b010000000000;
		14'b01100110011110: color_data = 12'b001000000000;
		14'b01100110011111: color_data = 12'b010000000000;
		14'b01100110100000: color_data = 12'b010000000000;
		14'b01100110100001: color_data = 12'b010000000000;
		14'b01100110100010: color_data = 12'b010000000000;
		14'b01100110100011: color_data = 12'b010000000000;
		14'b01100110101010: color_data = 12'b010000000000;
		14'b01100110101011: color_data = 12'b010000000000;
		14'b01100110101100: color_data = 12'b010000000000;
		14'b01100110101101: color_data = 12'b010000000000;
		14'b01100110101110: color_data = 12'b010000000000;
		14'b01100110101111: color_data = 12'b010000000000;
		14'b01100110110000: color_data = 12'b010000000000;
		14'b01100110110001: color_data = 12'b010000000000;
		14'b01100110110010: color_data = 12'b010000000000;
		14'b01100110110011: color_data = 12'b001000000000;
		14'b01100110110100: color_data = 12'b001000000000;
		14'b01100110110101: color_data = 12'b001000000000;
		14'b01100110110110: color_data = 12'b010000000000;
		14'b01100110110111: color_data = 12'b010000000000;
		14'b01100110111000: color_data = 12'b010000000000;
		14'b01100110111001: color_data = 12'b010000000000;
		14'b01100110111010: color_data = 12'b010000000000;
		14'b01100110111011: color_data = 12'b010000000000;
		14'b01100110111100: color_data = 12'b010000000000;
		14'b01100110111101: color_data = 12'b010000000000;
		14'b01100110111110: color_data = 12'b010000000000;
		14'b01100110111111: color_data = 12'b001000000000;
		14'b01100111000000: color_data = 12'b001000000000;
		14'b01100111000001: color_data = 12'b001000000000;
		14'b01100111000010: color_data = 12'b001000000000;
		14'b01100111000011: color_data = 12'b001000000000;
		14'b01100111000100: color_data = 12'b001000000000;
		14'b01100111100011: color_data = 12'b001000000000;
		14'b01100111100100: color_data = 12'b001000000000;
		14'b01100111100101: color_data = 12'b001000000000;
		14'b01100111100110: color_data = 12'b001000000000;
		14'b01100111100111: color_data = 12'b010000000000;
		14'b01100111101000: color_data = 12'b010000000000;
		14'b01100111101001: color_data = 12'b010000000000;
		14'b01100111101010: color_data = 12'b010000000000;
		14'b01100111101011: color_data = 12'b010000000000;
		14'b01100111101100: color_data = 12'b010000000000;
		14'b01100111101101: color_data = 12'b010000000000;
		14'b01101000010101: color_data = 12'b001000000000;
		14'b01101000010110: color_data = 12'b010000000000;
		14'b01101000010111: color_data = 12'b010000000000;
		14'b01101000011000: color_data = 12'b001000000000;
		14'b01101000011111: color_data = 12'b001000000000;
		14'b01101000100000: color_data = 12'b010000000000;
		14'b01101000100001: color_data = 12'b010000000000;
		14'b01101000100010: color_data = 12'b010000000000;
		14'b01101000100011: color_data = 12'b010000000000;
		14'b01101000100100: color_data = 12'b010000000000;
		14'b01101000100101: color_data = 12'b001000000000;
		14'b01101000101011: color_data = 12'b001000000000;
		14'b01101000101100: color_data = 12'b010000000000;
		14'b01101000101101: color_data = 12'b010000000000;
		14'b01101000101110: color_data = 12'b010000000000;
		14'b01101000101111: color_data = 12'b010000000000;
		14'b01101000110000: color_data = 12'b010000000000;
		14'b01101000110001: color_data = 12'b010000000000;
		14'b01101000110010: color_data = 12'b010000000000;
		14'b01101000110011: color_data = 12'b010000000000;
		14'b01101000110100: color_data = 12'b010000000000;
		14'b01101000110101: color_data = 12'b010000000000;
		14'b01101000110110: color_data = 12'b010000000000;
		14'b01101000110111: color_data = 12'b010000000000;
		14'b01101000111000: color_data = 12'b010000000000;
		14'b01101000111001: color_data = 12'b010000000000;
		14'b01101000111010: color_data = 12'b010000000000;
		14'b01101000111011: color_data = 12'b010000000000;
		14'b01101000111100: color_data = 12'b010000000000;
		14'b01101000111101: color_data = 12'b001000000000;
		14'b01101000111110: color_data = 12'b001000000000;
		14'b01101000111111: color_data = 12'b001000000000;
		14'b01101001000000: color_data = 12'b001000000000;
		14'b01101001000001: color_data = 12'b001000000000;
		14'b01101001000010: color_data = 12'b001000000000;
		14'b01101001000011: color_data = 12'b001000000000;
		14'b01101001100101: color_data = 12'b001000000000;
		14'b01101001100110: color_data = 12'b001000000000;
		14'b01101001100111: color_data = 12'b010000000000;
		14'b01101001101000: color_data = 12'b010000000000;
		14'b01101001101001: color_data = 12'b010000000000;
		14'b01101001101010: color_data = 12'b010000000000;
		14'b01101001101011: color_data = 12'b010000000000;
		14'b01101001101100: color_data = 12'b010000000000;
		14'b01101001101101: color_data = 12'b010000000000;
		14'b01101001101110: color_data = 12'b001000000000;
		14'b01101010010110: color_data = 12'b001000000000;
		14'b01101010010111: color_data = 12'b010000000000;
		14'b01101010011000: color_data = 12'b010000000000;
		14'b01101010011001: color_data = 12'b010000000000;
		14'b01101010100000: color_data = 12'b001000000000;
		14'b01101010100001: color_data = 12'b010000000000;
		14'b01101010100010: color_data = 12'b010000000000;
		14'b01101010100011: color_data = 12'b010000000000;
		14'b01101010100100: color_data = 12'b010000000000;
		14'b01101010100101: color_data = 12'b010000000000;
		14'b01101010100110: color_data = 12'b010000000000;
		14'b01101010101101: color_data = 12'b001000000000;
		14'b01101010101110: color_data = 12'b010000000000;
		14'b01101010101111: color_data = 12'b010000000000;
		14'b01101010110000: color_data = 12'b010000000000;
		14'b01101010110001: color_data = 12'b010000000000;
		14'b01101010110010: color_data = 12'b010000000000;
		14'b01101010110011: color_data = 12'b010000000000;
		14'b01101010110100: color_data = 12'b010000000000;
		14'b01101010110101: color_data = 12'b010000000000;
		14'b01101010110110: color_data = 12'b010000000000;
		14'b01101010110111: color_data = 12'b010000000000;
		14'b01101010111000: color_data = 12'b010000000000;
		14'b01101010111001: color_data = 12'b010000000000;
		14'b01101010111010: color_data = 12'b010000000000;
		14'b01101010111011: color_data = 12'b001000000000;
		14'b01101010111101: color_data = 12'b001000000000;
		14'b01101010111110: color_data = 12'b001000000000;
		14'b01101010111111: color_data = 12'b010000000000;
		14'b01101011000000: color_data = 12'b001000000000;
		14'b01101011000001: color_data = 12'b001000000000;
		14'b01101011000010: color_data = 12'b001000000000;
		14'b01101011100111: color_data = 12'b001000000000;
		14'b01101011101000: color_data = 12'b001000000000;
		14'b01101011101001: color_data = 12'b001000000000;
		14'b01101011101010: color_data = 12'b010000000000;
		14'b01101011101011: color_data = 12'b010000000000;
		14'b01101011101100: color_data = 12'b010000000000;
		14'b01101011101101: color_data = 12'b010000000000;
		14'b01101011101110: color_data = 12'b010000000000;
		14'b01101100010111: color_data = 12'b001000000000;
		14'b01101100011000: color_data = 12'b010000000000;
		14'b01101100011001: color_data = 12'b010000000000;
		14'b01101100011010: color_data = 12'b010000000000;
		14'b01101100100001: color_data = 12'b001000000000;
		14'b01101100100010: color_data = 12'b010000000000;
		14'b01101100100011: color_data = 12'b010000000000;
		14'b01101100100100: color_data = 12'b010000000000;
		14'b01101100100101: color_data = 12'b010000000000;
		14'b01101100100110: color_data = 12'b010000000000;
		14'b01101100100111: color_data = 12'b010000000000;
		14'b01101100101000: color_data = 12'b001000000000;
		14'b01101100101110: color_data = 12'b001000000000;
		14'b01101100101111: color_data = 12'b010000000000;
		14'b01101100110000: color_data = 12'b010000000000;
		14'b01101100110001: color_data = 12'b010000000000;
		14'b01101100110010: color_data = 12'b010000000000;
		14'b01101100110011: color_data = 12'b010000000000;
		14'b01101100110100: color_data = 12'b010000000000;
		14'b01101100110101: color_data = 12'b010000000000;
		14'b01101100110110: color_data = 12'b010000000000;
		14'b01101100110111: color_data = 12'b010000000000;
		14'b01101100111000: color_data = 12'b010000000000;
		14'b01101100111001: color_data = 12'b001000000000;
		14'b01101100111010: color_data = 12'b001000000000;
		14'b01101100111101: color_data = 12'b010000000000;
		14'b01101100111110: color_data = 12'b001000000000;
		14'b01101100111111: color_data = 12'b001000000000;
		14'b01101101000000: color_data = 12'b001000000000;
		14'b01101101000001: color_data = 12'b001000000000;
		14'b01101101000010: color_data = 12'b001000000000;
		14'b01101101101001: color_data = 12'b001000000000;
		14'b01101101101010: color_data = 12'b001000000000;
		14'b01101101101011: color_data = 12'b010000000000;
		14'b01101101101100: color_data = 12'b010000000000;
		14'b01101101101101: color_data = 12'b010000000000;
		14'b01101101101110: color_data = 12'b010000000000;
		14'b01101101101111: color_data = 12'b010000000000;
		14'b01101101110110: color_data = 12'b001000000000;
		14'b01101110011000: color_data = 12'b010000000000;
		14'b01101110011001: color_data = 12'b010000000000;
		14'b01101110011010: color_data = 12'b010000000000;
		14'b01101110011011: color_data = 12'b010000000000;
		14'b01101110011100: color_data = 12'b001000000000;
		14'b01101110100010: color_data = 12'b010000000000;
		14'b01101110100011: color_data = 12'b010000000000;
		14'b01101110100100: color_data = 12'b010000000000;
		14'b01101110100101: color_data = 12'b010000000000;
		14'b01101110100110: color_data = 12'b010000000000;
		14'b01101110100111: color_data = 12'b010000000000;
		14'b01101110101000: color_data = 12'b010000000000;
		14'b01101110101111: color_data = 12'b001000000000;
		14'b01101110110000: color_data = 12'b010000000000;
		14'b01101110110001: color_data = 12'b010000000000;
		14'b01101110110010: color_data = 12'b010000000000;
		14'b01101110110011: color_data = 12'b010000000000;
		14'b01101110110100: color_data = 12'b010000000000;
		14'b01101110110101: color_data = 12'b010000000000;
		14'b01101110110110: color_data = 12'b001000000000;
		14'b01101110110111: color_data = 12'b001000000000;
		14'b01101110111000: color_data = 12'b001000000000;
		14'b01101110111100: color_data = 12'b010000000000;
		14'b01101110111101: color_data = 12'b010000000000;
		14'b01101110111110: color_data = 12'b001000000000;
		14'b01101110111111: color_data = 12'b001000000000;
		14'b01101111000000: color_data = 12'b001000000000;
		14'b01101111101010: color_data = 12'b001000000000;
		14'b01101111101011: color_data = 12'b001000000000;
		14'b01101111101100: color_data = 12'b010000000000;
		14'b01101111101101: color_data = 12'b010000000000;
		14'b01101111101110: color_data = 12'b010000000000;
		14'b01101111101111: color_data = 12'b010000000000;
		14'b01101111110000: color_data = 12'b010000000000;
		14'b01101111110111: color_data = 12'b001000000000;
		14'b01110000011001: color_data = 12'b010000000000;
		14'b01110000011010: color_data = 12'b010000000000;
		14'b01110000011011: color_data = 12'b010000000000;
		14'b01110000011100: color_data = 12'b010000000000;
		14'b01110000011101: color_data = 12'b010000000000;
		14'b01110000100011: color_data = 12'b010000000000;
		14'b01110000100100: color_data = 12'b010000000000;
		14'b01110000100101: color_data = 12'b010000000000;
		14'b01110000100110: color_data = 12'b010000000000;
		14'b01110000100111: color_data = 12'b010000000000;
		14'b01110000101000: color_data = 12'b010000000000;
		14'b01110000101001: color_data = 12'b010000000000;
		14'b01110000101010: color_data = 12'b001000000000;
		14'b01110000101011: color_data = 12'b001000000000;
		14'b01110000101100: color_data = 12'b001000000000;
		14'b01110000110001: color_data = 12'b010000000000;
		14'b01110000110010: color_data = 12'b010000000000;
		14'b01110000110011: color_data = 12'b010000000000;
		14'b01110000110100: color_data = 12'b010000000000;
		14'b01110000111010: color_data = 12'b001000000000;
		14'b01110000111011: color_data = 12'b010000000000;
		14'b01110000111100: color_data = 12'b010000000000;
		14'b01110000111101: color_data = 12'b001000000000;
		14'b01110000111110: color_data = 12'b001000000000;
		14'b01110001101011: color_data = 12'b001000000000;
		14'b01110001101100: color_data = 12'b010000000000;
		14'b01110001101101: color_data = 12'b010000000000;
		14'b01110001101110: color_data = 12'b010000000000;
		14'b01110001101111: color_data = 12'b010000000000;
		14'b01110001110000: color_data = 12'b010000000000;
		14'b01110001110001: color_data = 12'b010000000000;
		14'b01110001111000: color_data = 12'b001000000000;
		14'b01110010011010: color_data = 12'b001000000000;
		14'b01110010011011: color_data = 12'b010000000000;
		14'b01110010011100: color_data = 12'b010000000000;
		14'b01110010011101: color_data = 12'b010000000000;
		14'b01110010011110: color_data = 12'b001000000000;
		14'b01110010100100: color_data = 12'b010000000000;
		14'b01110010100101: color_data = 12'b010000000000;
		14'b01110010100110: color_data = 12'b010000000000;
		14'b01110010100111: color_data = 12'b010000000000;
		14'b01110010101000: color_data = 12'b010000000000;
		14'b01110010101001: color_data = 12'b010000000000;
		14'b01110010101010: color_data = 12'b010000000000;
		14'b01110010101011: color_data = 12'b001000000000;
		14'b01110010101100: color_data = 12'b001000000000;
		14'b01110010101101: color_data = 12'b001000000000;
		14'b01110010110010: color_data = 12'b001000000000;
		14'b01110010111001: color_data = 12'b001000000000;
		14'b01110010111010: color_data = 12'b001000000000;
		14'b01110010111011: color_data = 12'b010000000000;
		14'b01110010111100: color_data = 12'b001000000000;
		14'b01110011010011: color_data = 12'b001000000000;
		14'b01110011101100: color_data = 12'b010000000000;
		14'b01110011101101: color_data = 12'b010000000000;
		14'b01110011101110: color_data = 12'b010000000000;
		14'b01110011101111: color_data = 12'b010000000000;
		14'b01110011110000: color_data = 12'b010000000000;
		14'b01110011110001: color_data = 12'b010000000000;
		14'b01110011110010: color_data = 12'b001000000000;
		14'b01110011111001: color_data = 12'b001000000000;
		14'b01110100011100: color_data = 12'b010000000000;
		14'b01110100011101: color_data = 12'b010000000000;
		14'b01110100011110: color_data = 12'b010000000000;
		14'b01110100011111: color_data = 12'b001000000000;
		14'b01110100100101: color_data = 12'b010000000000;
		14'b01110100100110: color_data = 12'b010000000000;
		14'b01110100100111: color_data = 12'b010000000000;
		14'b01110100101000: color_data = 12'b010000000000;
		14'b01110100101001: color_data = 12'b010000000000;
		14'b01110100101010: color_data = 12'b010000000000;
		14'b01110100101011: color_data = 12'b010000000000;
		14'b01110100101100: color_data = 12'b010000000000;
		14'b01110100101101: color_data = 12'b001000000000;
		14'b01110100101110: color_data = 12'b001000000000;
		14'b01110100110111: color_data = 12'b001000000000;
		14'b01110100111000: color_data = 12'b001000000000;
		14'b01110100111001: color_data = 12'b010000000000;
		14'b01110100111010: color_data = 12'b010000000000;
		14'b01110101010100: color_data = 12'b001000000000;
		14'b01110101010101: color_data = 12'b001000000000;
		14'b01110101010110: color_data = 12'b001000000000;
		14'b01110101101101: color_data = 12'b010000000000;
		14'b01110101101110: color_data = 12'b010000000000;
		14'b01110101101111: color_data = 12'b010000000000;
		14'b01110101110000: color_data = 12'b010000000000;
		14'b01110101110001: color_data = 12'b010000000000;
		14'b01110101110010: color_data = 12'b010000000000;
		14'b01110101110011: color_data = 12'b001000000000;
		14'b01110101111010: color_data = 12'b001000000000;
		14'b01110110011110: color_data = 12'b010000000000;
		14'b01110110011111: color_data = 12'b010000000000;
		14'b01110110100000: color_data = 12'b001000000000;
		14'b01110110100110: color_data = 12'b010000000000;
		14'b01110110100111: color_data = 12'b010000000000;
		14'b01110110101000: color_data = 12'b010000000000;
		14'b01110110101001: color_data = 12'b010000000000;
		14'b01110110101010: color_data = 12'b010000000000;
		14'b01110110101011: color_data = 12'b010000000000;
		14'b01110110101100: color_data = 12'b010000000000;
		14'b01110110101101: color_data = 12'b001000000000;
		14'b01110110101110: color_data = 12'b001000000000;
		14'b01110110101111: color_data = 12'b001000000000;
		14'b01110110110000: color_data = 12'b001000000000;
		14'b01110110110110: color_data = 12'b001000000000;
		14'b01110110110111: color_data = 12'b001000000000;
		14'b01110110111000: color_data = 12'b010000000000;
		14'b01110110111001: color_data = 12'b010000000000;
		14'b01110111010100: color_data = 12'b001000000000;
		14'b01110111010101: color_data = 12'b001000000000;
		14'b01110111010110: color_data = 12'b001000000000;
		14'b01110111010111: color_data = 12'b001000000000;
		14'b01110111101110: color_data = 12'b001000000000;
		14'b01110111101111: color_data = 12'b010000000000;
		14'b01110111110000: color_data = 12'b010000000000;
		14'b01110111110001: color_data = 12'b010000000000;
		14'b01110111110010: color_data = 12'b010000000000;
		14'b01110111110011: color_data = 12'b010000000000;
		14'b01110111110100: color_data = 12'b001000000000;
		14'b01110111111011: color_data = 12'b001000000000;
		14'b01111000011111: color_data = 12'b010000000000;
		14'b01111000100000: color_data = 12'b010000000000;
		14'b01111000100001: color_data = 12'b001000000000;
		14'b01111000100111: color_data = 12'b010000000000;
		14'b01111000101000: color_data = 12'b010000000000;
		14'b01111000101001: color_data = 12'b010000000000;
		14'b01111000101010: color_data = 12'b010000000000;
		14'b01111000101011: color_data = 12'b010000000000;
		14'b01111000101100: color_data = 12'b010000000000;
		14'b01111000101101: color_data = 12'b010000000000;
		14'b01111000101110: color_data = 12'b001000000000;
		14'b01111000101111: color_data = 12'b001000000000;
		14'b01111000110000: color_data = 12'b001000000000;
		14'b01111000110001: color_data = 12'b001000000000;
		14'b01111000110010: color_data = 12'b001000000000;
		14'b01111000110011: color_data = 12'b001000000000;
		14'b01111000110100: color_data = 12'b001000000000;
		14'b01111000110101: color_data = 12'b001000000000;
		14'b01111000110110: color_data = 12'b001000000000;
		14'b01111000110111: color_data = 12'b010000000000;
		14'b01111000111000: color_data = 12'b010000000000;
		14'b01111001010100: color_data = 12'b001000000000;
		14'b01111001010101: color_data = 12'b001000000000;
		14'b01111001010110: color_data = 12'b001000000000;
		14'b01111001010111: color_data = 12'b001000000000;
		14'b01111001101110: color_data = 12'b001000000000;
		14'b01111001110000: color_data = 12'b010000000000;
		14'b01111001110001: color_data = 12'b010000000000;
		14'b01111001110010: color_data = 12'b010000000000;
		14'b01111001110011: color_data = 12'b010000000000;
		14'b01111001110100: color_data = 12'b010000000000;
		14'b01111001110101: color_data = 12'b010000000000;
		14'b01111001111011: color_data = 12'b001000000000;
		14'b01111010011111: color_data = 12'b001000000000;
		14'b01111010100000: color_data = 12'b010000000000;
		14'b01111010100001: color_data = 12'b010000000000;
		14'b01111010100111: color_data = 12'b010000000000;
		14'b01111010101000: color_data = 12'b010000000000;
		14'b01111010101001: color_data = 12'b010000000000;
		14'b01111010101010: color_data = 12'b010000000000;
		14'b01111010101011: color_data = 12'b010000000000;
		14'b01111010101100: color_data = 12'b010000000000;
		14'b01111010101101: color_data = 12'b010000000000;
		14'b01111010101110: color_data = 12'b001000000000;
		14'b01111010101111: color_data = 12'b001000000000;
		14'b01111010110000: color_data = 12'b001000000000;
		14'b01111010110001: color_data = 12'b001000000000;
		14'b01111010110010: color_data = 12'b001000000000;
		14'b01111010110011: color_data = 12'b001000000000;
		14'b01111010110100: color_data = 12'b001000000000;
		14'b01111010110101: color_data = 12'b001000000000;
		14'b01111010110110: color_data = 12'b010000000000;
		14'b01111010110111: color_data = 12'b010000000000;
		14'b01111010111000: color_data = 12'b001000000000;
		14'b01111011000011: color_data = 12'b001000000000;
		14'b01111011000100: color_data = 12'b001000000000;
		14'b01111011000101: color_data = 12'b001000000000;
		14'b01111011001110: color_data = 12'b001000000000;
		14'b01111011001111: color_data = 12'b001000000000;
		14'b01111011010000: color_data = 12'b001000000000;
		14'b01111011010100: color_data = 12'b001000000000;
		14'b01111011010101: color_data = 12'b001000000000;
		14'b01111011010110: color_data = 12'b001000000000;
		14'b01111011010111: color_data = 12'b001000000000;
		14'b01111011011000: color_data = 12'b001000000000;
		14'b01111011110000: color_data = 12'b001000000000;
		14'b01111011110001: color_data = 12'b010000000000;
		14'b01111011110010: color_data = 12'b010000000000;
		14'b01111011110011: color_data = 12'b010000000000;
		14'b01111011110100: color_data = 12'b010000000000;
		14'b01111011110101: color_data = 12'b010000000000;
		14'b01111011110110: color_data = 12'b010000000000;
		14'b01111011110111: color_data = 12'b001000000000;
		14'b01111011111100: color_data = 12'b001000000000;
		14'b01111100100000: color_data = 12'b001000000000;
		14'b01111100100001: color_data = 12'b010000000000;
		14'b01111100100010: color_data = 12'b001000000000;
		14'b01111100100111: color_data = 12'b001000000000;
		14'b01111100101000: color_data = 12'b010000000000;
		14'b01111100101001: color_data = 12'b010000000000;
		14'b01111100101010: color_data = 12'b010000000000;
		14'b01111100101011: color_data = 12'b010000000000;
		14'b01111100101100: color_data = 12'b010000000000;
		14'b01111100101101: color_data = 12'b010000000000;
		14'b01111100101110: color_data = 12'b001000000000;
		14'b01111100101111: color_data = 12'b001000000000;
		14'b01111100110000: color_data = 12'b001000000000;
		14'b01111100110001: color_data = 12'b001000000000;
		14'b01111100110010: color_data = 12'b001000000000;
		14'b01111100110011: color_data = 12'b001000000000;
		14'b01111100110100: color_data = 12'b001000000000;
		14'b01111100110101: color_data = 12'b010000000000;
		14'b01111100110110: color_data = 12'b010000000000;
		14'b01111100110111: color_data = 12'b010000000000;
		14'b01111100111000: color_data = 12'b001000000000;
		14'b01111101000000: color_data = 12'b001000000000;
		14'b01111101000001: color_data = 12'b001000000000;
		14'b01111101000010: color_data = 12'b001000000000;
		14'b01111101000011: color_data = 12'b001000000000;
		14'b01111101000100: color_data = 12'b001000000000;
		14'b01111101000101: color_data = 12'b001000000000;
		14'b01111101000110: color_data = 12'b001000000000;
		14'b01111101000111: color_data = 12'b001000000000;
		14'b01111101001000: color_data = 12'b001000000000;
		14'b01111101001001: color_data = 12'b001000000000;
		14'b01111101001010: color_data = 12'b001000000000;
		14'b01111101001011: color_data = 12'b001000000000;
		14'b01111101001100: color_data = 12'b001000000000;
		14'b01111101001101: color_data = 12'b001000000000;
		14'b01111101001110: color_data = 12'b010000000000;
		14'b01111101001111: color_data = 12'b001000000000;
		14'b01111101010000: color_data = 12'b001000000000;
		14'b01111101010001: color_data = 12'b010000000000;
		14'b01111101010010: color_data = 12'b001000000000;
		14'b01111101010011: color_data = 12'b001000000000;
		14'b01111101010100: color_data = 12'b001000000000;
		14'b01111101010101: color_data = 12'b001000000000;
		14'b01111101010110: color_data = 12'b001000000000;
		14'b01111101010111: color_data = 12'b001000000000;
		14'b01111101011000: color_data = 12'b001000000000;
		14'b01111101110001: color_data = 12'b001000000000;
		14'b01111101110010: color_data = 12'b010000000000;
		14'b01111101110011: color_data = 12'b010000000000;
		14'b01111101110100: color_data = 12'b010000000000;
		14'b01111101110101: color_data = 12'b010000000000;
		14'b01111101110110: color_data = 12'b010000000000;
		14'b01111101110111: color_data = 12'b010000000000;
		14'b01111101111000: color_data = 12'b001000000000;
		14'b01111110100001: color_data = 12'b010000000000;
		14'b01111110100010: color_data = 12'b001000000000;
		14'b01111110101000: color_data = 12'b010000000000;
		14'b01111110101001: color_data = 12'b010000000000;
		14'b01111110101010: color_data = 12'b010000000000;
		14'b01111110101011: color_data = 12'b010000000000;
		14'b01111110101100: color_data = 12'b010000000000;
		14'b01111110101101: color_data = 12'b010000000000;
		14'b01111110101110: color_data = 12'b010000000000;
		14'b01111110101111: color_data = 12'b001000000000;
		14'b01111110110000: color_data = 12'b001000000000;
		14'b01111110110001: color_data = 12'b001000000000;
		14'b01111110110010: color_data = 12'b001000000000;
		14'b01111110110011: color_data = 12'b001000000000;
		14'b01111110110100: color_data = 12'b010000000000;
		14'b01111110110101: color_data = 12'b010000000000;
		14'b01111110110110: color_data = 12'b010000000000;
		14'b01111110110111: color_data = 12'b001000000000;
		14'b01111111000000: color_data = 12'b001000000000;
		14'b01111111000101: color_data = 12'b001000000000;
		14'b01111111000110: color_data = 12'b001000000000;
		14'b01111111000111: color_data = 12'b001000000000;
		14'b01111111001000: color_data = 12'b001000000000;
		14'b01111111001001: color_data = 12'b001000000000;
		14'b01111111001010: color_data = 12'b010000000000;
		14'b01111111001011: color_data = 12'b001000000000;
		14'b01111111001100: color_data = 12'b001000000000;
		14'b01111111001101: color_data = 12'b010000000000;
		14'b01111111001110: color_data = 12'b010000000000;
		14'b01111111001111: color_data = 12'b010000000000;
		14'b01111111010000: color_data = 12'b001000000000;
		14'b01111111010001: color_data = 12'b010000000000;
		14'b01111111010010: color_data = 12'b010000000000;
		14'b01111111010011: color_data = 12'b010000000000;
		14'b01111111010100: color_data = 12'b001000000000;
		14'b01111111010101: color_data = 12'b001000000000;
		14'b01111111010110: color_data = 12'b001000000000;
		14'b01111111010111: color_data = 12'b001000000000;
		14'b01111111011000: color_data = 12'b001000000000;
		14'b01111111011001: color_data = 12'b001000000000;
		14'b01111111110001: color_data = 12'b001000000000;
		14'b01111111110010: color_data = 12'b001000000000;
		14'b01111111110011: color_data = 12'b010000000000;
		14'b01111111110100: color_data = 12'b010000000000;
		14'b01111111110101: color_data = 12'b010000000000;
		14'b01111111110110: color_data = 12'b010000000000;
		14'b01111111110111: color_data = 12'b010000000000;
		14'b01111111111000: color_data = 12'b010000000000;
		14'b01111111111001: color_data = 12'b001000000000;
		14'b01111111111101: color_data = 12'b001000000000;
		14'b10000000100001: color_data = 12'b001000000000;
		14'b10000000100010: color_data = 12'b010000000000;
		14'b10000000101000: color_data = 12'b010000000000;
		14'b10000000101001: color_data = 12'b010000000000;
		14'b10000000101010: color_data = 12'b010000000000;
		14'b10000000101011: color_data = 12'b010000000000;
		14'b10000000101100: color_data = 12'b010000000000;
		14'b10000000101101: color_data = 12'b010000000000;
		14'b10000000101110: color_data = 12'b010000000000;
		14'b10000000101111: color_data = 12'b001000000000;
		14'b10000000110000: color_data = 12'b001000000000;
		14'b10000000110001: color_data = 12'b001000000000;
		14'b10000000110010: color_data = 12'b001000000000;
		14'b10000000110011: color_data = 12'b010000000000;
		14'b10000000110100: color_data = 12'b010000000000;
		14'b10000000110101: color_data = 12'b010000000000;
		14'b10000000110110: color_data = 12'b001000000000;
		14'b10000001000101: color_data = 12'b001000000000;
		14'b10000001000110: color_data = 12'b001000000000;
		14'b10000001000111: color_data = 12'b001000000000;
		14'b10000001001000: color_data = 12'b010000000000;
		14'b10000001001001: color_data = 12'b001000000000;
		14'b10000001001010: color_data = 12'b001000000000;
		14'b10000001001011: color_data = 12'b001000000000;
		14'b10000001001100: color_data = 12'b001000000000;
		14'b10000001001101: color_data = 12'b010000000000;
		14'b10000001001110: color_data = 12'b010000000000;
		14'b10000001001111: color_data = 12'b010000000000;
		14'b10000001010000: color_data = 12'b001000000000;
		14'b10000001010001: color_data = 12'b010000000000;
		14'b10000001010010: color_data = 12'b010000000000;
		14'b10000001010011: color_data = 12'b010000000000;
		14'b10000001010100: color_data = 12'b010000000000;
		14'b10000001010101: color_data = 12'b010000000000;
		14'b10000001010110: color_data = 12'b001000000000;
		14'b10000001010111: color_data = 12'b001000000000;
		14'b10000001011000: color_data = 12'b001000000000;
		14'b10000001011001: color_data = 12'b001000000000;
		14'b10000001110010: color_data = 12'b001000000000;
		14'b10000001110011: color_data = 12'b001000000000;
		14'b10000001110100: color_data = 12'b010000000000;
		14'b10000001110101: color_data = 12'b010000000000;
		14'b10000001110110: color_data = 12'b010000000000;
		14'b10000001110111: color_data = 12'b010000000000;
		14'b10000001111000: color_data = 12'b010000000000;
		14'b10000001111001: color_data = 12'b010000000000;
		14'b10000001111010: color_data = 12'b001000000000;
		14'b10000001111101: color_data = 12'b001000000000;
		14'b10000010100001: color_data = 12'b001000000000;
		14'b10000010100010: color_data = 12'b010000000000;
		14'b10000010101000: color_data = 12'b010000000000;
		14'b10000010101001: color_data = 12'b010000000000;
		14'b10000010101010: color_data = 12'b010000000000;
		14'b10000010101011: color_data = 12'b010000000000;
		14'b10000010101100: color_data = 12'b010000000000;
		14'b10000010101101: color_data = 12'b010000000000;
		14'b10000010101110: color_data = 12'b010000000000;
		14'b10000010101111: color_data = 12'b001000000000;
		14'b10000010110000: color_data = 12'b001000000000;
		14'b10000010110001: color_data = 12'b001000000000;
		14'b10000010110010: color_data = 12'b010000000000;
		14'b10000010110011: color_data = 12'b010000000000;
		14'b10000010110100: color_data = 12'b010000000000;
		14'b10000010110101: color_data = 12'b010000000000;
		14'b10000010110110: color_data = 12'b001000000000;
		14'b10000011000101: color_data = 12'b001000000000;
		14'b10000011000110: color_data = 12'b001000000000;
		14'b10000011000111: color_data = 12'b010000000000;
		14'b10000011001000: color_data = 12'b010000000000;
		14'b10000011001001: color_data = 12'b010000000000;
		14'b10000011001010: color_data = 12'b010000000000;
		14'b10000011001011: color_data = 12'b001000000000;
		14'b10000011001100: color_data = 12'b010000000000;
		14'b10000011001101: color_data = 12'b010000000000;
		14'b10000011001110: color_data = 12'b010000000000;
		14'b10000011001111: color_data = 12'b010000000000;
		14'b10000011010000: color_data = 12'b010000000000;
		14'b10000011010001: color_data = 12'b010000000000;
		14'b10000011010010: color_data = 12'b010000000000;
		14'b10000011010011: color_data = 12'b010000000000;
		14'b10000011010100: color_data = 12'b010000000000;
		14'b10000011010101: color_data = 12'b010000000000;
		14'b10000011010110: color_data = 12'b010000000000;
		14'b10000011010111: color_data = 12'b010000000000;
		14'b10000011011000: color_data = 12'b010000000000;
		14'b10000011011001: color_data = 12'b001000000000;
		14'b10000011011010: color_data = 12'b001000000000;
		14'b10000011110011: color_data = 12'b001000000000;
		14'b10000011110100: color_data = 12'b001000000000;
		14'b10000011110101: color_data = 12'b010000000000;
		14'b10000011110110: color_data = 12'b010000000000;
		14'b10000011110111: color_data = 12'b010000000000;
		14'b10000011111000: color_data = 12'b010000000000;
		14'b10000011111001: color_data = 12'b010000000000;
		14'b10000011111010: color_data = 12'b010000000000;
		14'b10000011111011: color_data = 12'b001000000000;
		14'b10000100100001: color_data = 12'b001000000000;
		14'b10000100100010: color_data = 12'b001000000000;
		14'b10000100101000: color_data = 12'b010000000000;
		14'b10000100101001: color_data = 12'b010000000000;
		14'b10000100101010: color_data = 12'b010000000000;
		14'b10000100101011: color_data = 12'b010000000000;
		14'b10000100101100: color_data = 12'b010000000000;
		14'b10000100101101: color_data = 12'b010000000000;
		14'b10000100101110: color_data = 12'b001000000000;
		14'b10000100101111: color_data = 12'b001000000000;
		14'b10000100110000: color_data = 12'b001000000000;
		14'b10000100110001: color_data = 12'b001000000000;
		14'b10000100110010: color_data = 12'b010000000000;
		14'b10000100110011: color_data = 12'b010000000000;
		14'b10000100110100: color_data = 12'b010000000000;
		14'b10000100110101: color_data = 12'b001000000000;
		14'b10000101000100: color_data = 12'b001000000000;
		14'b10000101000101: color_data = 12'b001000000000;
		14'b10000101000110: color_data = 12'b010000000000;
		14'b10000101000111: color_data = 12'b010000000000;
		14'b10000101001000: color_data = 12'b010000000000;
		14'b10000101001001: color_data = 12'b010000000000;
		14'b10000101001010: color_data = 12'b010000000000;
		14'b10000101001011: color_data = 12'b010000000000;
		14'b10000101001100: color_data = 12'b010000000000;
		14'b10000101001101: color_data = 12'b010000000000;
		14'b10000101001110: color_data = 12'b010000000000;
		14'b10000101001111: color_data = 12'b010000000000;
		14'b10000101010000: color_data = 12'b010000000000;
		14'b10000101010001: color_data = 12'b010000000000;
		14'b10000101010010: color_data = 12'b010000000000;
		14'b10000101010011: color_data = 12'b010000000000;
		14'b10000101010100: color_data = 12'b010000000000;
		14'b10000101010101: color_data = 12'b010000000000;
		14'b10000101010110: color_data = 12'b010000000000;
		14'b10000101010111: color_data = 12'b010000000000;
		14'b10000101011000: color_data = 12'b010000000000;
		14'b10000101011001: color_data = 12'b010000000000;
		14'b10000101011010: color_data = 12'b001000000000;
		14'b10000101110100: color_data = 12'b001000000000;
		14'b10000101110101: color_data = 12'b010000000000;
		14'b10000101110110: color_data = 12'b010000000000;
		14'b10000101110111: color_data = 12'b010000000000;
		14'b10000101111000: color_data = 12'b010000000000;
		14'b10000101111001: color_data = 12'b010000000000;
		14'b10000101111010: color_data = 12'b010000000000;
		14'b10000101111011: color_data = 12'b010000000000;
		14'b10000101111100: color_data = 12'b001000000000;
		14'b10000110100001: color_data = 12'b001000000000;
		14'b10000110100010: color_data = 12'b001000000000;
		14'b10000110101000: color_data = 12'b010000000000;
		14'b10000110101001: color_data = 12'b010000000000;
		14'b10000110101010: color_data = 12'b010000000000;
		14'b10000110101011: color_data = 12'b010000000000;
		14'b10000110101100: color_data = 12'b010000000000;
		14'b10000110101101: color_data = 12'b010000000000;
		14'b10000110101110: color_data = 12'b001000000000;
		14'b10000110101111: color_data = 12'b001000000000;
		14'b10000110110000: color_data = 12'b001000000000;
		14'b10000110110001: color_data = 12'b010000000000;
		14'b10000110110010: color_data = 12'b010000000000;
		14'b10000110110011: color_data = 12'b010000000000;
		14'b10000110110100: color_data = 12'b010000000000;
		14'b10000110110101: color_data = 12'b001000000000;
		14'b10000111000011: color_data = 12'b010000000000;
		14'b10000111000100: color_data = 12'b010000000000;
		14'b10000111000101: color_data = 12'b010000000000;
		14'b10000111000110: color_data = 12'b010000000000;
		14'b10000111000111: color_data = 12'b010000000000;
		14'b10000111001000: color_data = 12'b010000000000;
		14'b10000111001001: color_data = 12'b010000000000;
		14'b10000111001010: color_data = 12'b010000000000;
		14'b10000111001011: color_data = 12'b010000000000;
		14'b10000111001100: color_data = 12'b010000000000;
		14'b10000111001101: color_data = 12'b010000000000;
		14'b10000111001110: color_data = 12'b010000000000;
		14'b10000111001111: color_data = 12'b010000000000;
		14'b10000111010000: color_data = 12'b010000000000;
		14'b10000111010001: color_data = 12'b010000000000;
		14'b10000111010010: color_data = 12'b010000000000;
		14'b10000111010011: color_data = 12'b001000000000;
		14'b10000111010100: color_data = 12'b010000000000;
		14'b10000111010101: color_data = 12'b010000000000;
		14'b10000111010110: color_data = 12'b010000000000;
		14'b10000111010111: color_data = 12'b010000000000;
		14'b10000111011000: color_data = 12'b010000000000;
		14'b10000111011001: color_data = 12'b010000000000;
		14'b10000111011010: color_data = 12'b010000000000;
		14'b10000111110100: color_data = 12'b001000000000;
		14'b10000111110101: color_data = 12'b001000000000;
		14'b10000111110110: color_data = 12'b010000000000;
		14'b10000111110111: color_data = 12'b010000000000;
		14'b10000111111000: color_data = 12'b010000000000;
		14'b10000111111001: color_data = 12'b010000000000;
		14'b10000111111010: color_data = 12'b010000000000;
		14'b10000111111011: color_data = 12'b010000000000;
		14'b10000111111100: color_data = 12'b001000000000;
		14'b10001000100001: color_data = 12'b001000000000;
		14'b10001000100010: color_data = 12'b001000000000;
		14'b10001000101000: color_data = 12'b010000000000;
		14'b10001000101001: color_data = 12'b010000000000;
		14'b10001000101010: color_data = 12'b010000000000;
		14'b10001000101011: color_data = 12'b010000000000;
		14'b10001000101100: color_data = 12'b010000000000;
		14'b10001000101101: color_data = 12'b001000000000;
		14'b10001000101110: color_data = 12'b001000000000;
		14'b10001000101111: color_data = 12'b001000000000;
		14'b10001000110000: color_data = 12'b010000000000;
		14'b10001000110001: color_data = 12'b010000000000;
		14'b10001000110010: color_data = 12'b010000000000;
		14'b10001000110011: color_data = 12'b010000000000;
		14'b10001000110100: color_data = 12'b001000000000;
		14'b10001001000010: color_data = 12'b010000000000;
		14'b10001001000011: color_data = 12'b010000000000;
		14'b10001001000100: color_data = 12'b010000000000;
		14'b10001001000101: color_data = 12'b010000000000;
		14'b10001001000110: color_data = 12'b010000000000;
		14'b10001001000111: color_data = 12'b010000000000;
		14'b10001001001000: color_data = 12'b010000000000;
		14'b10001001001001: color_data = 12'b010000000000;
		14'b10001001001010: color_data = 12'b010000000000;
		14'b10001001001011: color_data = 12'b010000000000;
		14'b10001001001100: color_data = 12'b010000000000;
		14'b10001001001101: color_data = 12'b010000000000;
		14'b10001001001110: color_data = 12'b010000000000;
		14'b10001001001111: color_data = 12'b010000000000;
		14'b10001001010000: color_data = 12'b010000000000;
		14'b10001001010001: color_data = 12'b010000000000;
		14'b10001001010010: color_data = 12'b010000000000;
		14'b10001001010011: color_data = 12'b001000000000;
		14'b10001001010100: color_data = 12'b001000000000;
		14'b10001001010101: color_data = 12'b001000000000;
		14'b10001001010110: color_data = 12'b010000000000;
		14'b10001001010111: color_data = 12'b010000000000;
		14'b10001001011000: color_data = 12'b010000000000;
		14'b10001001011001: color_data = 12'b010000000000;
		14'b10001001011010: color_data = 12'b010000000000;
		14'b10001001011011: color_data = 12'b010000000000;
		14'b10001001110101: color_data = 12'b001000000000;
		14'b10001001110110: color_data = 12'b001000000000;
		14'b10001001110111: color_data = 12'b010000000000;
		14'b10001001111000: color_data = 12'b010000000000;
		14'b10001001111001: color_data = 12'b010000000000;
		14'b10001001111010: color_data = 12'b010000000000;
		14'b10001001111011: color_data = 12'b010000000000;
		14'b10001001111100: color_data = 12'b001000000000;
		14'b10001010100001: color_data = 12'b001000000000;
		14'b10001010100010: color_data = 12'b001000000000;
		14'b10001010101000: color_data = 12'b010000000000;
		14'b10001010101001: color_data = 12'b010000000000;
		14'b10001010101010: color_data = 12'b010000000000;
		14'b10001010101011: color_data = 12'b010000000000;
		14'b10001010101100: color_data = 12'b010000000000;
		14'b10001010101101: color_data = 12'b001000000000;
		14'b10001010101110: color_data = 12'b001000000000;
		14'b10001010101111: color_data = 12'b001000000000;
		14'b10001010110000: color_data = 12'b010000000000;
		14'b10001010110001: color_data = 12'b010000000000;
		14'b10001010110010: color_data = 12'b010000000000;
		14'b10001010110011: color_data = 12'b010000000000;
		14'b10001010110100: color_data = 12'b001000000000;
		14'b10001011000001: color_data = 12'b001000000000;
		14'b10001011000010: color_data = 12'b010000000000;
		14'b10001011000011: color_data = 12'b001000000000;
		14'b10001011000100: color_data = 12'b001000000000;
		14'b10001011000101: color_data = 12'b001000000000;
		14'b10001011000110: color_data = 12'b001000000000;
		14'b10001011000111: color_data = 12'b010000000000;
		14'b10001011001000: color_data = 12'b010000000000;
		14'b10001011001001: color_data = 12'b010000000000;
		14'b10001011001010: color_data = 12'b010000000000;
		14'b10001011001011: color_data = 12'b001000000000;
		14'b10001011001100: color_data = 12'b001000000000;
		14'b10001011001111: color_data = 12'b001000000000;
		14'b10001011010000: color_data = 12'b001000000000;
		14'b10001011010001: color_data = 12'b010000000000;
		14'b10001011010010: color_data = 12'b010000000000;
		14'b10001011010011: color_data = 12'b010000000000;
		14'b10001011010111: color_data = 12'b001000000000;
		14'b10001011011000: color_data = 12'b010000000000;
		14'b10001011011001: color_data = 12'b010000000000;
		14'b10001011011010: color_data = 12'b010000000000;
		14'b10001011011011: color_data = 12'b010000000000;
		14'b10001011011100: color_data = 12'b010000000000;
		14'b10001011110110: color_data = 12'b001000000000;
		14'b10001011110111: color_data = 12'b010000000000;
		14'b10001011111000: color_data = 12'b010000000000;
		14'b10001011111001: color_data = 12'b010000000000;
		14'b10001011111010: color_data = 12'b010000000000;
		14'b10001011111011: color_data = 12'b010000000000;
		14'b10001011111100: color_data = 12'b001000000000;
		14'b10001100100001: color_data = 12'b001000000000;
		14'b10001100100010: color_data = 12'b001000000000;
		14'b10001100100011: color_data = 12'b001000000000;
		14'b10001100101000: color_data = 12'b010000000000;
		14'b10001100101001: color_data = 12'b010000000000;
		14'b10001100101010: color_data = 12'b010000000000;
		14'b10001100101011: color_data = 12'b010000000000;
		14'b10001100101100: color_data = 12'b001000000000;
		14'b10001100101101: color_data = 12'b001000000000;
		14'b10001100101110: color_data = 12'b001000000000;
		14'b10001100101111: color_data = 12'b001000000000;
		14'b10001100110000: color_data = 12'b010000000000;
		14'b10001100110001: color_data = 12'b010000000000;
		14'b10001100110010: color_data = 12'b010000000000;
		14'b10001100110011: color_data = 12'b001000000000;
		14'b10001101000001: color_data = 12'b001000000000;
		14'b10001101000010: color_data = 12'b001000000000;
		14'b10001101000011: color_data = 12'b001000000000;
		14'b10001101000100: color_data = 12'b001000000000;
		14'b10001101000101: color_data = 12'b001000000000;
		14'b10001101000110: color_data = 12'b001000000000;
		14'b10001101000111: color_data = 12'b010000000000;
		14'b10001101001000: color_data = 12'b010000000000;
		14'b10001101001001: color_data = 12'b010000000000;
		14'b10001101001010: color_data = 12'b001000000000;
		14'b10001101010001: color_data = 12'b010000000000;
		14'b10001101010010: color_data = 12'b010000000000;
		14'b10001101010011: color_data = 12'b010000000000;
		14'b10001101011000: color_data = 12'b001000000000;
		14'b10001101011001: color_data = 12'b001000000000;
		14'b10001101011010: color_data = 12'b010000000000;
		14'b10001101011011: color_data = 12'b010000000000;
		14'b10001101011100: color_data = 12'b010000000000;
		14'b10001101011101: color_data = 12'b001000000000;
		14'b10001101110110: color_data = 12'b001000000000;
		14'b10001101110111: color_data = 12'b001000000000;
		14'b10001101111000: color_data = 12'b010000000000;
		14'b10001101111001: color_data = 12'b010000000000;
		14'b10001101111010: color_data = 12'b010000000000;
		14'b10001101111011: color_data = 12'b010000000000;
		14'b10001101111100: color_data = 12'b001000000000;
		14'b10001110100001: color_data = 12'b001000000000;
		14'b10001110100010: color_data = 12'b001000000000;
		14'b10001110101000: color_data = 12'b010000000000;
		14'b10001110101001: color_data = 12'b010000000000;
		14'b10001110101010: color_data = 12'b010000000000;
		14'b10001110101011: color_data = 12'b001000000000;
		14'b10001110101100: color_data = 12'b001000000000;
		14'b10001110101101: color_data = 12'b001000000000;
		14'b10001110101110: color_data = 12'b001000000000;
		14'b10001110101111: color_data = 12'b001000000000;
		14'b10001110110000: color_data = 12'b010000000000;
		14'b10001110110001: color_data = 12'b010000000000;
		14'b10001110110010: color_data = 12'b010000000000;
		14'b10001110110011: color_data = 12'b001000000000;
		14'b10001111000000: color_data = 12'b001000000000;
		14'b10001111000100: color_data = 12'b001000000000;
		14'b10001111000101: color_data = 12'b001000000000;
		14'b10001111000110: color_data = 12'b010000000000;
		14'b10001111000111: color_data = 12'b010000000000;
		14'b10001111001000: color_data = 12'b010000000000;
		14'b10001111001001: color_data = 12'b010000000000;
		14'b10001111010001: color_data = 12'b010000000000;
		14'b10001111010010: color_data = 12'b010000000000;
		14'b10001111010011: color_data = 12'b010000000000;
		14'b10001111010100: color_data = 12'b010000000000;
		14'b10001111011010: color_data = 12'b010000000000;
		14'b10001111011011: color_data = 12'b010000000000;
		14'b10001111011100: color_data = 12'b010000000000;
		14'b10001111011101: color_data = 12'b010000000000;
		14'b10001111011110: color_data = 12'b001000000000;
		14'b10001111110111: color_data = 12'b001000000000;
		14'b10001111111000: color_data = 12'b010000000000;
		14'b10001111111001: color_data = 12'b010000000000;
		14'b10001111111010: color_data = 12'b010000000000;
		14'b10001111111011: color_data = 12'b010000000000;
		14'b10001111111100: color_data = 12'b001000000000;
		14'b10010000100000: color_data = 12'b001000000000;
		14'b10010000100111: color_data = 12'b001000000000;
		14'b10010000101000: color_data = 12'b010000000000;
		14'b10010000101001: color_data = 12'b010000000000;
		14'b10010000101010: color_data = 12'b010000000000;
		14'b10010000101011: color_data = 12'b001000000000;
		14'b10010000101100: color_data = 12'b001000000000;
		14'b10010000101101: color_data = 12'b001000000000;
		14'b10010000101110: color_data = 12'b001000000000;
		14'b10010000101111: color_data = 12'b001000000000;
		14'b10010000110000: color_data = 12'b010000000000;
		14'b10010000110001: color_data = 12'b010000000000;
		14'b10010000110010: color_data = 12'b010000000000;
		14'b10010000110011: color_data = 12'b001000000000;
		14'b10010000111111: color_data = 12'b001000000000;
		14'b10010001000000: color_data = 12'b001000000000;
		14'b10010001000100: color_data = 12'b001000000000;
		14'b10010001000101: color_data = 12'b001000000000;
		14'b10010001000110: color_data = 12'b010000000000;
		14'b10010001000111: color_data = 12'b010000000000;
		14'b10010001001000: color_data = 12'b010000000000;
		14'b10010001010000: color_data = 12'b001000000000;
		14'b10010001010001: color_data = 12'b010000000000;
		14'b10010001010010: color_data = 12'b010000000000;
		14'b10010001010011: color_data = 12'b010000000000;
		14'b10010001010100: color_data = 12'b010000000000;
		14'b10010001010101: color_data = 12'b010000000000;
		14'b10010001011011: color_data = 12'b010000000000;
		14'b10010001011100: color_data = 12'b010000000000;
		14'b10010001011101: color_data = 12'b010000000000;
		14'b10010001011110: color_data = 12'b001000000000;
		14'b10010001011111: color_data = 12'b001000000000;
		14'b10010001111000: color_data = 12'b010000000000;
		14'b10010001111001: color_data = 12'b010000000000;
		14'b10010001111010: color_data = 12'b010000000000;
		14'b10010001111011: color_data = 12'b010000000000;
		14'b10010001111100: color_data = 12'b001000000000;
		14'b10010010100111: color_data = 12'b001000000000;
		14'b10010010101000: color_data = 12'b010000000000;
		14'b10010010101001: color_data = 12'b001000000000;
		14'b10010010101010: color_data = 12'b001000000000;
		14'b10010010101011: color_data = 12'b001000000000;
		14'b10010010101100: color_data = 12'b001000000000;
		14'b10010010101101: color_data = 12'b001000000000;
		14'b10010010101110: color_data = 12'b001000000000;
		14'b10010010101111: color_data = 12'b010000000000;
		14'b10010010110000: color_data = 12'b010000000000;
		14'b10010010110001: color_data = 12'b010000000000;
		14'b10010010110010: color_data = 12'b001000000000;
		14'b10010010111111: color_data = 12'b001000000000;
		14'b10010011000100: color_data = 12'b001000000000;
		14'b10010011000101: color_data = 12'b010000000000;
		14'b10010011000110: color_data = 12'b010000000000;
		14'b10010011000111: color_data = 12'b010000000000;
		14'b10010011001111: color_data = 12'b001000000000;
		14'b10010011010000: color_data = 12'b001000000000;
		14'b10010011010001: color_data = 12'b010000000000;
		14'b10010011010010: color_data = 12'b010000000000;
		14'b10010011010011: color_data = 12'b010000000000;
		14'b10010011010100: color_data = 12'b010000000000;
		14'b10010011010101: color_data = 12'b010000000000;
		14'b10010011010110: color_data = 12'b001000000000;
		14'b10010011010111: color_data = 12'b001000000000;
		14'b10010011011100: color_data = 12'b010000000000;
		14'b10010011011101: color_data = 12'b010000000000;
		14'b10010011011110: color_data = 12'b001000000000;
		14'b10010011011111: color_data = 12'b001000000000;
		14'b10010011111000: color_data = 12'b001000000000;
		14'b10010011111001: color_data = 12'b010000000000;
		14'b10010011111010: color_data = 12'b010000000000;
		14'b10010011111011: color_data = 12'b010000000000;
		14'b10010011111100: color_data = 12'b010000000000;
		14'b10010011111101: color_data = 12'b001000000000;
		14'b10010100100110: color_data = 12'b001000000000;
		14'b10010100100111: color_data = 12'b010000000000;
		14'b10010100101000: color_data = 12'b001000000000;
		14'b10010100101001: color_data = 12'b001000000000;
		14'b10010100101010: color_data = 12'b001000000000;
		14'b10010100101011: color_data = 12'b001000000000;
		14'b10010100101100: color_data = 12'b001000000000;
		14'b10010100101101: color_data = 12'b001000000000;
		14'b10010100101110: color_data = 12'b001000000000;
		14'b10010100101111: color_data = 12'b010000000000;
		14'b10010100110000: color_data = 12'b010000000000;
		14'b10010100110001: color_data = 12'b010000000000;
		14'b10010100110010: color_data = 12'b001000000000;
		14'b10010101000011: color_data = 12'b001000000000;
		14'b10010101000100: color_data = 12'b010000000000;
		14'b10010101000101: color_data = 12'b010000000000;
		14'b10010101000110: color_data = 12'b010000000000;
		14'b10010101000111: color_data = 12'b001000000000;
		14'b10010101001011: color_data = 12'b001000000000;
		14'b10010101001100: color_data = 12'b001000000000;
		14'b10010101001101: color_data = 12'b001000000000;
		14'b10010101001110: color_data = 12'b001000000000;
		14'b10010101001111: color_data = 12'b010000000000;
		14'b10010101010000: color_data = 12'b010000000000;
		14'b10010101010001: color_data = 12'b010000000000;
		14'b10010101010010: color_data = 12'b010000000000;
		14'b10010101010011: color_data = 12'b010000000000;
		14'b10010101010100: color_data = 12'b010000000000;
		14'b10010101010101: color_data = 12'b010000000000;
		14'b10010101010110: color_data = 12'b010000000000;
		14'b10010101010111: color_data = 12'b010000000000;
		14'b10010101011000: color_data = 12'b001000000000;
		14'b10010101011101: color_data = 12'b010000000000;
		14'b10010101011110: color_data = 12'b001000000000;
		14'b10010101011111: color_data = 12'b001000000000;
		14'b10010101100000: color_data = 12'b001000000000;
		14'b10010101111001: color_data = 12'b010000000000;
		14'b10010101111010: color_data = 12'b010000000000;
		14'b10010101111011: color_data = 12'b010000000000;
		14'b10010101111100: color_data = 12'b010000000000;
		14'b10010101111101: color_data = 12'b001000000000;
		14'b10010110100010: color_data = 12'b001000000000;
		14'b10010110100110: color_data = 12'b001000000000;
		14'b10010110100111: color_data = 12'b001000000000;
		14'b10010110101000: color_data = 12'b001000000000;
		14'b10010110101001: color_data = 12'b001000000000;
		14'b10010110101010: color_data = 12'b010000000000;
		14'b10010110101011: color_data = 12'b010000000000;
		14'b10010110101100: color_data = 12'b001000000000;
		14'b10010110101101: color_data = 12'b001000000000;
		14'b10010110101110: color_data = 12'b001000000000;
		14'b10010110101111: color_data = 12'b010000000000;
		14'b10010110110000: color_data = 12'b010000000000;
		14'b10010110110001: color_data = 12'b001000000000;
		14'b10010110110010: color_data = 12'b001000000000;
		14'b10010111000010: color_data = 12'b001000000000;
		14'b10010111000101: color_data = 12'b001000000000;
		14'b10010111000110: color_data = 12'b001000000000;
		14'b10010111000111: color_data = 12'b001000000000;
		14'b10010111001000: color_data = 12'b001000000000;
		14'b10010111001001: color_data = 12'b001000000000;
		14'b10010111001010: color_data = 12'b010000000000;
		14'b10010111001011: color_data = 12'b010000000000;
		14'b10010111001100: color_data = 12'b010000000000;
		14'b10010111001101: color_data = 12'b010000000000;
		14'b10010111001110: color_data = 12'b010000000000;
		14'b10010111001111: color_data = 12'b010000000000;
		14'b10010111010000: color_data = 12'b010000000000;
		14'b10010111010001: color_data = 12'b010000000000;
		14'b10010111010010: color_data = 12'b010000000000;
		14'b10010111010011: color_data = 12'b010000000000;
		14'b10010111010100: color_data = 12'b010000000000;
		14'b10010111010101: color_data = 12'b010000000000;
		14'b10010111010110: color_data = 12'b010000000000;
		14'b10010111010111: color_data = 12'b010000000000;
		14'b10010111011000: color_data = 12'b010000000000;
		14'b10010111011001: color_data = 12'b001000000000;
		14'b10010111011110: color_data = 12'b001000000000;
		14'b10010111011111: color_data = 12'b001000000000;
		14'b10010111100001: color_data = 12'b001000000000;
		14'b10010111111001: color_data = 12'b001000000000;
		14'b10010111111010: color_data = 12'b010000000000;
		14'b10010111111011: color_data = 12'b010000000000;
		14'b10010111111100: color_data = 12'b010000000000;
		14'b10010111111101: color_data = 12'b010000000000;
		14'b10010111111110: color_data = 12'b001000000000;
		14'b10011000011110: color_data = 12'b001000000000;
		14'b10011000100001: color_data = 12'b001000000000;
		14'b10011000100010: color_data = 12'b001000000000;
		14'b10011000100101: color_data = 12'b001000000000;
		14'b10011000100110: color_data = 12'b010000000000;
		14'b10011000100111: color_data = 12'b010000000000;
		14'b10011000101000: color_data = 12'b010000000000;
		14'b10011000101001: color_data = 12'b010000000000;
		14'b10011000101010: color_data = 12'b010000000000;
		14'b10011000101011: color_data = 12'b001000000000;
		14'b10011000101100: color_data = 12'b001000000000;
		14'b10011000101101: color_data = 12'b001000000000;
		14'b10011000101110: color_data = 12'b010000000000;
		14'b10011000101111: color_data = 12'b010000000000;
		14'b10011000110000: color_data = 12'b010000000000;
		14'b10011000110001: color_data = 12'b001000000000;
		14'b10011000110010: color_data = 12'b001000000000;
		14'b10011001000001: color_data = 12'b001000000000;
		14'b10011001000010: color_data = 12'b001000000000;
		14'b10011001000101: color_data = 12'b001000000000;
		14'b10011001000110: color_data = 12'b001000000000;
		14'b10011001000111: color_data = 12'b001000000000;
		14'b10011001001000: color_data = 12'b010000000000;
		14'b10011001001001: color_data = 12'b010000000000;
		14'b10011001001010: color_data = 12'b010000000000;
		14'b10011001001011: color_data = 12'b010000000000;
		14'b10011001001100: color_data = 12'b010000000000;
		14'b10011001001101: color_data = 12'b010000000000;
		14'b10011001001110: color_data = 12'b010000000000;
		14'b10011001001111: color_data = 12'b010000000000;
		14'b10011001010000: color_data = 12'b010000000000;
		14'b10011001010001: color_data = 12'b010000000000;
		14'b10011001010010: color_data = 12'b010000000000;
		14'b10011001010011: color_data = 12'b010000000000;
		14'b10011001010100: color_data = 12'b010000000000;
		14'b10011001010101: color_data = 12'b010000000000;
		14'b10011001010110: color_data = 12'b010000000000;
		14'b10011001010111: color_data = 12'b010000000000;
		14'b10011001011000: color_data = 12'b010000000000;
		14'b10011001011001: color_data = 12'b010000000000;
		14'b10011001011010: color_data = 12'b001000000000;
		14'b10011001011110: color_data = 12'b001000000000;
		14'b10011001011111: color_data = 12'b001000000000;
		14'b10011001100001: color_data = 12'b001000000000;
		14'b10011001111001: color_data = 12'b001000000000;
		14'b10011001111010: color_data = 12'b001000000000;
		14'b10011001111011: color_data = 12'b010000000000;
		14'b10011001111100: color_data = 12'b010000000000;
		14'b10011001111101: color_data = 12'b010000000000;
		14'b10011001111110: color_data = 12'b001000000000;
		14'b10011010011110: color_data = 12'b001000000000;
		14'b10011010100000: color_data = 12'b001000000000;
		14'b10011010100001: color_data = 12'b001000000000;
		14'b10011010100100: color_data = 12'b001000000000;
		14'b10011010100101: color_data = 12'b010000000000;
		14'b10011010100110: color_data = 12'b010000000000;
		14'b10011010100111: color_data = 12'b010000000000;
		14'b10011010101000: color_data = 12'b010000000000;
		14'b10011010101001: color_data = 12'b010000000000;
		14'b10011010101010: color_data = 12'b010000000000;
		14'b10011010101011: color_data = 12'b001000000000;
		14'b10011010101100: color_data = 12'b001000000000;
		14'b10011010101101: color_data = 12'b001000000000;
		14'b10011010101110: color_data = 12'b010000000000;
		14'b10011010101111: color_data = 12'b010000000000;
		14'b10011010110000: color_data = 12'b001000000000;
		14'b10011010110001: color_data = 12'b001000000000;
		14'b10011010110010: color_data = 12'b001000000000;
		14'b10011011000001: color_data = 12'b001000000000;
		14'b10011011000101: color_data = 12'b001000000000;
		14'b10011011000110: color_data = 12'b001000000000;
		14'b10011011000111: color_data = 12'b010000000000;
		14'b10011011001000: color_data = 12'b010000000000;
		14'b10011011001001: color_data = 12'b010000000000;
		14'b10011011001010: color_data = 12'b010000000000;
		14'b10011011001011: color_data = 12'b010000000000;
		14'b10011011001100: color_data = 12'b001000000000;
		14'b10011011001101: color_data = 12'b001000000000;
		14'b10011011001110: color_data = 12'b010000000000;
		14'b10011011001111: color_data = 12'b010000000000;
		14'b10011011010000: color_data = 12'b010000000000;
		14'b10011011010001: color_data = 12'b010000000000;
		14'b10011011010010: color_data = 12'b010000000000;
		14'b10011011010011: color_data = 12'b010000000000;
		14'b10011011010100: color_data = 12'b010000000000;
		14'b10011011010101: color_data = 12'b010000000000;
		14'b10011011010110: color_data = 12'b010000000000;
		14'b10011011010111: color_data = 12'b010000000000;
		14'b10011011011000: color_data = 12'b010000000000;
		14'b10011011011001: color_data = 12'b010000000000;
		14'b10011011011010: color_data = 12'b010000000000;
		14'b10011011011011: color_data = 12'b001000000000;
		14'b10011011011100: color_data = 12'b001000000000;
		14'b10011011011110: color_data = 12'b001000000000;
		14'b10011011011111: color_data = 12'b001000000000;
		14'b10011011111010: color_data = 12'b001000000000;
		14'b10011011111011: color_data = 12'b010000000000;
		14'b10011011111100: color_data = 12'b010000000000;
		14'b10011011111101: color_data = 12'b010000000000;
		14'b10011011111110: color_data = 12'b001000000000;
		14'b10011011111111: color_data = 12'b001000000000;
		14'b10011100000000: color_data = 12'b001000000000;
		14'b10011100100000: color_data = 12'b001000000000;
		14'b10011100100011: color_data = 12'b001000000000;
		14'b10011100100100: color_data = 12'b010000000000;
		14'b10011100100101: color_data = 12'b010000000000;
		14'b10011100100110: color_data = 12'b010000000000;
		14'b10011100100111: color_data = 12'b010000000000;
		14'b10011100101000: color_data = 12'b010000000000;
		14'b10011100101001: color_data = 12'b010000000000;
		14'b10011100101010: color_data = 12'b010000000000;
		14'b10011100101011: color_data = 12'b010000000000;
		14'b10011100101100: color_data = 12'b001000000000;
		14'b10011100101101: color_data = 12'b001000000000;
		14'b10011100101110: color_data = 12'b010000000000;
		14'b10011100101111: color_data = 12'b010000000000;
		14'b10011100110000: color_data = 12'b001000000000;
		14'b10011100110001: color_data = 12'b001000000000;
		14'b10011100110010: color_data = 12'b001000000000;
		14'b10011101000101: color_data = 12'b001000000000;
		14'b10011101000110: color_data = 12'b010000000000;
		14'b10011101000111: color_data = 12'b010000000000;
		14'b10011101001000: color_data = 12'b010000000000;
		14'b10011101001001: color_data = 12'b010000000000;
		14'b10011101001010: color_data = 12'b001000000000;
		14'b10011101001011: color_data = 12'b001000000000;
		14'b10011101001100: color_data = 12'b001000000000;
		14'b10011101001101: color_data = 12'b001000000000;
		14'b10011101001110: color_data = 12'b010000000000;
		14'b10011101001111: color_data = 12'b010000000000;
		14'b10011101010000: color_data = 12'b010000000000;
		14'b10011101010001: color_data = 12'b010000000000;
		14'b10011101010010: color_data = 12'b010000000000;
		14'b10011101010011: color_data = 12'b010000000000;
		14'b10011101010100: color_data = 12'b001000000000;
		14'b10011101010101: color_data = 12'b001000000000;
		14'b10011101010110: color_data = 12'b010000000000;
		14'b10011101010111: color_data = 12'b010000000000;
		14'b10011101011000: color_data = 12'b010000000000;
		14'b10011101011001: color_data = 12'b010000000000;
		14'b10011101011010: color_data = 12'b010000000000;
		14'b10011101011011: color_data = 12'b010000000000;
		14'b10011101011100: color_data = 12'b010000000000;
		14'b10011101011111: color_data = 12'b010000000000;
		14'b10011101100000: color_data = 12'b001000000000;
		14'b10011101111010: color_data = 12'b001000000000;
		14'b10011101111011: color_data = 12'b001000000000;
		14'b10011101111100: color_data = 12'b010000000000;
		14'b10011101111101: color_data = 12'b010000000000;
		14'b10011101111110: color_data = 12'b010000000000;
		14'b10011101111111: color_data = 12'b001000000000;
		14'b10011110000000: color_data = 12'b001000000000;
		14'b10011110100011: color_data = 12'b010000000000;
		14'b10011110100100: color_data = 12'b010000000000;
		14'b10011110100101: color_data = 12'b010000000000;
		14'b10011110100110: color_data = 12'b010000000000;
		14'b10011110100111: color_data = 12'b010000000000;
		14'b10011110101000: color_data = 12'b010000000000;
		14'b10011110101001: color_data = 12'b010000000000;
		14'b10011110101010: color_data = 12'b010000000000;
		14'b10011110101011: color_data = 12'b010000000000;
		14'b10011110101100: color_data = 12'b001000000000;
		14'b10011110101101: color_data = 12'b001000000000;
		14'b10011110101110: color_data = 12'b010000000000;
		14'b10011110101111: color_data = 12'b001000000000;
		14'b10011110110000: color_data = 12'b001000000000;
		14'b10011110110001: color_data = 12'b010000000000;
		14'b10011110110010: color_data = 12'b001000000000;
		14'b10011111000100: color_data = 12'b001000000000;
		14'b10011111000101: color_data = 12'b001000000000;
		14'b10011111000110: color_data = 12'b001000000000;
		14'b10011111000111: color_data = 12'b001000000000;
		14'b10011111001000: color_data = 12'b001000000000;
		14'b10011111001001: color_data = 12'b001000000000;
		14'b10011111001011: color_data = 12'b001000000000;
		14'b10011111001100: color_data = 12'b001000000000;
		14'b10011111001101: color_data = 12'b010000000000;
		14'b10011111001110: color_data = 12'b010000000000;
		14'b10011111001111: color_data = 12'b010000000000;
		14'b10011111010000: color_data = 12'b010000000000;
		14'b10011111010001: color_data = 12'b010000000000;
		14'b10011111010010: color_data = 12'b001000000000;
		14'b10011111010011: color_data = 12'b001000000000;
		14'b10011111010110: color_data = 12'b001000000000;
		14'b10011111010111: color_data = 12'b010000000000;
		14'b10011111011000: color_data = 12'b001000000000;
		14'b10011111011001: color_data = 12'b010000000000;
		14'b10011111011010: color_data = 12'b010000000000;
		14'b10011111011011: color_data = 12'b010000000000;
		14'b10011111011100: color_data = 12'b010000000000;
		14'b10011111011101: color_data = 12'b001000000000;
		14'b10011111011110: color_data = 12'b001000000000;
		14'b10011111011111: color_data = 12'b001000000000;
		14'b10011111100000: color_data = 12'b010000000000;
		14'b10011111100001: color_data = 12'b001000000000;
		14'b10011111111011: color_data = 12'b001000000000;
		14'b10011111111100: color_data = 12'b010000000000;
		14'b10011111111101: color_data = 12'b010000000000;
		14'b10011111111110: color_data = 12'b010000000000;
		14'b10011111111111: color_data = 12'b001000000000;
		14'b10100000000000: color_data = 12'b001000000000;
		14'b10100000010011: color_data = 12'b001000000000;
		14'b10100000010100: color_data = 12'b001000000000;
		14'b10100000100010: color_data = 12'b001000000000;
		14'b10100000100011: color_data = 12'b010000000000;
		14'b10100000100100: color_data = 12'b010000000000;
		14'b10100000100101: color_data = 12'b010000000000;
		14'b10100000100110: color_data = 12'b010000000000;
		14'b10100000100111: color_data = 12'b010000000000;
		14'b10100000101000: color_data = 12'b010000000000;
		14'b10100000101001: color_data = 12'b010000000000;
		14'b10100000101010: color_data = 12'b010000000000;
		14'b10100000101011: color_data = 12'b010000000000;
		14'b10100000101100: color_data = 12'b001000000000;
		14'b10100000101101: color_data = 12'b001000000000;
		14'b10100000101110: color_data = 12'b001000000000;
		14'b10100000101111: color_data = 12'b001000000000;
		14'b10100000110000: color_data = 12'b001000000000;
		14'b10100000110001: color_data = 12'b010000000000;
		14'b10100000110010: color_data = 12'b001000000000;
		14'b10100001000011: color_data = 12'b001000000000;
		14'b10100001000100: color_data = 12'b001000000000;
		14'b10100001001011: color_data = 12'b001000000000;
		14'b10100001001100: color_data = 12'b010000000000;
		14'b10100001001101: color_data = 12'b010000000000;
		14'b10100001001110: color_data = 12'b010000000000;
		14'b10100001001111: color_data = 12'b010000000000;
		14'b10100001010000: color_data = 12'b001000000000;
		14'b10100001010001: color_data = 12'b001000000000;
		14'b10100001010110: color_data = 12'b010000000000;
		14'b10100001010111: color_data = 12'b001000000000;
		14'b10100001011001: color_data = 12'b001000000000;
		14'b10100001011010: color_data = 12'b010000000000;
		14'b10100001011011: color_data = 12'b010000000000;
		14'b10100001011100: color_data = 12'b010000000000;
		14'b10100001011101: color_data = 12'b010000000000;
		14'b10100001011110: color_data = 12'b001000000000;
		14'b10100001011111: color_data = 12'b001000000000;
		14'b10100001100000: color_data = 12'b010000000000;
		14'b10100001100001: color_data = 12'b010000000000;
		14'b10100001111011: color_data = 12'b001000000000;
		14'b10100001111100: color_data = 12'b001000000000;
		14'b10100001111101: color_data = 12'b010000000000;
		14'b10100001111110: color_data = 12'b010000000000;
		14'b10100001111111: color_data = 12'b010000000000;
		14'b10100010000000: color_data = 12'b001000000000;
		14'b10100010010110: color_data = 12'b001000000000;
		14'b10100010011110: color_data = 12'b001000000000;
		14'b10100010100010: color_data = 12'b001000000000;
		14'b10100010100011: color_data = 12'b010000000000;
		14'b10100010100100: color_data = 12'b010000000000;
		14'b10100010100101: color_data = 12'b010000000000;
		14'b10100010100110: color_data = 12'b010000000000;
		14'b10100010100111: color_data = 12'b010000000000;
		14'b10100010101000: color_data = 12'b010000000000;
		14'b10100010101001: color_data = 12'b010000000000;
		14'b10100010101010: color_data = 12'b010000000000;
		14'b10100010101011: color_data = 12'b001000000000;
		14'b10100010101100: color_data = 12'b001000000000;
		14'b10100010101101: color_data = 12'b001000000000;
		14'b10100010101110: color_data = 12'b001000000000;
		14'b10100010101111: color_data = 12'b001000000000;
		14'b10100010110000: color_data = 12'b010000000000;
		14'b10100010110001: color_data = 12'b010000000000;
		14'b10100010110010: color_data = 12'b010000000000;
		14'b10100011001001: color_data = 12'b001000000000;
		14'b10100011001010: color_data = 12'b001000000000;
		14'b10100011001011: color_data = 12'b010000000000;
		14'b10100011001100: color_data = 12'b010000000000;
		14'b10100011001101: color_data = 12'b010000000000;
		14'b10100011001110: color_data = 12'b010000000000;
		14'b10100011001111: color_data = 12'b001000000000;
		14'b10100011010100: color_data = 12'b001000000000;
		14'b10100011010101: color_data = 12'b001000000000;
		14'b10100011010110: color_data = 12'b010000000000;
		14'b10100011010111: color_data = 12'b010000000000;
		14'b10100011011010: color_data = 12'b001000000000;
		14'b10100011011011: color_data = 12'b010000000000;
		14'b10100011011100: color_data = 12'b010000000000;
		14'b10100011011101: color_data = 12'b010000000000;
		14'b10100011011110: color_data = 12'b010000000000;
		14'b10100011011111: color_data = 12'b001000000000;
		14'b10100011100000: color_data = 12'b001000000000;
		14'b10100011100001: color_data = 12'b010000000000;
		14'b10100011100010: color_data = 12'b001000000000;
		14'b10100011111011: color_data = 12'b001000000000;
		14'b10100011111100: color_data = 12'b001000000000;
		14'b10100011111101: color_data = 12'b010000000000;
		14'b10100011111110: color_data = 12'b010000000000;
		14'b10100011111111: color_data = 12'b010000000000;
		14'b10100100000000: color_data = 12'b001000000000;
		14'b10100100000001: color_data = 12'b001000000000;
		14'b10100100011000: color_data = 12'b001000000000;
		14'b10100100011110: color_data = 12'b001000000000;
		14'b10100100100010: color_data = 12'b001000000000;
		14'b10100100100011: color_data = 12'b010000000000;
		14'b10100100100100: color_data = 12'b010000000000;
		14'b10100100100101: color_data = 12'b010000000000;
		14'b10100100100110: color_data = 12'b010000000000;
		14'b10100100100111: color_data = 12'b010000000000;
		14'b10100100101000: color_data = 12'b010000000000;
		14'b10100100101001: color_data = 12'b010000000000;
		14'b10100100101010: color_data = 12'b001000000000;
		14'b10100100101011: color_data = 12'b001000000000;
		14'b10100100101100: color_data = 12'b001000000000;
		14'b10100100101101: color_data = 12'b001000000000;
		14'b10100100101110: color_data = 12'b001000000000;
		14'b10100100101111: color_data = 12'b010000000000;
		14'b10100100110000: color_data = 12'b010000000000;
		14'b10100100110001: color_data = 12'b010000000000;
		14'b10100100110010: color_data = 12'b001000000000;
		14'b10100101001000: color_data = 12'b001000000000;
		14'b10100101001001: color_data = 12'b001000000000;
		14'b10100101001010: color_data = 12'b010000000000;
		14'b10100101001011: color_data = 12'b010000000000;
		14'b10100101001100: color_data = 12'b010000000000;
		14'b10100101001101: color_data = 12'b010000000000;
		14'b10100101001110: color_data = 12'b001000000000;
		14'b10100101001111: color_data = 12'b001000000000;
		14'b10100101010000: color_data = 12'b001000000000;
		14'b10100101010001: color_data = 12'b001000000000;
		14'b10100101010010: color_data = 12'b001000000000;
		14'b10100101010011: color_data = 12'b010000000000;
		14'b10100101010100: color_data = 12'b010000000000;
		14'b10100101010101: color_data = 12'b010000000000;
		14'b10100101010110: color_data = 12'b010000000000;
		14'b10100101010111: color_data = 12'b010000000000;
		14'b10100101011000: color_data = 12'b001000000000;
		14'b10100101011010: color_data = 12'b001000000000;
		14'b10100101011011: color_data = 12'b010000000000;
		14'b10100101011100: color_data = 12'b010000000000;
		14'b10100101011101: color_data = 12'b010000000000;
		14'b10100101011110: color_data = 12'b010000000000;
		14'b10100101011111: color_data = 12'b010000000000;
		14'b10100101100000: color_data = 12'b001000000000;
		14'b10100101100001: color_data = 12'b001000000000;
		14'b10100101100010: color_data = 12'b001000000000;
		14'b10100101111100: color_data = 12'b001000000000;
		14'b10100101111101: color_data = 12'b010000000000;
		14'b10100101111110: color_data = 12'b010000000000;
		14'b10100101111111: color_data = 12'b010000000000;
		14'b10100110000000: color_data = 12'b001000000000;
		14'b10100110000001: color_data = 12'b001000000000;
		14'b10100110011000: color_data = 12'b001000000000;
		14'b10100110011001: color_data = 12'b001000000000;
		14'b10100110011110: color_data = 12'b001000000000;
		14'b10100110100010: color_data = 12'b001000000000;
		14'b10100110100011: color_data = 12'b010000000000;
		14'b10100110100100: color_data = 12'b010000000000;
		14'b10100110100101: color_data = 12'b010000000000;
		14'b10100110100110: color_data = 12'b010000000000;
		14'b10100110100111: color_data = 12'b010000000000;
		14'b10100110101000: color_data = 12'b001000000000;
		14'b10100110101001: color_data = 12'b001000000000;
		14'b10100110101010: color_data = 12'b001000000000;
		14'b10100110101011: color_data = 12'b001000000000;
		14'b10100110101100: color_data = 12'b001000000000;
		14'b10100110101101: color_data = 12'b010000000000;
		14'b10100110101110: color_data = 12'b010000000000;
		14'b10100110101111: color_data = 12'b010000000000;
		14'b10100110110000: color_data = 12'b010000000000;
		14'b10100110110001: color_data = 12'b010000000000;
		14'b10100110110010: color_data = 12'b001000000000;
		14'b10100111000110: color_data = 12'b001000000000;
		14'b10100111001000: color_data = 12'b010000000000;
		14'b10100111001001: color_data = 12'b010000000000;
		14'b10100111001010: color_data = 12'b010000000000;
		14'b10100111001011: color_data = 12'b010000000000;
		14'b10100111001100: color_data = 12'b010000000000;
		14'b10100111001101: color_data = 12'b010000000000;
		14'b10100111001110: color_data = 12'b010000000000;
		14'b10100111001111: color_data = 12'b010000000000;
		14'b10100111010000: color_data = 12'b010000000000;
		14'b10100111010001: color_data = 12'b010000000000;
		14'b10100111010010: color_data = 12'b010000000000;
		14'b10100111010011: color_data = 12'b001000000000;
		14'b10100111010100: color_data = 12'b010000000000;
		14'b10100111010101: color_data = 12'b010000000000;
		14'b10100111010110: color_data = 12'b010000000000;
		14'b10100111010111: color_data = 12'b010000000000;
		14'b10100111011000: color_data = 12'b010000000000;
		14'b10100111011010: color_data = 12'b001000000000;
		14'b10100111011011: color_data = 12'b010000000000;
		14'b10100111011100: color_data = 12'b010000000000;
		14'b10100111011101: color_data = 12'b010000000000;
		14'b10100111011110: color_data = 12'b010000000000;
		14'b10100111011111: color_data = 12'b010000000000;
		14'b10100111100000: color_data = 12'b001000000000;
		14'b10100111111100: color_data = 12'b001000000000;
		14'b10100111111101: color_data = 12'b010000000000;
		14'b10100111111110: color_data = 12'b010000000000;
		14'b10100111111111: color_data = 12'b010000000000;
		14'b10101000000000: color_data = 12'b001000000000;
		14'b10101000000001: color_data = 12'b001000000000;
		14'b10101000011000: color_data = 12'b001000000000;
		14'b10101000011001: color_data = 12'b001000000000;
		14'b10101000100010: color_data = 12'b001000000000;
		14'b10101000100011: color_data = 12'b010000000000;
		14'b10101000100100: color_data = 12'b010000000000;
		14'b10101000100101: color_data = 12'b010000000000;
		14'b10101000100110: color_data = 12'b010000000000;
		14'b10101000100111: color_data = 12'b001000000000;
		14'b10101000101000: color_data = 12'b001000000000;
		14'b10101000101001: color_data = 12'b001000000000;
		14'b10101000101010: color_data = 12'b001000000000;
		14'b10101000101011: color_data = 12'b010000000000;
		14'b10101000101100: color_data = 12'b010000000000;
		14'b10101000101101: color_data = 12'b010000000000;
		14'b10101000101110: color_data = 12'b010000000000;
		14'b10101000101111: color_data = 12'b010000000000;
		14'b10101000110000: color_data = 12'b010000000000;
		14'b10101000110001: color_data = 12'b010000000000;
		14'b10101000110010: color_data = 12'b001000000000;
		14'b10101001000110: color_data = 12'b001000000000;
		14'b10101001000111: color_data = 12'b010000000000;
		14'b10101001001000: color_data = 12'b010000000000;
		14'b10101001001001: color_data = 12'b010000000000;
		14'b10101001001010: color_data = 12'b010000000000;
		14'b10101001001011: color_data = 12'b010000000000;
		14'b10101001001100: color_data = 12'b010000000000;
		14'b10101001001101: color_data = 12'b010000000000;
		14'b10101001001110: color_data = 12'b010000000000;
		14'b10101001001111: color_data = 12'b010000000000;
		14'b10101001010000: color_data = 12'b010000000000;
		14'b10101001010001: color_data = 12'b001000000000;
		14'b10101001010010: color_data = 12'b001000000000;
		14'b10101001010100: color_data = 12'b001000000000;
		14'b10101001010101: color_data = 12'b010000000000;
		14'b10101001010110: color_data = 12'b010000000000;
		14'b10101001010111: color_data = 12'b010000000000;
		14'b10101001011000: color_data = 12'b010000000000;
		14'b10101001011001: color_data = 12'b010000000000;
		14'b10101001011010: color_data = 12'b010000000000;
		14'b10101001011011: color_data = 12'b010000000000;
		14'b10101001011100: color_data = 12'b010000000000;
		14'b10101001011101: color_data = 12'b010000000000;
		14'b10101001011110: color_data = 12'b010000000000;
		14'b10101001011111: color_data = 12'b010000000000;
		14'b10101001100000: color_data = 12'b001000000000;
		14'b10101001111100: color_data = 12'b001000000000;
		14'b10101001111101: color_data = 12'b010000000000;
		14'b10101001111110: color_data = 12'b010000000000;
		14'b10101001111111: color_data = 12'b010000000000;
		14'b10101010000000: color_data = 12'b001000000000;
		14'b10101010000001: color_data = 12'b001000000000;
		14'b10101010001111: color_data = 12'b001000000000;
		14'b10101010010101: color_data = 12'b010000000000;
		14'b10101010011000: color_data = 12'b001000000000;
		14'b10101010011001: color_data = 12'b001000000000;
		14'b10101010100001: color_data = 12'b001000000000;
		14'b10101010100010: color_data = 12'b001000000000;
		14'b10101010100011: color_data = 12'b010000000000;
		14'b10101010100100: color_data = 12'b010000000000;
		14'b10101010100101: color_data = 12'b010000000000;
		14'b10101010100110: color_data = 12'b001000000000;
		14'b10101010100111: color_data = 12'b001000000000;
		14'b10101010101000: color_data = 12'b001000000000;
		14'b10101010101001: color_data = 12'b001000000000;
		14'b10101010101010: color_data = 12'b010000000000;
		14'b10101010101011: color_data = 12'b010000000000;
		14'b10101010101100: color_data = 12'b010000000000;
		14'b10101010101101: color_data = 12'b010000000000;
		14'b10101010101110: color_data = 12'b010000000000;
		14'b10101010101111: color_data = 12'b010000000000;
		14'b10101010110000: color_data = 12'b010000000000;
		14'b10101010110001: color_data = 12'b010000000000;
		14'b10101010110010: color_data = 12'b001000000000;
		14'b10101011000101: color_data = 12'b010000000000;
		14'b10101011000110: color_data = 12'b010000000000;
		14'b10101011000111: color_data = 12'b010000000000;
		14'b10101011001000: color_data = 12'b010000000000;
		14'b10101011001001: color_data = 12'b010000000000;
		14'b10101011001010: color_data = 12'b010000000000;
		14'b10101011001011: color_data = 12'b010000000000;
		14'b10101011001100: color_data = 12'b010000000000;
		14'b10101011001101: color_data = 12'b010000000000;
		14'b10101011001110: color_data = 12'b001000000000;
		14'b10101011001111: color_data = 12'b001000000000;
		14'b10101011010000: color_data = 12'b001000000000;
		14'b10101011010001: color_data = 12'b001000000000;
		14'b10101011010100: color_data = 12'b001000000000;
		14'b10101011010101: color_data = 12'b010000000000;
		14'b10101011010110: color_data = 12'b010000000000;
		14'b10101011010111: color_data = 12'b010000000000;
		14'b10101011011000: color_data = 12'b010000000000;
		14'b10101011011001: color_data = 12'b010000000000;
		14'b10101011011010: color_data = 12'b010000000000;
		14'b10101011011011: color_data = 12'b010000000000;
		14'b10101011011100: color_data = 12'b010000000000;
		14'b10101011011101: color_data = 12'b010000000000;
		14'b10101011011110: color_data = 12'b001000000000;
		14'b10101011011111: color_data = 12'b010000000000;
		14'b10101011100000: color_data = 12'b010000000000;
		14'b10101011111100: color_data = 12'b001000000000;
		14'b10101011111101: color_data = 12'b010000000000;
		14'b10101011111110: color_data = 12'b010000000000;
		14'b10101011111111: color_data = 12'b010000000000;
		14'b10101100000000: color_data = 12'b001000000000;
		14'b10101100000001: color_data = 12'b001000000000;
		14'b10101100010000: color_data = 12'b001000000000;
		14'b10101100010001: color_data = 12'b001000000000;
		14'b10101100010010: color_data = 12'b001000000000;
		14'b10101100010011: color_data = 12'b001000000000;
		14'b10101100010100: color_data = 12'b010000000000;
		14'b10101100010101: color_data = 12'b010000000000;
		14'b10101100010110: color_data = 12'b010000000000;
		14'b10101100010111: color_data = 12'b010000000000;
		14'b10101100011000: color_data = 12'b001000000000;
		14'b10101100011001: color_data = 12'b001000000000;
		14'b10101100100010: color_data = 12'b001000000000;
		14'b10101100100011: color_data = 12'b010000000000;
		14'b10101100100100: color_data = 12'b010000000000;
		14'b10101100100101: color_data = 12'b001000000000;
		14'b10101100100110: color_data = 12'b001000000000;
		14'b10101100100111: color_data = 12'b001000000000;
		14'b10101100101000: color_data = 12'b010000000000;
		14'b10101100101001: color_data = 12'b010000000000;
		14'b10101100101010: color_data = 12'b010000000000;
		14'b10101100101011: color_data = 12'b010000000000;
		14'b10101100101100: color_data = 12'b010000000000;
		14'b10101100101101: color_data = 12'b010000000000;
		14'b10101100101110: color_data = 12'b010000000000;
		14'b10101100101111: color_data = 12'b010000000000;
		14'b10101100110000: color_data = 12'b001000000000;
		14'b10101100110001: color_data = 12'b001000000000;
		14'b10101100110010: color_data = 12'b001000000000;
		14'b10101101000100: color_data = 12'b010000000000;
		14'b10101101000101: color_data = 12'b010000000000;
		14'b10101101000110: color_data = 12'b010000000000;
		14'b10101101000111: color_data = 12'b010000000000;
		14'b10101101001000: color_data = 12'b010000000000;
		14'b10101101001001: color_data = 12'b010000000000;
		14'b10101101001010: color_data = 12'b010000000000;
		14'b10101101001011: color_data = 12'b001000000000;
		14'b10101101001100: color_data = 12'b001000000000;
		14'b10101101001101: color_data = 12'b001000000000;
		14'b10101101001110: color_data = 12'b001000000000;
		14'b10101101010100: color_data = 12'b001000000000;
		14'b10101101010101: color_data = 12'b001000000000;
		14'b10101101010110: color_data = 12'b010000000000;
		14'b10101101010111: color_data = 12'b010000000000;
		14'b10101101011000: color_data = 12'b010000000000;
		14'b10101101011001: color_data = 12'b010000000000;
		14'b10101101011010: color_data = 12'b010000000000;
		14'b10101101011011: color_data = 12'b010000000000;
		14'b10101101011100: color_data = 12'b010000000000;
		14'b10101101011101: color_data = 12'b010000000000;
		14'b10101101011110: color_data = 12'b001000000000;
		14'b10101101011111: color_data = 12'b010000000000;
		14'b10101101100000: color_data = 12'b010000000000;
		14'b10101101100001: color_data = 12'b001000000000;
		14'b10101101111100: color_data = 12'b001000000000;
		14'b10101101111101: color_data = 12'b010000000000;
		14'b10101101111110: color_data = 12'b010000000000;
		14'b10101101111111: color_data = 12'b010000000000;
		14'b10101110000000: color_data = 12'b001000000000;
		14'b10101110000001: color_data = 12'b001000000000;
		14'b10101110010000: color_data = 12'b010000000000;
		14'b10101110010001: color_data = 12'b010000000000;
		14'b10101110010010: color_data = 12'b010000000000;
		14'b10101110010011: color_data = 12'b010000000000;
		14'b10101110010100: color_data = 12'b010000000000;
		14'b10101110010101: color_data = 12'b010000000000;
		14'b10101110010110: color_data = 12'b010000000000;
		14'b10101110010111: color_data = 12'b010000000000;
		14'b10101110011000: color_data = 12'b010000000000;
		14'b10101110011001: color_data = 12'b010000000000;
		14'b10101110011010: color_data = 12'b001000000000;
		14'b10101110100010: color_data = 12'b001000000000;
		14'b10101110100011: color_data = 12'b010000000000;
		14'b10101110100100: color_data = 12'b010000000000;
		14'b10101110100101: color_data = 12'b001000000000;
		14'b10101110100110: color_data = 12'b001000000000;
		14'b10101110100111: color_data = 12'b010000000000;
		14'b10101110101000: color_data = 12'b010000000000;
		14'b10101110101001: color_data = 12'b010000000000;
		14'b10101110101010: color_data = 12'b010000000000;
		14'b10101110101011: color_data = 12'b010000000000;
		14'b10101110101100: color_data = 12'b010000000000;
		14'b10101110101101: color_data = 12'b010000000000;
		14'b10101110101110: color_data = 12'b010000000000;
		14'b10101110101111: color_data = 12'b010000000000;
		14'b10101110110000: color_data = 12'b001000000000;
		14'b10101110110001: color_data = 12'b001000000000;
		14'b10101111000011: color_data = 12'b010000000000;
		14'b10101111000100: color_data = 12'b010000000000;
		14'b10101111000101: color_data = 12'b010000000000;
		14'b10101111000110: color_data = 12'b010000000000;
		14'b10101111000111: color_data = 12'b010000000000;
		14'b10101111001000: color_data = 12'b010000000000;
		14'b10101111001001: color_data = 12'b010000000000;
		14'b10101111001010: color_data = 12'b010000000000;
		14'b10101111010100: color_data = 12'b001000000000;
		14'b10101111010101: color_data = 12'b001000000000;
		14'b10101111010110: color_data = 12'b010000000000;
		14'b10101111010111: color_data = 12'b010000000000;
		14'b10101111011000: color_data = 12'b010000000000;
		14'b10101111011001: color_data = 12'b010000000000;
		14'b10101111011010: color_data = 12'b010000000000;
		14'b10101111011011: color_data = 12'b010000000000;
		14'b10101111011100: color_data = 12'b010000000000;
		14'b10101111011101: color_data = 12'b010000000000;
		14'b10101111011110: color_data = 12'b001000000000;
		14'b10101111011111: color_data = 12'b010000000000;
		14'b10101111100000: color_data = 12'b010000000000;
		14'b10101111100001: color_data = 12'b001000000000;
		14'b10101111111100: color_data = 12'b001000000000;
		14'b10101111111101: color_data = 12'b010000000000;
		14'b10101111111110: color_data = 12'b010000000000;
		14'b10101111111111: color_data = 12'b010000000000;
		14'b10110000000000: color_data = 12'b001000000000;
		14'b10110000000001: color_data = 12'b001000000000;
		14'b10110000001111: color_data = 12'b010000000000;
		14'b10110000010000: color_data = 12'b010000000000;
		14'b10110000010001: color_data = 12'b010000000000;
		14'b10110000010010: color_data = 12'b010000000000;
		14'b10110000010011: color_data = 12'b010000000000;
		14'b10110000010100: color_data = 12'b010000000000;
		14'b10110000010101: color_data = 12'b010000000000;
		14'b10110000010110: color_data = 12'b010000000000;
		14'b10110000010111: color_data = 12'b010000000000;
		14'b10110000011000: color_data = 12'b010000000000;
		14'b10110000011001: color_data = 12'b010000000000;
		14'b10110000011010: color_data = 12'b001000000000;
		14'b10110000100010: color_data = 12'b001000000000;
		14'b10110000100011: color_data = 12'b010000000000;
		14'b10110000100100: color_data = 12'b010000000000;
		14'b10110000100101: color_data = 12'b001000000000;
		14'b10110000100110: color_data = 12'b001000000000;
		14'b10110000100111: color_data = 12'b010000000000;
		14'b10110000101000: color_data = 12'b010000000000;
		14'b10110000101001: color_data = 12'b010000000000;
		14'b10110000101010: color_data = 12'b010000000000;
		14'b10110000101011: color_data = 12'b010000000000;
		14'b10110000101100: color_data = 12'b010000000000;
		14'b10110000101101: color_data = 12'b010000000000;
		14'b10110000101110: color_data = 12'b010000000000;
		14'b10110001000010: color_data = 12'b010000000000;
		14'b10110001000011: color_data = 12'b010000000000;
		14'b10110001000100: color_data = 12'b010000000000;
		14'b10110001000101: color_data = 12'b010000000000;
		14'b10110001000110: color_data = 12'b010000000000;
		14'b10110001000111: color_data = 12'b010000000000;
		14'b10110001001000: color_data = 12'b001000000000;
		14'b10110001010100: color_data = 12'b001000000000;
		14'b10110001010101: color_data = 12'b001000000000;
		14'b10110001010110: color_data = 12'b010000000000;
		14'b10110001010111: color_data = 12'b010000000000;
		14'b10110001011000: color_data = 12'b010000000000;
		14'b10110001011001: color_data = 12'b010000000000;
		14'b10110001011010: color_data = 12'b010000000000;
		14'b10110001011011: color_data = 12'b010000000000;
		14'b10110001011100: color_data = 12'b010000000000;
		14'b10110001011101: color_data = 12'b010000000000;
		14'b10110001100000: color_data = 12'b010000000000;
		14'b10110001100001: color_data = 12'b001000000000;
		14'b10110001111100: color_data = 12'b001000000000;
		14'b10110001111101: color_data = 12'b010000000000;
		14'b10110001111110: color_data = 12'b010000000000;
		14'b10110001111111: color_data = 12'b010000000000;
		14'b10110010000000: color_data = 12'b001000000000;
		14'b10110010000001: color_data = 12'b001000000000;
		14'b10110010001110: color_data = 12'b010000000000;
		14'b10110010001111: color_data = 12'b010000000000;
		14'b10110010010000: color_data = 12'b010000000000;
		14'b10110010010001: color_data = 12'b010000000000;
		14'b10110010010010: color_data = 12'b010000000000;
		14'b10110010010011: color_data = 12'b010000000000;
		14'b10110010010100: color_data = 12'b010000000000;
		14'b10110010010101: color_data = 12'b010000000000;
		14'b10110010010110: color_data = 12'b010000000000;
		14'b10110010010111: color_data = 12'b010000000000;
		14'b10110010011000: color_data = 12'b010000000000;
		14'b10110010011001: color_data = 12'b010000000000;
		14'b10110010011010: color_data = 12'b010000000000;
		14'b10110010011011: color_data = 12'b001000000000;
		14'b10110010100010: color_data = 12'b001000000000;
		14'b10110010100011: color_data = 12'b010000000000;
		14'b10110010100100: color_data = 12'b010000000000;
		14'b10110010100101: color_data = 12'b010000000000;
		14'b10110010100110: color_data = 12'b010000000000;
		14'b10110010100111: color_data = 12'b010000000000;
		14'b10110010101000: color_data = 12'b010000000000;
		14'b10110010101001: color_data = 12'b010000000000;
		14'b10110010101010: color_data = 12'b010000000000;
		14'b10110010101011: color_data = 12'b010000000000;
		14'b10110010101100: color_data = 12'b001000000000;
		14'b10110011000001: color_data = 12'b001000000000;
		14'b10110011000010: color_data = 12'b010000000000;
		14'b10110011000011: color_data = 12'b010000000000;
		14'b10110011000100: color_data = 12'b010000000000;
		14'b10110011000101: color_data = 12'b010000000000;
		14'b10110011010100: color_data = 12'b001000000000;
		14'b10110011010101: color_data = 12'b001000000000;
		14'b10110011010110: color_data = 12'b010000000000;
		14'b10110011010111: color_data = 12'b010000000000;
		14'b10110011011000: color_data = 12'b010000000000;
		14'b10110011011001: color_data = 12'b010000000000;
		14'b10110011011010: color_data = 12'b010000000000;
		14'b10110011011011: color_data = 12'b010000000000;
		14'b10110011011100: color_data = 12'b010000000000;
		14'b10110011011101: color_data = 12'b010000000000;
		14'b10110011100000: color_data = 12'b010000000000;
		14'b10110011100001: color_data = 12'b001000000000;
		14'b10110011111100: color_data = 12'b001000000000;
		14'b10110011111101: color_data = 12'b010000000000;
		14'b10110011111110: color_data = 12'b010000000000;
		14'b10110011111111: color_data = 12'b010000000000;
		14'b10110100000000: color_data = 12'b001000000000;
		14'b10110100000001: color_data = 12'b001000000000;
		14'b10110100001101: color_data = 12'b001000000000;
		14'b10110100001110: color_data = 12'b010000000000;
		14'b10110100001111: color_data = 12'b010000000000;
		14'b10110100010000: color_data = 12'b010000000000;
		14'b10110100010001: color_data = 12'b010000000000;
		14'b10110100010010: color_data = 12'b010000000000;
		14'b10110100010100: color_data = 12'b001000000000;
		14'b10110100010101: color_data = 12'b010000000000;
		14'b10110100010110: color_data = 12'b010000000000;
		14'b10110100010111: color_data = 12'b001000000000;
		14'b10110100011001: color_data = 12'b010000000000;
		14'b10110100011010: color_data = 12'b010000000000;
		14'b10110100011011: color_data = 12'b010000000000;
		14'b10110100100000: color_data = 12'b001000000000;
		14'b10110100100010: color_data = 12'b001000000000;
		14'b10110100100011: color_data = 12'b010000000000;
		14'b10110100100100: color_data = 12'b010000000000;
		14'b10110100100101: color_data = 12'b010000000000;
		14'b10110100100110: color_data = 12'b010000000000;
		14'b10110100100111: color_data = 12'b010000000000;
		14'b10110100101000: color_data = 12'b010000000000;
		14'b10110100101001: color_data = 12'b010000000000;
		14'b10110100101010: color_data = 12'b010000000000;
		14'b10110101000000: color_data = 12'b001000000000;
		14'b10110101000001: color_data = 12'b001000000000;
		14'b10110101000010: color_data = 12'b010000000000;
		14'b10110101000011: color_data = 12'b010000000000;
		14'b10110101000100: color_data = 12'b001000000000;
		14'b10110101010100: color_data = 12'b001000000000;
		14'b10110101010101: color_data = 12'b001000000000;
		14'b10110101010110: color_data = 12'b001000000000;
		14'b10110101010111: color_data = 12'b010000000000;
		14'b10110101011000: color_data = 12'b001000000000;
		14'b10110101011001: color_data = 12'b001000000000;
		14'b10110101011011: color_data = 12'b001000000000;
		14'b10110101011100: color_data = 12'b010000000000;
		14'b10110101011101: color_data = 12'b010000000000;
		14'b10110101100000: color_data = 12'b001000000000;
		14'b10110101100001: color_data = 12'b001000000000;
		14'b10110101111100: color_data = 12'b001000000000;
		14'b10110101111101: color_data = 12'b010000000000;
		14'b10110101111110: color_data = 12'b010000000000;
		14'b10110101111111: color_data = 12'b010000000000;
		14'b10110110000000: color_data = 12'b001000000000;
		14'b10110110000001: color_data = 12'b001000000000;
		14'b10110110001100: color_data = 12'b001000000000;
		14'b10110110001110: color_data = 12'b001000000000;
		14'b10110110001111: color_data = 12'b001000000000;
		14'b10110110010000: color_data = 12'b010000000000;
		14'b10110110010001: color_data = 12'b010000000000;
		14'b10110110010101: color_data = 12'b001000000000;
		14'b10110110010110: color_data = 12'b010000000000;
		14'b10110110010111: color_data = 12'b001000000000;
		14'b10110110011010: color_data = 12'b010000000000;
		14'b10110110011011: color_data = 12'b010000000000;
		14'b10110110011100: color_data = 12'b001000000000;
		14'b10110110100000: color_data = 12'b001000000000;
		14'b10110110100010: color_data = 12'b001000000000;
		14'b10110110100011: color_data = 12'b010000000000;
		14'b10110110100100: color_data = 12'b010000000000;
		14'b10110110100101: color_data = 12'b010000000000;
		14'b10110110100110: color_data = 12'b010000000000;
		14'b10110110100111: color_data = 12'b010000000000;
		14'b10110110101000: color_data = 12'b010000000000;
		14'b10110110101001: color_data = 12'b010000000000;
		14'b10110110101010: color_data = 12'b001000000000;
		14'b10110110111110: color_data = 12'b001000000000;
		14'b10110110111111: color_data = 12'b001000000000;
		14'b10110111000000: color_data = 12'b001000000000;
		14'b10110111000001: color_data = 12'b010000000000;
		14'b10110111000010: color_data = 12'b010000000000;
		14'b10110111000011: color_data = 12'b001000000000;
		14'b10110111010001: color_data = 12'b001000000000;
		14'b10110111010101: color_data = 12'b001000000000;
		14'b10110111010110: color_data = 12'b001000000000;
		14'b10110111010111: color_data = 12'b001000000000;
		14'b10110111011011: color_data = 12'b001000000000;
		14'b10110111011100: color_data = 12'b010000000000;
		14'b10110111011101: color_data = 12'b010000000000;
		14'b10110111100000: color_data = 12'b001000000000;
		14'b10110111100001: color_data = 12'b001000000000;
		14'b10110111111100: color_data = 12'b001000000000;
		14'b10110111111101: color_data = 12'b010000000000;
		14'b10110111111110: color_data = 12'b010000000000;
		14'b10110111111111: color_data = 12'b010000000000;
		14'b10111000000000: color_data = 12'b001000000000;
		14'b10111000000001: color_data = 12'b001000000000;
		14'b10111000001100: color_data = 12'b001000000000;
		14'b10111000001110: color_data = 12'b001000000000;
		14'b10111000001111: color_data = 12'b010000000000;
		14'b10111000010000: color_data = 12'b010000000000;
		14'b10111000010101: color_data = 12'b001000000000;
		14'b10111000010110: color_data = 12'b010000000000;
		14'b10111000010111: color_data = 12'b010000000000;
		14'b10111000011011: color_data = 12'b010000000000;
		14'b10111000011100: color_data = 12'b010000000000;
		14'b10111000011101: color_data = 12'b001000000000;
		14'b10111000100000: color_data = 12'b001000000000;
		14'b10111000100001: color_data = 12'b001000000000;
		14'b10111000100010: color_data = 12'b001000000000;
		14'b10111000100011: color_data = 12'b010000000000;
		14'b10111000100100: color_data = 12'b010000000000;
		14'b10111000100101: color_data = 12'b010000000000;
		14'b10111000100110: color_data = 12'b010000000000;
		14'b10111000100111: color_data = 12'b010000000000;
		14'b10111000101000: color_data = 12'b010000000000;
		14'b10111000101001: color_data = 12'b001000000000;
		14'b10111000101010: color_data = 12'b001000000000;
		14'b10111000111110: color_data = 12'b001000000000;
		14'b10111000111111: color_data = 12'b001000000000;
		14'b10111001000000: color_data = 12'b010000000000;
		14'b10111001000001: color_data = 12'b010000000000;
		14'b10111001000010: color_data = 12'b010000000000;
		14'b10111001000011: color_data = 12'b001000000000;
		14'b10111001010000: color_data = 12'b001000000000;
		14'b10111001010001: color_data = 12'b010000000000;
		14'b10111001010101: color_data = 12'b001000000000;
		14'b10111001010110: color_data = 12'b001000000000;
		14'b10111001010111: color_data = 12'b001000000000;
		14'b10111001011011: color_data = 12'b001000000000;
		14'b10111001011100: color_data = 12'b010000000000;
		14'b10111001011101: color_data = 12'b010000000000;
		14'b10111001100000: color_data = 12'b001000000000;
		14'b10111001100001: color_data = 12'b001000000000;
		14'b10111001111100: color_data = 12'b001000000000;
		14'b10111001111101: color_data = 12'b010000000000;
		14'b10111001111110: color_data = 12'b010000000000;
		14'b10111001111111: color_data = 12'b010000000000;
		14'b10111010000000: color_data = 12'b001000000000;
		14'b10111010000001: color_data = 12'b001000000000;
		14'b10111010001011: color_data = 12'b001000000000;
		14'b10111010001110: color_data = 12'b001000000000;
		14'b10111010001111: color_data = 12'b010000000000;
		14'b10111010010000: color_data = 12'b001000000000;
		14'b10111010010100: color_data = 12'b001000000000;
		14'b10111010010101: color_data = 12'b010000000000;
		14'b10111010010110: color_data = 12'b010000000000;
		14'b10111010010111: color_data = 12'b010000000000;
		14'b10111010011000: color_data = 12'b001000000000;
		14'b10111010011011: color_data = 12'b001000000000;
		14'b10111010011100: color_data = 12'b010000000000;
		14'b10111010011101: color_data = 12'b001000000000;
		14'b10111010100000: color_data = 12'b001000000000;
		14'b10111010100001: color_data = 12'b001000000000;
		14'b10111010100010: color_data = 12'b001000000000;
		14'b10111010100011: color_data = 12'b010000000000;
		14'b10111010100100: color_data = 12'b010000000000;
		14'b10111010100101: color_data = 12'b010000000000;
		14'b10111010100110: color_data = 12'b010000000000;
		14'b10111010100111: color_data = 12'b010000000000;
		14'b10111010101000: color_data = 12'b010000000000;
		14'b10111010101001: color_data = 12'b010000000000;
		14'b10111010101010: color_data = 12'b001000000000;
		14'b10111010111101: color_data = 12'b001000000000;
		14'b10111010111110: color_data = 12'b001000000000;
		14'b10111010111111: color_data = 12'b010000000000;
		14'b10111011000000: color_data = 12'b010000000000;
		14'b10111011000001: color_data = 12'b010000000000;
		14'b10111011000010: color_data = 12'b001000000000;
		14'b10111011011010: color_data = 12'b001000000000;
		14'b10111011011011: color_data = 12'b010000000000;
		14'b10111011011100: color_data = 12'b010000000000;
		14'b10111011011101: color_data = 12'b001000000000;
		14'b10111011100000: color_data = 12'b001000000000;
		14'b10111011100001: color_data = 12'b001000000000;
		14'b10111011111100: color_data = 12'b001000000000;
		14'b10111011111101: color_data = 12'b010000000000;
		14'b10111011111110: color_data = 12'b010000000000;
		14'b10111011111111: color_data = 12'b010000000000;
		14'b10111100000000: color_data = 12'b001000000000;
		14'b10111100000001: color_data = 12'b001000000000;
		14'b10111100001101: color_data = 12'b001000000000;
		14'b10111100001110: color_data = 12'b001000000000;
		14'b10111100001111: color_data = 12'b001000000000;
		14'b10111100010000: color_data = 12'b001000000000;
		14'b10111100010001: color_data = 12'b001000000000;
		14'b10111100010010: color_data = 12'b010000000000;
		14'b10111100010011: color_data = 12'b010000000000;
		14'b10111100010100: color_data = 12'b010000000000;
		14'b10111100010101: color_data = 12'b010000000000;
		14'b10111100010110: color_data = 12'b010000000000;
		14'b10111100010111: color_data = 12'b010000000000;
		14'b10111100011000: color_data = 12'b010000000000;
		14'b10111100011001: color_data = 12'b001000000000;
		14'b10111100011100: color_data = 12'b001000000000;
		14'b10111100011101: color_data = 12'b001000000000;
		14'b10111100100001: color_data = 12'b001000000000;
		14'b10111100100010: color_data = 12'b001000000000;
		14'b10111100100011: color_data = 12'b010000000000;
		14'b10111100100100: color_data = 12'b010000000000;
		14'b10111100100101: color_data = 12'b010000000000;
		14'b10111100100110: color_data = 12'b010000000000;
		14'b10111100100111: color_data = 12'b010000000000;
		14'b10111100101000: color_data = 12'b010000000000;
		14'b10111100101001: color_data = 12'b010000000000;
		14'b10111100101010: color_data = 12'b001000000000;
		14'b10111100111101: color_data = 12'b001000000000;
		14'b10111100111110: color_data = 12'b010000000000;
		14'b10111100111111: color_data = 12'b010000000000;
		14'b10111101000000: color_data = 12'b001000000000;
		14'b10111101000001: color_data = 12'b001000000000;
		14'b10111101010010: color_data = 12'b001000000000;
		14'b10111101010011: color_data = 12'b010000000000;
		14'b10111101011001: color_data = 12'b001000000000;
		14'b10111101011010: color_data = 12'b010000000000;
		14'b10111101011011: color_data = 12'b010000000000;
		14'b10111101011100: color_data = 12'b010000000000;
		14'b10111101011101: color_data = 12'b001000000000;
		14'b10111101100000: color_data = 12'b001000000000;
		14'b10111101111100: color_data = 12'b001000000000;
		14'b10111101111101: color_data = 12'b010000000000;
		14'b10111101111110: color_data = 12'b010000000000;
		14'b10111101111111: color_data = 12'b010000000000;
		14'b10111110000000: color_data = 12'b001000000000;
		14'b10111110000001: color_data = 12'b001000000000;
		14'b10111110001110: color_data = 12'b001000000000;
		14'b10111110001111: color_data = 12'b001000000000;
		14'b10111110010000: color_data = 12'b010000000000;
		14'b10111110010001: color_data = 12'b010000000000;
		14'b10111110010010: color_data = 12'b010000000000;
		14'b10111110010011: color_data = 12'b010000000000;
		14'b10111110010100: color_data = 12'b010000000000;
		14'b10111110010101: color_data = 12'b010000000000;
		14'b10111110010110: color_data = 12'b010000000000;
		14'b10111110010111: color_data = 12'b010000000000;
		14'b10111110011000: color_data = 12'b010000000000;
		14'b10111110011001: color_data = 12'b010000000000;
		14'b10111110011010: color_data = 12'b001000000000;
		14'b10111110011100: color_data = 12'b001000000000;
		14'b10111110011101: color_data = 12'b001000000000;
		14'b10111110100001: color_data = 12'b001000000000;
		14'b10111110100010: color_data = 12'b010000000000;
		14'b10111110100011: color_data = 12'b010000000000;
		14'b10111110100100: color_data = 12'b010000000000;
		14'b10111110100101: color_data = 12'b010000000000;
		14'b10111110100110: color_data = 12'b010000000000;
		14'b10111110100111: color_data = 12'b010000000000;
		14'b10111110101000: color_data = 12'b010000000000;
		14'b10111110101001: color_data = 12'b010000000000;
		14'b10111110101010: color_data = 12'b001000000000;
		14'b10111110111100: color_data = 12'b001000000000;
		14'b10111110111101: color_data = 12'b001000000000;
		14'b10111110111110: color_data = 12'b010000000000;
		14'b10111110111111: color_data = 12'b001000000000;
		14'b10111111000000: color_data = 12'b001000000000;
		14'b10111111000001: color_data = 12'b001000000000;
		14'b10111111010010: color_data = 12'b010000000000;
		14'b10111111010011: color_data = 12'b010000000000;
		14'b10111111011001: color_data = 12'b001000000000;
		14'b10111111011010: color_data = 12'b010000000000;
		14'b10111111011011: color_data = 12'b010000000000;
		14'b10111111011100: color_data = 12'b010000000000;
		14'b10111111011101: color_data = 12'b001000000000;
		14'b10111111111100: color_data = 12'b001000000000;
		14'b10111111111101: color_data = 12'b010000000000;
		14'b10111111111110: color_data = 12'b010000000000;
		14'b10111111111111: color_data = 12'b010000000000;
		14'b11000000000000: color_data = 12'b001000000000;
		14'b11000000000001: color_data = 12'b001000000000;
		14'b11000000001110: color_data = 12'b001000000000;
		14'b11000000001111: color_data = 12'b010000000000;
		14'b11000000010000: color_data = 12'b010000000000;
		14'b11000000010001: color_data = 12'b001000000000;
		14'b11000000010010: color_data = 12'b001000000000;
		14'b11000000010011: color_data = 12'b010000000000;
		14'b11000000010100: color_data = 12'b010000000000;
		14'b11000000010101: color_data = 12'b010000000000;
		14'b11000000010110: color_data = 12'b010000000000;
		14'b11000000010111: color_data = 12'b010000000000;
		14'b11000000011000: color_data = 12'b010000000000;
		14'b11000000011001: color_data = 12'b010000000000;
		14'b11000000011010: color_data = 12'b010000000000;
		14'b11000000011011: color_data = 12'b001000000000;
		14'b11000000011100: color_data = 12'b001000000000;
		14'b11000000011101: color_data = 12'b001000000000;
		14'b11000000100010: color_data = 12'b001000000000;
		14'b11000000100011: color_data = 12'b010000000000;
		14'b11000000100100: color_data = 12'b010000000000;
		14'b11000000100101: color_data = 12'b010000000000;
		14'b11000000100110: color_data = 12'b010000000000;
		14'b11000000100111: color_data = 12'b010000000000;
		14'b11000000101000: color_data = 12'b010000000000;
		14'b11000000101001: color_data = 12'b010000000000;
		14'b11000000101010: color_data = 12'b010000000000;
		14'b11000000101011: color_data = 12'b001000000000;
		14'b11000000111100: color_data = 12'b001000000000;
		14'b11000000111101: color_data = 12'b001000000000;
		14'b11000000111110: color_data = 12'b010000000000;
		14'b11000000111111: color_data = 12'b001000000000;
		14'b11000001000000: color_data = 12'b001000000000;
		14'b11000001000001: color_data = 12'b001000000000;
		14'b11000001011000: color_data = 12'b001000000000;
		14'b11000001011001: color_data = 12'b010000000000;
		14'b11000001011010: color_data = 12'b010000000000;
		14'b11000001011011: color_data = 12'b010000000000;
		14'b11000001011100: color_data = 12'b010000000000;
		14'b11000001111011: color_data = 12'b001000000000;
		14'b11000001111100: color_data = 12'b010000000000;
		14'b11000001111101: color_data = 12'b010000000000;
		14'b11000001111110: color_data = 12'b010000000000;
		14'b11000001111111: color_data = 12'b010000000000;
		14'b11000010000000: color_data = 12'b001000000000;
		14'b11000010000001: color_data = 12'b001000000000;
		14'b11000010001110: color_data = 12'b001000000000;
		14'b11000010001111: color_data = 12'b001000000000;
		14'b11000010010001: color_data = 12'b001000000000;
		14'b11000010010010: color_data = 12'b010000000000;
		14'b11000010010011: color_data = 12'b010000000000;
		14'b11000010010100: color_data = 12'b010000000000;
		14'b11000010010101: color_data = 12'b001000000000;
		14'b11000010010111: color_data = 12'b001000000000;
		14'b11000010011000: color_data = 12'b010000000000;
		14'b11000010011001: color_data = 12'b010000000000;
		14'b11000010011010: color_data = 12'b010000000000;
		14'b11000010011011: color_data = 12'b001000000000;
		14'b11000010011100: color_data = 12'b001000000000;
		14'b11000010011101: color_data = 12'b001000000000;
		14'b11000010100010: color_data = 12'b001000000000;
		14'b11000010100011: color_data = 12'b010000000000;
		14'b11000010100100: color_data = 12'b010000000000;
		14'b11000010100101: color_data = 12'b010000000000;
		14'b11000010100110: color_data = 12'b010000000000;
		14'b11000010100111: color_data = 12'b010000000000;
		14'b11000010101000: color_data = 12'b010000000000;
		14'b11000010101001: color_data = 12'b010000000000;
		14'b11000010101010: color_data = 12'b010000000000;
		14'b11000010101011: color_data = 12'b001000000000;
		14'b11000010111100: color_data = 12'b001000000000;
		14'b11000010111101: color_data = 12'b001000000000;
		14'b11000010111110: color_data = 12'b001000000000;
		14'b11000011000000: color_data = 12'b001000000000;
		14'b11000011000001: color_data = 12'b001000000000;
		14'b11000011010110: color_data = 12'b001000000000;
		14'b11000011010111: color_data = 12'b001000000000;
		14'b11000011011000: color_data = 12'b010000000000;
		14'b11000011011001: color_data = 12'b010000000000;
		14'b11000011011010: color_data = 12'b010000000000;
		14'b11000011011011: color_data = 12'b010000000000;
		14'b11000011011100: color_data = 12'b001000000000;
		14'b11000011111011: color_data = 12'b001000000000;
		14'b11000011111100: color_data = 12'b010000000000;
		14'b11000011111101: color_data = 12'b010000000000;
		14'b11000011111110: color_data = 12'b010000000000;
		14'b11000011111111: color_data = 12'b010000000000;
		14'b11000100000000: color_data = 12'b001000000000;
		14'b11000100000001: color_data = 12'b001000000000;
		14'b11000100010001: color_data = 12'b001000000000;
		14'b11000100010010: color_data = 12'b010000000000;
		14'b11000100010011: color_data = 12'b010000000000;
		14'b11000100010100: color_data = 12'b001000000000;
		14'b11000100010111: color_data = 12'b001000000000;
		14'b11000100011000: color_data = 12'b001000000000;
		14'b11000100011001: color_data = 12'b001000000000;
		14'b11000100011010: color_data = 12'b010000000000;
		14'b11000100011011: color_data = 12'b010000000000;
		14'b11000100011100: color_data = 12'b001000000000;
		14'b11000100011101: color_data = 12'b001000000000;
		14'b11000100100011: color_data = 12'b001000000000;
		14'b11000100100100: color_data = 12'b010000000000;
		14'b11000100100101: color_data = 12'b010000000000;
		14'b11000100100110: color_data = 12'b010000000000;
		14'b11000100100111: color_data = 12'b010000000000;
		14'b11000100101000: color_data = 12'b010000000000;
		14'b11000100101001: color_data = 12'b010000000000;
		14'b11000100101010: color_data = 12'b001000000000;
		14'b11000100101011: color_data = 12'b001000000000;
		14'b11000100111011: color_data = 12'b001000000000;
		14'b11000100111100: color_data = 12'b001000000000;
		14'b11000100111101: color_data = 12'b001000000000;
		14'b11000100111110: color_data = 12'b001000000000;
		14'b11000101000001: color_data = 12'b001000000000;
		14'b11000101010101: color_data = 12'b001000000000;
		14'b11000101010110: color_data = 12'b001000000000;
		14'b11000101010111: color_data = 12'b010000000000;
		14'b11000101011000: color_data = 12'b010000000000;
		14'b11000101011001: color_data = 12'b010000000000;
		14'b11000101011010: color_data = 12'b010000000000;
		14'b11000101011011: color_data = 12'b010000000000;
		14'b11000101011100: color_data = 12'b001000000000;
		14'b11000101111100: color_data = 12'b010000000000;
		14'b11000101111101: color_data = 12'b010000000000;
		14'b11000101111110: color_data = 12'b010000000000;
		14'b11000101111111: color_data = 12'b010000000000;
		14'b11000110000000: color_data = 12'b001000000000;
		14'b11000110010000: color_data = 12'b010000000000;
		14'b11000110010001: color_data = 12'b010000000000;
		14'b11000110010010: color_data = 12'b010000000000;
		14'b11000110010011: color_data = 12'b001000000000;
		14'b11000110010100: color_data = 12'b001000000000;
		14'b11000110010110: color_data = 12'b010000000000;
		14'b11000110010111: color_data = 12'b010000000000;
		14'b11000110011000: color_data = 12'b001000000000;
		14'b11000110011001: color_data = 12'b001000000000;
		14'b11000110011010: color_data = 12'b010000000000;
		14'b11000110011011: color_data = 12'b010000000000;
		14'b11000110011100: color_data = 12'b010000000000;
		14'b11000110011101: color_data = 12'b001000000000;
		14'b11000110100011: color_data = 12'b001000000000;
		14'b11000110100100: color_data = 12'b010000000000;
		14'b11000110100101: color_data = 12'b010000000000;
		14'b11000110100110: color_data = 12'b010000000000;
		14'b11000110100111: color_data = 12'b010000000000;
		14'b11000110101000: color_data = 12'b010000000000;
		14'b11000110101001: color_data = 12'b001000000000;
		14'b11000110101010: color_data = 12'b001000000000;
		14'b11000110111011: color_data = 12'b001000000000;
		14'b11000110111100: color_data = 12'b001000000000;
		14'b11000110111101: color_data = 12'b001000000000;
		14'b11000110111110: color_data = 12'b001000000000;
		14'b11000111000001: color_data = 12'b001000000000;
		14'b11000111000010: color_data = 12'b001000000000;
		14'b11000111010010: color_data = 12'b001000000000;
		14'b11000111010100: color_data = 12'b001000000000;
		14'b11000111010101: color_data = 12'b001000000000;
		14'b11000111010110: color_data = 12'b010000000000;
		14'b11000111010111: color_data = 12'b010000000000;
		14'b11000111011000: color_data = 12'b010000000000;
		14'b11000111011001: color_data = 12'b010000000000;
		14'b11000111011010: color_data = 12'b010000000000;
		14'b11000111011011: color_data = 12'b001000000000;
		14'b11000111111100: color_data = 12'b010000000000;
		14'b11000111111101: color_data = 12'b010000000000;
		14'b11000111111110: color_data = 12'b010000000000;
		14'b11000111111111: color_data = 12'b010000000000;
		14'b11001000000000: color_data = 12'b001000000000;
		14'b11001000001111: color_data = 12'b010000000000;
		14'b11001000010000: color_data = 12'b010000000000;
		14'b11001000010001: color_data = 12'b010000000000;
		14'b11001000010010: color_data = 12'b010000000000;
		14'b11001000010011: color_data = 12'b010000000000;
		14'b11001000010100: color_data = 12'b010000000000;
		14'b11001000010101: color_data = 12'b001000000000;
		14'b11001000010110: color_data = 12'b010000000000;
		14'b11001000010111: color_data = 12'b010000000000;
		14'b11001000011000: color_data = 12'b010000000000;
		14'b11001000011001: color_data = 12'b010000000000;
		14'b11001000011010: color_data = 12'b010000000000;
		14'b11001000011011: color_data = 12'b010000000000;
		14'b11001000011100: color_data = 12'b010000000000;
		14'b11001000011101: color_data = 12'b001000000000;
		14'b11001000100011: color_data = 12'b001000000000;
		14'b11001000100100: color_data = 12'b010000000000;
		14'b11001000100101: color_data = 12'b010000000000;
		14'b11001000100110: color_data = 12'b010000000000;
		14'b11001000100111: color_data = 12'b010000000000;
		14'b11001000101000: color_data = 12'b010000000000;
		14'b11001000101001: color_data = 12'b001000000000;
		14'b11001000111011: color_data = 12'b001000000000;
		14'b11001000111100: color_data = 12'b001000000000;
		14'b11001000111101: color_data = 12'b001000000000;
		14'b11001001000001: color_data = 12'b001000000000;
		14'b11001001000010: color_data = 12'b001000000000;
		14'b11001001010010: color_data = 12'b001000000000;
		14'b11001001010100: color_data = 12'b001000000000;
		14'b11001001010101: color_data = 12'b010000000000;
		14'b11001001010110: color_data = 12'b010000000000;
		14'b11001001010111: color_data = 12'b010000000000;
		14'b11001001011000: color_data = 12'b010000000000;
		14'b11001001011001: color_data = 12'b010000000000;
		14'b11001001011010: color_data = 12'b001000000000;
		14'b11001001111011: color_data = 12'b010000000000;
		14'b11001001111100: color_data = 12'b010000000000;
		14'b11001001111101: color_data = 12'b010000000000;
		14'b11001001111110: color_data = 12'b010000000000;
		14'b11001001111111: color_data = 12'b001000000000;
		14'b11001010000000: color_data = 12'b001000000000;
		14'b11001010001110: color_data = 12'b010000000000;
		14'b11001010001111: color_data = 12'b010000000000;
		14'b11001010010000: color_data = 12'b010000000000;
		14'b11001010010001: color_data = 12'b010000000000;
		14'b11001010010010: color_data = 12'b010000000000;
		14'b11001010010011: color_data = 12'b001000000000;
		14'b11001010010100: color_data = 12'b001000000000;
		14'b11001010010110: color_data = 12'b001000000000;
		14'b11001010010111: color_data = 12'b010000000000;
		14'b11001010011000: color_data = 12'b010000000000;
		14'b11001010011001: color_data = 12'b010000000000;
		14'b11001010011010: color_data = 12'b010000000000;
		14'b11001010011011: color_data = 12'b010000000000;
		14'b11001010011100: color_data = 12'b010000000000;
		14'b11001010011101: color_data = 12'b001000000000;
		14'b11001010100100: color_data = 12'b001000000000;
		14'b11001010100101: color_data = 12'b010000000000;
		14'b11001010100110: color_data = 12'b010000000000;
		14'b11001010100111: color_data = 12'b010000000000;
		14'b11001010101000: color_data = 12'b001000000000;
		14'b11001010111011: color_data = 12'b001000000000;
		14'b11001010111100: color_data = 12'b001000000000;
		14'b11001010111101: color_data = 12'b001000000000;
		14'b11001011000011: color_data = 12'b001000000000;
		14'b11001011010010: color_data = 12'b001000000000;
		14'b11001011010011: color_data = 12'b001000000000;
		14'b11001011010100: color_data = 12'b010000000000;
		14'b11001011010101: color_data = 12'b010000000000;
		14'b11001011010110: color_data = 12'b010000000000;
		14'b11001011010111: color_data = 12'b010000000000;
		14'b11001011011000: color_data = 12'b010000000000;
		14'b11001011011001: color_data = 12'b001000000000;
		14'b11001011111010: color_data = 12'b001000000000;
		14'b11001011111011: color_data = 12'b010000000000;
		14'b11001011111100: color_data = 12'b010000000000;
		14'b11001011111101: color_data = 12'b010000000000;
		14'b11001011111110: color_data = 12'b010000000000;
		14'b11001011111111: color_data = 12'b001000000000;
		14'b11001100001101: color_data = 12'b010000000000;
		14'b11001100001110: color_data = 12'b010000000000;
		14'b11001100001111: color_data = 12'b010000000000;
		14'b11001100010000: color_data = 12'b001000000000;
		14'b11001100010001: color_data = 12'b001000000000;
		14'b11001100010010: color_data = 12'b001000000000;
		14'b11001100010110: color_data = 12'b001000000000;
		14'b11001100010111: color_data = 12'b010000000000;
		14'b11001100011000: color_data = 12'b010000000000;
		14'b11001100011001: color_data = 12'b010000000000;
		14'b11001100011010: color_data = 12'b010000000000;
		14'b11001100011011: color_data = 12'b001000000000;
		14'b11001100011100: color_data = 12'b001000000000;
		14'b11001100011101: color_data = 12'b001000000000;
		14'b11001100100100: color_data = 12'b001000000000;
		14'b11001100100101: color_data = 12'b010000000000;
		14'b11001100100110: color_data = 12'b010000000000;
		14'b11001100100111: color_data = 12'b010000000000;
		14'b11001100101000: color_data = 12'b001000000000;
		14'b11001100111011: color_data = 12'b001000000000;
		14'b11001100111100: color_data = 12'b001000000000;
		14'b11001101010010: color_data = 12'b010000000000;
		14'b11001101010011: color_data = 12'b010000000000;
		14'b11001101010100: color_data = 12'b010000000000;
		14'b11001101010101: color_data = 12'b010000000000;
		14'b11001101010110: color_data = 12'b010000000000;
		14'b11001101010111: color_data = 12'b010000000000;
		14'b11001101011000: color_data = 12'b001000000000;
		14'b11001101111010: color_data = 12'b001000000000;
		14'b11001101111011: color_data = 12'b010000000000;
		14'b11001101111100: color_data = 12'b010000000000;
		14'b11001101111101: color_data = 12'b010000000000;
		14'b11001101111110: color_data = 12'b001000000000;
		14'b11001101111111: color_data = 12'b001000000000;
		14'b11001110001100: color_data = 12'b010000000000;
		14'b11001110001101: color_data = 12'b010000000000;
		14'b11001110001110: color_data = 12'b010000000000;
		14'b11001110001111: color_data = 12'b010000000000;
		14'b11001110010110: color_data = 12'b001000000000;
		14'b11001110010111: color_data = 12'b010000000000;
		14'b11001110011000: color_data = 12'b010000000000;
		14'b11001110011001: color_data = 12'b010000000000;
		14'b11001110011010: color_data = 12'b010000000000;
		14'b11001110011011: color_data = 12'b001000000000;
		14'b11001110011100: color_data = 12'b001000000000;
		14'b11001110100100: color_data = 12'b001000000000;
		14'b11001110100101: color_data = 12'b010000000000;
		14'b11001110100110: color_data = 12'b010000000000;
		14'b11001110100111: color_data = 12'b010000000000;
		14'b11001110101000: color_data = 12'b001000000000;
		14'b11001110111011: color_data = 12'b001000000000;
		14'b11001110111100: color_data = 12'b001000000000;
		14'b11001111010001: color_data = 12'b010000000000;
		14'b11001111010010: color_data = 12'b010000000000;
		14'b11001111010011: color_data = 12'b010000000000;
		14'b11001111010100: color_data = 12'b010000000000;
		14'b11001111010101: color_data = 12'b010000000000;
		14'b11001111010110: color_data = 12'b010000000000;
		14'b11001111010111: color_data = 12'b010000000000;
		14'b11001111111010: color_data = 12'b010000000000;
		14'b11001111111011: color_data = 12'b010000000000;
		14'b11001111111100: color_data = 12'b010000000000;
		14'b11001111111101: color_data = 12'b010000000000;
		14'b11001111111110: color_data = 12'b001000000000;
		14'b11001111111111: color_data = 12'b001000000000;
		14'b11010000001011: color_data = 12'b010000000000;
		14'b11010000001100: color_data = 12'b010000000000;
		14'b11010000001101: color_data = 12'b010000000000;
		14'b11010000010110: color_data = 12'b001000000000;
		14'b11010000010111: color_data = 12'b010000000000;
		14'b11010000011000: color_data = 12'b010000000000;
		14'b11010000011001: color_data = 12'b010000000000;
		14'b11010000011010: color_data = 12'b010000000000;
		14'b11010000011011: color_data = 12'b001000000000;
		14'b11010000011100: color_data = 12'b001000000000;
		14'b11010000100101: color_data = 12'b010000000000;
		14'b11010000100110: color_data = 12'b010000000000;
		14'b11010000100111: color_data = 12'b010000000000;
		14'b11010000101000: color_data = 12'b001000000000;
		14'b11010000111011: color_data = 12'b001000000000;
		14'b11010000111100: color_data = 12'b001000000000;
		14'b11010001010000: color_data = 12'b001000000000;
		14'b11010001010001: color_data = 12'b010000000000;
		14'b11010001010010: color_data = 12'b010000000000;
		14'b11010001010011: color_data = 12'b010000000000;
		14'b11010001010100: color_data = 12'b010000000000;
		14'b11010001010101: color_data = 12'b010000000000;
		14'b11010001010110: color_data = 12'b010000000000;
		14'b11010001111001: color_data = 12'b010000000000;
		14'b11010001111010: color_data = 12'b010000000000;
		14'b11010001111011: color_data = 12'b010000000000;
		14'b11010001111100: color_data = 12'b010000000000;
		14'b11010001111101: color_data = 12'b010000000000;
		14'b11010001111110: color_data = 12'b001000000000;
		14'b11010010001010: color_data = 12'b001000000000;
		14'b11010010001011: color_data = 12'b010000000000;
		14'b11010010001100: color_data = 12'b001000000000;
		14'b11010010010110: color_data = 12'b001000000000;
		14'b11010010011001: color_data = 12'b001000000000;
		14'b11010010011010: color_data = 12'b001000000000;
		14'b11010010100101: color_data = 12'b010000000000;
		14'b11010010100110: color_data = 12'b010000000000;
		14'b11010010100111: color_data = 12'b010000000000;
		14'b11010010101000: color_data = 12'b001000000000;
		14'b11010010111011: color_data = 12'b001000000000;
		14'b11010010111100: color_data = 12'b001000000000;
		14'b11010011001110: color_data = 12'b001000000000;
		14'b11010011001111: color_data = 12'b001000000000;
		14'b11010011010000: color_data = 12'b001000000000;
		14'b11010011010001: color_data = 12'b010000000000;
		14'b11010011010010: color_data = 12'b010000000000;
		14'b11010011010011: color_data = 12'b010000000000;
		14'b11010011010100: color_data = 12'b010000000000;
		14'b11010011010101: color_data = 12'b001000000000;
		14'b11010011111000: color_data = 12'b001000000000;
		14'b11010011111001: color_data = 12'b010000000000;
		14'b11010011111010: color_data = 12'b010000000000;
		14'b11010011111011: color_data = 12'b010000000000;
		14'b11010011111100: color_data = 12'b010000000000;
		14'b11010011111101: color_data = 12'b001000000000;
		14'b11010100001001: color_data = 12'b001000000000;
		14'b11010100001010: color_data = 12'b010000000000;
		14'b11010100001011: color_data = 12'b010000000000;
		14'b11010100011001: color_data = 12'b001000000000;
		14'b11010100011010: color_data = 12'b001000000000;
		14'b11010100100101: color_data = 12'b001000000000;
		14'b11010100100110: color_data = 12'b010000000000;
		14'b11010100100111: color_data = 12'b010000000000;
		14'b11010100101000: color_data = 12'b001000000000;
		14'b11010100101001: color_data = 12'b001000000000;
		14'b11010100111011: color_data = 12'b001000000000;
		14'b11010100111100: color_data = 12'b001000000000;
		14'b11010101001101: color_data = 12'b001000000000;
		14'b11010101001110: color_data = 12'b001000000000;
		14'b11010101001111: color_data = 12'b001000000000;
		14'b11010101010000: color_data = 12'b010000000000;
		14'b11010101010001: color_data = 12'b010000000000;
		14'b11010101010010: color_data = 12'b010000000000;
		14'b11010101010011: color_data = 12'b001000000000;
		14'b11010101010100: color_data = 12'b001000000000;
		14'b11010101110111: color_data = 12'b001000000000;
		14'b11010101111000: color_data = 12'b001000000000;
		14'b11010101111001: color_data = 12'b010000000000;
		14'b11010101111010: color_data = 12'b010000000000;
		14'b11010101111011: color_data = 12'b001000000000;
		14'b11010101111100: color_data = 12'b001000000000;
		14'b11010110001000: color_data = 12'b001000000000;
		14'b11010110001001: color_data = 12'b010000000000;
		14'b11010110001010: color_data = 12'b010000000000;
		14'b11010110010100: color_data = 12'b001000000000;
		14'b11010110011000: color_data = 12'b001000000000;
		14'b11010110011001: color_data = 12'b010000000000;
		14'b11010110011010: color_data = 12'b001000000000;
		14'b11010110100101: color_data = 12'b001000000000;
		14'b11010110100110: color_data = 12'b010000000000;
		14'b11010110100111: color_data = 12'b010000000000;
		14'b11010110101000: color_data = 12'b001000000000;
		14'b11010110101001: color_data = 12'b001000000000;
		14'b11010110111100: color_data = 12'b001000000000;
		14'b11010111001101: color_data = 12'b001000000000;
		14'b11010111001110: color_data = 12'b001000000000;
		14'b11010111001111: color_data = 12'b001000000000;
		14'b11010111010000: color_data = 12'b001000000000;
		14'b11010111010001: color_data = 12'b001000000000;
		14'b11010111010010: color_data = 12'b001000000000;
		14'b11010111110110: color_data = 12'b001000000000;
		14'b11010111110111: color_data = 12'b001000000000;
		14'b11010111111000: color_data = 12'b010000000000;
		14'b11010111111001: color_data = 12'b010000000000;
		14'b11010111111010: color_data = 12'b001000000000;
		14'b11010111111011: color_data = 12'b001000000000;
		14'b11010111111100: color_data = 12'b001000000000;
		14'b11011000001000: color_data = 12'b001000000000;
		14'b11011000001001: color_data = 12'b010000000000;
		14'b11011000010100: color_data = 12'b001000000000;
		14'b11011000011000: color_data = 12'b010000000000;
		14'b11011000011001: color_data = 12'b010000000000;
		14'b11011000011010: color_data = 12'b001000000000;
		14'b11011000100101: color_data = 12'b001000000000;
		14'b11011000100110: color_data = 12'b010000000000;
		14'b11011000100111: color_data = 12'b010000000000;
		14'b11011000101000: color_data = 12'b001000000000;
		14'b11011000101001: color_data = 12'b001000000000;
		14'b11011000111100: color_data = 12'b001000000000;
		14'b11011001001100: color_data = 12'b001000000000;
		14'b11011001001101: color_data = 12'b001000000000;
		14'b11011001001110: color_data = 12'b001000000000;
		14'b11011001001111: color_data = 12'b001000000000;
		14'b11011001010000: color_data = 12'b001000000000;
		14'b11011001010001: color_data = 12'b001000000000;
		14'b11011001010010: color_data = 12'b001000000000;
		14'b11011001110110: color_data = 12'b001000000000;
		14'b11011001110111: color_data = 12'b001000000000;
		14'b11011001111000: color_data = 12'b010000000000;
		14'b11011001111001: color_data = 12'b001000000000;
		14'b11011001111010: color_data = 12'b001000000000;
		14'b11011001111011: color_data = 12'b001000000000;
		14'b11011001111100: color_data = 12'b010000000000;
		14'b11011001111101: color_data = 12'b001000000000;
		14'b11011010000111: color_data = 12'b001000000000;
		14'b11011010001000: color_data = 12'b001000000000;
		14'b11011010001001: color_data = 12'b001000000000;
		14'b11011010010111: color_data = 12'b001000000000;
		14'b11011010011000: color_data = 12'b010000000000;
		14'b11011010011001: color_data = 12'b010000000000;
		14'b11011010100101: color_data = 12'b001000000000;
		14'b11011010100110: color_data = 12'b010000000000;
		14'b11011010100111: color_data = 12'b010000000000;
		14'b11011010101000: color_data = 12'b001000000000;
		14'b11011010101001: color_data = 12'b001000000000;
		14'b11011010111100: color_data = 12'b001000000000;
		14'b11011011001011: color_data = 12'b001000000000;
		14'b11011011001100: color_data = 12'b001000000000;
		14'b11011011001101: color_data = 12'b001000000000;
		14'b11011011001110: color_data = 12'b001000000000;
		14'b11011011001111: color_data = 12'b001000000000;
		14'b11011011010000: color_data = 12'b001000000000;
		14'b11011011010001: color_data = 12'b001000000000;
		14'b11011011110111: color_data = 12'b001000000000;
		14'b11011011111000: color_data = 12'b010000000000;
		14'b11011011111001: color_data = 12'b001000000000;
		14'b11011011111010: color_data = 12'b001000000000;
		14'b11011011111011: color_data = 12'b010000000000;
		14'b11011011111100: color_data = 12'b010000000000;
		14'b11011100000111: color_data = 12'b001000000000;
		14'b11011100001000: color_data = 12'b001000000000;
		14'b11011100001001: color_data = 12'b001000000000;
		14'b11011100010110: color_data = 12'b001000000000;
		14'b11011100010111: color_data = 12'b010000000000;
		14'b11011100011000: color_data = 12'b010000000000;
		14'b11011100011001: color_data = 12'b001000000000;
		14'b11011100100110: color_data = 12'b010000000000;
		14'b11011100100111: color_data = 12'b010000000000;
		14'b11011100101000: color_data = 12'b001000000000;
		14'b11011100101001: color_data = 12'b001000000000;
		14'b11011101001011: color_data = 12'b001000000000;
		14'b11011101001100: color_data = 12'b001000000000;
		14'b11011101001101: color_data = 12'b001000000000;
		14'b11011101001110: color_data = 12'b001000000000;
		14'b11011101001111: color_data = 12'b001000000000;
		14'b11011101110111: color_data = 12'b001000000000;
		14'b11011101111000: color_data = 12'b001000000000;
		14'b11011101111001: color_data = 12'b001000000000;
		14'b11011101111010: color_data = 12'b001000000000;
		14'b11011101111011: color_data = 12'b001000000000;
		14'b11011101111100: color_data = 12'b001000000000;
		14'b11011110000111: color_data = 12'b001000000000;
		14'b11011110001000: color_data = 12'b001000000000;
		14'b11011110001010: color_data = 12'b001000000000;
		14'b11011110010101: color_data = 12'b001000000000;
		14'b11011110010110: color_data = 12'b010000000000;
		14'b11011110010111: color_data = 12'b010000000000;
		14'b11011110011000: color_data = 12'b010000000000;
		14'b11011110100110: color_data = 12'b010000000000;
		14'b11011110100111: color_data = 12'b010000000000;
		14'b11011110101000: color_data = 12'b010000000000;
		14'b11011110101001: color_data = 12'b001000000000;
		14'b11011110101010: color_data = 12'b001000000000;
		14'b11011111001011: color_data = 12'b001000000000;
		14'b11011111001100: color_data = 12'b001000000000;
		14'b11011111001101: color_data = 12'b001000000000;
		14'b11011111110101: color_data = 12'b001000000000;
		14'b11011111110110: color_data = 12'b001000000000;
		14'b11011111110111: color_data = 12'b001000000000;
		14'b11011111111000: color_data = 12'b001000000000;
		14'b11011111111001: color_data = 12'b001000000000;
		14'b11011111111010: color_data = 12'b001000000000;
		14'b11100000000111: color_data = 12'b001000000000;
		14'b11100000001010: color_data = 12'b001000000000;
		14'b11100000001011: color_data = 12'b001000000000;
		14'b11100000010100: color_data = 12'b001000000000;
		14'b11100000010101: color_data = 12'b010000000000;
		14'b11100000010110: color_data = 12'b010000000000;
		14'b11100000010111: color_data = 12'b010000000000;
		14'b11100000100101: color_data = 12'b001000000000;
		14'b11100000100110: color_data = 12'b010000000000;
		14'b11100000100111: color_data = 12'b010000000000;
		14'b11100000101000: color_data = 12'b010000000000;
		14'b11100000101001: color_data = 12'b001000000000;
		14'b11100000101010: color_data = 12'b001000000000;
		14'b11100000101011: color_data = 12'b001000000000;
		14'b11100001001011: color_data = 12'b001000000000;
		14'b11100001110100: color_data = 12'b001000000000;
		14'b11100001110101: color_data = 12'b001000000000;
		14'b11100001110110: color_data = 12'b001000000000;
		14'b11100001110111: color_data = 12'b001000000000;
		14'b11100001111000: color_data = 12'b001000000000;
		14'b11100010000111: color_data = 12'b001000000000;
		14'b11100010010011: color_data = 12'b001000000000;
		14'b11100010010100: color_data = 12'b010000000000;
		14'b11100010010101: color_data = 12'b010000000000;
		14'b11100010010110: color_data = 12'b010000000000;
		14'b11100010010111: color_data = 12'b001000000000;
		14'b11100010100101: color_data = 12'b001000000000;
		14'b11100010100110: color_data = 12'b010000000000;
		14'b11100010100111: color_data = 12'b010000000000;
		14'b11100010101000: color_data = 12'b010000000000;
		14'b11100010101001: color_data = 12'b010000000000;
		14'b11100010101010: color_data = 12'b001000000000;
		14'b11100010101011: color_data = 12'b001000000000;
		14'b11100010101100: color_data = 12'b001000000000;
		14'b11100011001010: color_data = 12'b001000000000;
		14'b11100011001011: color_data = 12'b001000000000;
		14'b11100011110011: color_data = 12'b001000000000;
		14'b11100011110100: color_data = 12'b010000000000;
		14'b11100011110101: color_data = 12'b001000000000;
		14'b11100011110110: color_data = 12'b001000000000;
		14'b11100100010010: color_data = 12'b001000000000;
		14'b11100100010011: color_data = 12'b010000000000;
		14'b11100100010100: color_data = 12'b010000000000;
		14'b11100100010101: color_data = 12'b010000000000;
		14'b11100100100101: color_data = 12'b001000000000;
		14'b11100100100110: color_data = 12'b010000000000;
		14'b11100100100111: color_data = 12'b010000000000;
		14'b11100100101000: color_data = 12'b010000000000;
		14'b11100100101001: color_data = 12'b010000000000;
		14'b11100100101010: color_data = 12'b010000000000;
		14'b11100100101011: color_data = 12'b001000000000;
		14'b11100100101100: color_data = 12'b001000000000;
		14'b11100100101101: color_data = 12'b001000000000;
		14'b11100100101110: color_data = 12'b001000000000;
		14'b11100101001011: color_data = 12'b001000000000;
		14'b11100101110010: color_data = 12'b001000000000;
		14'b11100101110011: color_data = 12'b010000000000;
		14'b11100101110100: color_data = 12'b010000000000;
		14'b11100101110101: color_data = 12'b001000000000;
		14'b11100110010001: color_data = 12'b001000000000;
		14'b11100110010010: color_data = 12'b010000000000;
		14'b11100110010011: color_data = 12'b010000000000;
		14'b11100110010100: color_data = 12'b001000000000;
		14'b11100110100101: color_data = 12'b010000000000;
		14'b11100110100110: color_data = 12'b010000000000;
		14'b11100110100111: color_data = 12'b001000000000;
		14'b11100110101000: color_data = 12'b010000000000;
		14'b11100110101001: color_data = 12'b010000000000;
		14'b11100110101010: color_data = 12'b010000000000;
		14'b11100110101011: color_data = 12'b001000000000;
		14'b11100110101100: color_data = 12'b001000000000;
		14'b11100110101101: color_data = 12'b001000000000;
		14'b11100110101110: color_data = 12'b001000000000;
		14'b11100110101111: color_data = 12'b001000000000;
		14'b11100111001011: color_data = 12'b001000000000;
		14'b11100111110001: color_data = 12'b001000000000;
		14'b11100111110010: color_data = 12'b010000000000;
		14'b11100111110011: color_data = 12'b010000000000;
		14'b11100111110100: color_data = 12'b001000000000;
		14'b11101000010001: color_data = 12'b001000000000;
		14'b11101000010010: color_data = 12'b001000000000;
		14'b11101000010011: color_data = 12'b001000000000;
		14'b11101000100100: color_data = 12'b010000000000;
		14'b11101000100101: color_data = 12'b010000000000;
		14'b11101000100110: color_data = 12'b010000000000;
		14'b11101000100111: color_data = 12'b001000000000;
		14'b11101000101000: color_data = 12'b001000000000;
		14'b11101000101001: color_data = 12'b010000000000;
		14'b11101000101010: color_data = 12'b010000000000;
		14'b11101000101011: color_data = 12'b010000000000;
		14'b11101000101100: color_data = 12'b010000000000;
		14'b11101000101101: color_data = 12'b001000000000;
		14'b11101000101110: color_data = 12'b001000000000;
		14'b11101000101111: color_data = 12'b001000000000;
		14'b11101001001011: color_data = 12'b001000000000;
		14'b11101001110001: color_data = 12'b001000000000;
		14'b11101001110010: color_data = 12'b010000000000;
		14'b11101001110011: color_data = 12'b010000000000;
		14'b11101010010000: color_data = 12'b001000000000;
		14'b11101010010001: color_data = 12'b001000000000;
		14'b11101010010010: color_data = 12'b001000000000;
		14'b11101010100011: color_data = 12'b010000000000;
		14'b11101010100100: color_data = 12'b010000000000;
		14'b11101010100101: color_data = 12'b010000000000;
		14'b11101010100110: color_data = 12'b010000000000;
		14'b11101010100111: color_data = 12'b001000000000;
		14'b11101010101000: color_data = 12'b001000000000;
		14'b11101010101001: color_data = 12'b010000000000;
		14'b11101010101010: color_data = 12'b010000000000;
		14'b11101010101011: color_data = 12'b010000000000;
		14'b11101010101100: color_data = 12'b010000000000;
		14'b11101010101101: color_data = 12'b010000000000;
		14'b11101010101110: color_data = 12'b001000000000;
		14'b11101010101111: color_data = 12'b001000000000;
		14'b11101010110000: color_data = 12'b001000000000;
		14'b11101011001100: color_data = 12'b001000000000;
		14'b11101011110000: color_data = 12'b001000000000;
		14'b11101011110001: color_data = 12'b010000000000;
		14'b11101011110010: color_data = 12'b010000000000;
		14'b11101011110011: color_data = 12'b001000000000;
		14'b11101100001111: color_data = 12'b001000000000;
		14'b11101100010000: color_data = 12'b001000000000;
		14'b11101100100001: color_data = 12'b010000000000;
		14'b11101100100010: color_data = 12'b010000000000;
		14'b11101100100011: color_data = 12'b010000000000;
		14'b11101100100100: color_data = 12'b010000000000;
		14'b11101100100101: color_data = 12'b010000000000;
		14'b11101100100110: color_data = 12'b010000000000;
		14'b11101100100111: color_data = 12'b001000000000;
		14'b11101100101000: color_data = 12'b001000000000;
		14'b11101100101001: color_data = 12'b010000000000;
		14'b11101100101010: color_data = 12'b010000000000;
		14'b11101100101011: color_data = 12'b010000000000;
		14'b11101100101100: color_data = 12'b010000000000;
		14'b11101100101101: color_data = 12'b010000000000;
		14'b11101100101110: color_data = 12'b010000000000;
		14'b11101100101111: color_data = 12'b001000000000;
		14'b11101100110000: color_data = 12'b001000000000;
		14'b11101101101110: color_data = 12'b001000000000;
		14'b11101101101111: color_data = 12'b001000000000;
		14'b11101101110000: color_data = 12'b010000000000;
		14'b11101101110001: color_data = 12'b010000000000;
		14'b11101101110010: color_data = 12'b010000000000;
		14'b11101101110011: color_data = 12'b001000000000;
		14'b11101110001111: color_data = 12'b001000000000;
		14'b11101110011110: color_data = 12'b010000000000;
		14'b11101110011111: color_data = 12'b010000000000;
		14'b11101110100000: color_data = 12'b010000000000;
		14'b11101110100001: color_data = 12'b010000000000;
		14'b11101110100010: color_data = 12'b010000000000;
		14'b11101110100011: color_data = 12'b010000000000;
		14'b11101110100100: color_data = 12'b010000000000;
		14'b11101110100101: color_data = 12'b010000000000;
		14'b11101110100110: color_data = 12'b001000000000;
		14'b11101110100111: color_data = 12'b001000000000;
		14'b11101110101000: color_data = 12'b010000000000;
		14'b11101110101001: color_data = 12'b010000000000;
		14'b11101110101010: color_data = 12'b010000000000;
		14'b11101110101011: color_data = 12'b010000000000;
		14'b11101110101100: color_data = 12'b010000000000;
		14'b11101110101101: color_data = 12'b010000000000;
		14'b11101110101110: color_data = 12'b010000000000;
		14'b11101110101111: color_data = 12'b001000000000;
		14'b11101110110000: color_data = 12'b001000000000;
		14'b11101111101100: color_data = 12'b001000000000;
		14'b11101111101101: color_data = 12'b001000000000;
		14'b11101111101110: color_data = 12'b001000000000;
		14'b11101111101111: color_data = 12'b010000000000;
		14'b11101111110000: color_data = 12'b010000000000;
		14'b11101111110001: color_data = 12'b010000000000;
		14'b11101111110010: color_data = 12'b001000000000;
		14'b11101111110011: color_data = 12'b001000000000;
		14'b11110000011010: color_data = 12'b001000000000;
		14'b11110000011011: color_data = 12'b010000000000;
		14'b11110000011100: color_data = 12'b010000000000;
		14'b11110000011101: color_data = 12'b010000000000;
		14'b11110000011110: color_data = 12'b010000000000;
		14'b11110000011111: color_data = 12'b010000000000;
		14'b11110000100000: color_data = 12'b010000000000;
		14'b11110000100001: color_data = 12'b010000000000;
		14'b11110000100010: color_data = 12'b010000000000;
		14'b11110000100011: color_data = 12'b010000000000;
		14'b11110000100100: color_data = 12'b010000000000;
		14'b11110000100101: color_data = 12'b001000000000;
		14'b11110000100110: color_data = 12'b001000000000;
		14'b11110000100111: color_data = 12'b001000000000;
		14'b11110000101000: color_data = 12'b010000000000;
		14'b11110000101001: color_data = 12'b010000000000;
		14'b11110000101010: color_data = 12'b010000000000;
		14'b11110000101011: color_data = 12'b010000000000;
		14'b11110000101100: color_data = 12'b010000000000;
		14'b11110000101101: color_data = 12'b010000000000;
		14'b11110000101110: color_data = 12'b010000000000;
		14'b11110000101111: color_data = 12'b001000000000;
		14'b11110000110000: color_data = 12'b001000000000;
		14'b11110001101010: color_data = 12'b001000000000;
		14'b11110001101011: color_data = 12'b001000000000;
		14'b11110001101100: color_data = 12'b001000000000;
		14'b11110001101101: color_data = 12'b001000000000;
		14'b11110001101110: color_data = 12'b001000000000;
		14'b11110001101111: color_data = 12'b010000000000;
		14'b11110001110000: color_data = 12'b010000000000;
		14'b11110001110001: color_data = 12'b010000000000;
		14'b11110001110010: color_data = 12'b001000000000;
		14'b11110001110011: color_data = 12'b001000000000;
		14'b11110010010111: color_data = 12'b001000000000;
		14'b11110010011000: color_data = 12'b010000000000;
		14'b11110010011001: color_data = 12'b010000000000;
		14'b11110010011010: color_data = 12'b010000000000;
		14'b11110010011011: color_data = 12'b010000000000;
		14'b11110010011100: color_data = 12'b010000000000;
		14'b11110010011101: color_data = 12'b010000000000;
		14'b11110010011110: color_data = 12'b010000000000;
		14'b11110010011111: color_data = 12'b010000000000;
		14'b11110010100000: color_data = 12'b010000000000;
		14'b11110010100001: color_data = 12'b010000000000;
		14'b11110010100010: color_data = 12'b010000000000;
		14'b11110010100011: color_data = 12'b010000000000;
		14'b11110010100100: color_data = 12'b010000000000;
		14'b11110010100101: color_data = 12'b001000000000;
		14'b11110010100110: color_data = 12'b001000000000;
		14'b11110010100111: color_data = 12'b010000000000;
		14'b11110010101000: color_data = 12'b010000000000;
		14'b11110010101001: color_data = 12'b010000000000;
		14'b11110010101010: color_data = 12'b010000000000;
		14'b11110010101011: color_data = 12'b010000000000;
		14'b11110010101100: color_data = 12'b010000000000;
		14'b11110010101101: color_data = 12'b001000000000;
		14'b11110010101110: color_data = 12'b001000000000;
		14'b11110010101111: color_data = 12'b001000000000;
		14'b11110011100111: color_data = 12'b001000000000;
		14'b11110011101000: color_data = 12'b001000000000;
		14'b11110011101001: color_data = 12'b001000000000;
		14'b11110011101010: color_data = 12'b001000000000;
		14'b11110011101011: color_data = 12'b001000000000;
		14'b11110011101100: color_data = 12'b001000000000;
		14'b11110011101101: color_data = 12'b001000000000;
		14'b11110011101110: color_data = 12'b010000000000;
		14'b11110011101111: color_data = 12'b010000000000;
		14'b11110011110000: color_data = 12'b010000000000;
		14'b11110011110001: color_data = 12'b010000000000;
		14'b11110011110010: color_data = 12'b001000000000;
		14'b11110100010001: color_data = 12'b001000000000;
		14'b11110100010110: color_data = 12'b001000000000;
		14'b11110100010111: color_data = 12'b001000000000;
		14'b11110100011000: color_data = 12'b010000000000;
		14'b11110100011001: color_data = 12'b010000000000;
		14'b11110100011010: color_data = 12'b010000000000;
		14'b11110100011011: color_data = 12'b010000000000;
		14'b11110100011100: color_data = 12'b010000000000;
		14'b11110100011101: color_data = 12'b010000000000;
		14'b11110100011110: color_data = 12'b010000000000;
		14'b11110100011111: color_data = 12'b010000000000;
		14'b11110100100000: color_data = 12'b010000000000;
		14'b11110100100001: color_data = 12'b010000000000;
		14'b11110100100010: color_data = 12'b010000000000;
		14'b11110100100011: color_data = 12'b010000000000;
		14'b11110100100100: color_data = 12'b010000000000;
		14'b11110100100101: color_data = 12'b010000000000;
		14'b11110100100110: color_data = 12'b010000000000;
		14'b11110100100111: color_data = 12'b010000000000;
		14'b11110100101000: color_data = 12'b010000000000;
		14'b11110100101001: color_data = 12'b010000000000;
		14'b11110100101010: color_data = 12'b010000000000;
		14'b11110100101011: color_data = 12'b001000000000;
		14'b11110100101100: color_data = 12'b001000000000;
		14'b11110100101101: color_data = 12'b001000000000;
		14'b11110100101110: color_data = 12'b001000000000;
		14'b11110101100011: color_data = 12'b001000000000;
		14'b11110101100100: color_data = 12'b001000000000;
		14'b11110101100101: color_data = 12'b001000000000;
		14'b11110101100110: color_data = 12'b001000000000;
		14'b11110101100111: color_data = 12'b001000000000;
		14'b11110101101000: color_data = 12'b001000000000;
		14'b11110101101001: color_data = 12'b001000000000;
		14'b11110101101010: color_data = 12'b001000000000;
		14'b11110101101011: color_data = 12'b001000000000;
		14'b11110101101100: color_data = 12'b001000000000;
		14'b11110101101101: color_data = 12'b010000000000;
		14'b11110101101110: color_data = 12'b010000000000;
		14'b11110101101111: color_data = 12'b010000000000;
		14'b11110101110000: color_data = 12'b010000000000;
		14'b11110101110001: color_data = 12'b001000000000;
		14'b11110110001000: color_data = 12'b001000000000;
		14'b11110110001001: color_data = 12'b001000000000;
		14'b11110110010001: color_data = 12'b001000000000;
		14'b11110110010010: color_data = 12'b001000000000;
		14'b11110110010011: color_data = 12'b001000000000;
		14'b11110110010100: color_data = 12'b001000000000;
		14'b11110110010101: color_data = 12'b001000000000;
		14'b11110110010110: color_data = 12'b001000000000;
		14'b11110110010111: color_data = 12'b001000000000;
		14'b11110110011000: color_data = 12'b001000000000;
		14'b11110110011001: color_data = 12'b001000000000;
		14'b11110110011010: color_data = 12'b001000000000;
		14'b11110110011011: color_data = 12'b010000000000;
		14'b11110110011100: color_data = 12'b010000000000;
		14'b11110110011101: color_data = 12'b010000000000;
		14'b11110110011110: color_data = 12'b010000000000;
		14'b11110110011111: color_data = 12'b010000000000;
		14'b11110110100000: color_data = 12'b010000000000;
		14'b11110110100001: color_data = 12'b010000000000;
		14'b11110110100010: color_data = 12'b010000000000;
		14'b11110110100011: color_data = 12'b010000000000;
		14'b11110110100100: color_data = 12'b010000000000;
		14'b11110110100101: color_data = 12'b010000000000;
		14'b11110110100110: color_data = 12'b010000000000;
		14'b11110110100111: color_data = 12'b001000000000;
		14'b11110110101000: color_data = 12'b001000000000;
		14'b11110110101001: color_data = 12'b001000000000;
		14'b11110110101010: color_data = 12'b001000000000;
		14'b11110110101011: color_data = 12'b001000000000;
		14'b11110111100000: color_data = 12'b001000000000;
		14'b11110111100001: color_data = 12'b001000000000;
		14'b11110111100010: color_data = 12'b001000000000;
		14'b11110111100011: color_data = 12'b001000000000;
		14'b11110111100100: color_data = 12'b001000000000;
		14'b11110111100101: color_data = 12'b001000000000;
		14'b11110111100110: color_data = 12'b001000000000;
		14'b11110111100111: color_data = 12'b001000000000;
		14'b11110111101000: color_data = 12'b001000000000;
		14'b11110111101001: color_data = 12'b001000000000;
		14'b11110111101010: color_data = 12'b001000000000;
		14'b11110111101011: color_data = 12'b001000000000;
		14'b11110111101100: color_data = 12'b010000000000;
		14'b11110111101101: color_data = 12'b010000000000;
		14'b11110111101110: color_data = 12'b010000000000;
		14'b11110111101111: color_data = 12'b010000000000;
		14'b11110111110000: color_data = 12'b001000000000;
		14'b11111000001001: color_data = 12'b001000000000;
		14'b11111000001010: color_data = 12'b001000000000;
		14'b11111000001011: color_data = 12'b001000000000;
		14'b11111000010001: color_data = 12'b001000000000;
		14'b11111000010010: color_data = 12'b001000000000;
		14'b11111000010011: color_data = 12'b001000000000;
		14'b11111000010100: color_data = 12'b001000000000;
		14'b11111000010101: color_data = 12'b001000000000;
		14'b11111000010110: color_data = 12'b001000000000;
		14'b11111000010111: color_data = 12'b001000000000;
		14'b11111000011000: color_data = 12'b010000000000;
		14'b11111000011001: color_data = 12'b010000000000;
		14'b11111000011010: color_data = 12'b010000000000;
		14'b11111000011011: color_data = 12'b010000000000;
		14'b11111000011100: color_data = 12'b010000000000;
		14'b11111000011101: color_data = 12'b010000000000;
		14'b11111000011110: color_data = 12'b001000000000;
		14'b11111000011111: color_data = 12'b001000000000;
		14'b11111000100000: color_data = 12'b001000000000;
		14'b11111000100001: color_data = 12'b001000000000;
		14'b11111000100010: color_data = 12'b001000000000;
		14'b11111000100011: color_data = 12'b001000000000;
		14'b11111000100100: color_data = 12'b001000000000;
		14'b11111000100101: color_data = 12'b001000000000;
		14'b11111000100111: color_data = 12'b001000000000;
		14'b11111000101000: color_data = 12'b001000000000;
		14'b11111000101001: color_data = 12'b001000000000;
		14'b11111000101010: color_data = 12'b001000000000;
		14'b11111000101011: color_data = 12'b001000000000;
		14'b11111001001111: color_data = 12'b001000000000;
		14'b11111001010000: color_data = 12'b001000000000;
		14'b11111001011101: color_data = 12'b001000000000;
		14'b11111001011110: color_data = 12'b001000000000;
		14'b11111001011111: color_data = 12'b001000000000;
		14'b11111001100000: color_data = 12'b001000000000;
		14'b11111001100001: color_data = 12'b001000000000;
		14'b11111001100010: color_data = 12'b001000000000;
		14'b11111001100011: color_data = 12'b001000000000;
		14'b11111001100100: color_data = 12'b001000000000;
		14'b11111001100101: color_data = 12'b001000000000;
		14'b11111001100110: color_data = 12'b001000000000;
		14'b11111001100111: color_data = 12'b001000000000;
		14'b11111001101000: color_data = 12'b001000000000;
		14'b11111001101001: color_data = 12'b001000000000;
		14'b11111001101010: color_data = 12'b010000000000;
		14'b11111001101011: color_data = 12'b010000000000;
		14'b11111001101100: color_data = 12'b010000000000;
		14'b11111001101101: color_data = 12'b001000000000;
		14'b11111001101110: color_data = 12'b001000000000;
		14'b11111001101111: color_data = 12'b001000000000;
		14'b11111001110000: color_data = 12'b001000000000;
		14'b11111010001100: color_data = 12'b001000000000;
		14'b11111010001101: color_data = 12'b001000000000;
		14'b11111010001110: color_data = 12'b001000000000;
		14'b11111010001111: color_data = 12'b001000000000;
		14'b11111010010000: color_data = 12'b001000000000;
		14'b11111010010001: color_data = 12'b001000000000;
		14'b11111010010010: color_data = 12'b001000000000;
		14'b11111010010011: color_data = 12'b001000000000;
		14'b11111010010100: color_data = 12'b001000000000;
		14'b11111010010101: color_data = 12'b001000000000;
		14'b11111010010110: color_data = 12'b001000000000;
		14'b11111010010111: color_data = 12'b001000000000;
		14'b11111010011000: color_data = 12'b001000000000;
		14'b11111010011001: color_data = 12'b001000000000;
		14'b11111010011010: color_data = 12'b001000000000;
		14'b11111010011011: color_data = 12'b001000000000;
		14'b11111010011100: color_data = 12'b001000000000;
		14'b11111010011101: color_data = 12'b001000000000;
		14'b11111010011110: color_data = 12'b001000000000;
		14'b11111010011111: color_data = 12'b001000000000;
		14'b11111010100000: color_data = 12'b001000000000;
		14'b11111010100001: color_data = 12'b001000000000;
		14'b11111010100010: color_data = 12'b001000000000;
		14'b11111010100011: color_data = 12'b001000000000;
		14'b11111010100100: color_data = 12'b001000000000;
		14'b11111010100101: color_data = 12'b001000000000;
		14'b11111011010000: color_data = 12'b001000000000;
		14'b11111011010001: color_data = 12'b010000000000;
		14'b11111011010010: color_data = 12'b001000000000;
		14'b11111011010011: color_data = 12'b001000000000;
		14'b11111011010100: color_data = 12'b001000000000;
		14'b11111011010101: color_data = 12'b001000000000;
		14'b11111011010110: color_data = 12'b001000000000;
		14'b11111011010111: color_data = 12'b001000000000;
		14'b11111011011000: color_data = 12'b001000000000;
		14'b11111011011001: color_data = 12'b001000000000;
		14'b11111011011010: color_data = 12'b001000000000;
		14'b11111011011011: color_data = 12'b001000000000;
		14'b11111011011100: color_data = 12'b001000000000;
		14'b11111011011101: color_data = 12'b010000000000;
		14'b11111011011110: color_data = 12'b010000000000;
		14'b11111011011111: color_data = 12'b010000000000;
		14'b11111011100000: color_data = 12'b010000000000;
		14'b11111011100001: color_data = 12'b010000000000;
		14'b11111011100010: color_data = 12'b010000000000;
		14'b11111011100011: color_data = 12'b010000000000;
		14'b11111011100100: color_data = 12'b001000000000;
		14'b11111011100101: color_data = 12'b001000000000;
		14'b11111011100110: color_data = 12'b001000000000;
		14'b11111011100111: color_data = 12'b001000000000;
		14'b11111011101000: color_data = 12'b010000000000;
		14'b11111011101001: color_data = 12'b010000000000;
		14'b11111011101010: color_data = 12'b010000000000;
		14'b11111011101011: color_data = 12'b001000000000;
		14'b11111011101100: color_data = 12'b001000000000;
		14'b11111011101101: color_data = 12'b001000000000;
		14'b11111011101110: color_data = 12'b001000000000;
		14'b11111011101111: color_data = 12'b001000000000;
		14'b11111011111111: color_data = 12'b001000000000;
		14'b11111100010001: color_data = 12'b001000000000;
		14'b11111100010010: color_data = 12'b001000000000;
		14'b11111100010011: color_data = 12'b001000000000;
		14'b11111100010100: color_data = 12'b001000000000;
		14'b11111100010101: color_data = 12'b001000000000;
		14'b11111100010110: color_data = 12'b001000000000;
		14'b11111100010111: color_data = 12'b001000000000;
		14'b11111100011000: color_data = 12'b001000000000;
		14'b11111100111100: color_data = 12'b001000000000;
		14'b11111100111101: color_data = 12'b001000000000;
		14'b11111100111110: color_data = 12'b001000000000;
		14'b11111101010001: color_data = 12'b001000000000;
		14'b11111101010010: color_data = 12'b010000000000;
		14'b11111101010011: color_data = 12'b010000000000;
		14'b11111101010100: color_data = 12'b010000000000;
		14'b11111101010101: color_data = 12'b010000000000;
		14'b11111101010110: color_data = 12'b010000000000;
		14'b11111101010111: color_data = 12'b010000000000;
		14'b11111101011000: color_data = 12'b010000000000;
		14'b11111101011001: color_data = 12'b010000000000;
		14'b11111101011010: color_data = 12'b010000000000;
		14'b11111101011011: color_data = 12'b010000000000;
		14'b11111101011100: color_data = 12'b010000000000;
		14'b11111101011101: color_data = 12'b010000000000;
		14'b11111101011110: color_data = 12'b010000000000;
		14'b11111101011111: color_data = 12'b010000000000;
		14'b11111101100000: color_data = 12'b010000000000;
		14'b11111101100001: color_data = 12'b010000000000;
		14'b11111101100010: color_data = 12'b010000000000;
		14'b11111101100011: color_data = 12'b010000000000;
		14'b11111101100100: color_data = 12'b001000000000;
		14'b11111101100101: color_data = 12'b001000000000;
		14'b11111101100110: color_data = 12'b001000000000;
		14'b11111101100111: color_data = 12'b001000000000;
		14'b11111101101000: color_data = 12'b001000000000;
		14'b11111101101001: color_data = 12'b001000000000;
		14'b11111101101010: color_data = 12'b001000000000;
		14'b11111110111111: color_data = 12'b001000000000;
		14'b11111111000000: color_data = 12'b001000000000;
		14'b11111111010011: color_data = 12'b001000000000;
		14'b11111111010100: color_data = 12'b001000000000;
		14'b11111111010101: color_data = 12'b001000000000;
		14'b11111111010110: color_data = 12'b001000000000;
		14'b11111111010111: color_data = 12'b001000000000;
		14'b11111111011000: color_data = 12'b010000000000;
		14'b11111111011001: color_data = 12'b010000000000;
		14'b11111111011010: color_data = 12'b010000000000;
		14'b11111111011011: color_data = 12'b010000000000;
		14'b11111111011100: color_data = 12'b010000000000;
		14'b11111111011101: color_data = 12'b010000000000;
		14'b11111111011110: color_data = 12'b010000000000;
		14'b11111111011111: color_data = 12'b010000000000;
		14'b11111111100000: color_data = 12'b010000000000;
		14'b11111111100001: color_data = 12'b010000000000;
		14'b11111111100010: color_data = 12'b010000000000;
		14'b11111111100011: color_data = 12'b010000000000;
		14'b11111111100100: color_data = 12'b010000000000;
		14'b11111111100101: color_data = 12'b001000000000;
		14'b11111111100110: color_data = 12'b001000000000;
		14'b11111111100111: color_data = 12'b001000000000;
		default: color_data = 12'b000000000000;
	endcase
endmodule