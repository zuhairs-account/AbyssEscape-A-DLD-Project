module death_1_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);
parameter Z = 12'b111111111111;
		
	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		19'b0110101100100111111: color_data = Z;
		19'b0110101100101000000: color_data = Z;
		19'b0110101100101000001: color_data = Z;
		19'b0110101100101000010: color_data = Z;
		19'b0110101100101000011: color_data = Z;
		19'b0110101110100111100: color_data = Z;
		19'b0110101110100111101: color_data = Z;
		19'b0110101110100111110: color_data = Z;
		19'b0110101110100111111: color_data = Z;
		19'b0110101110101000000: color_data = Z;
		19'b0110101110101000001: color_data = Z;
		19'b0110101110101000010: color_data = Z;
		19'b0110101110101000011: color_data = Z;
		19'b0110101110101000100: color_data = Z;
		19'b0110101110101000101: color_data = Z;
		19'b0110101110101000110: color_data = Z;
		19'b0110110000100111010: color_data = Z;
		19'b0110110000100111011: color_data = Z;
		19'b0110110000100111100: color_data = Z;
		19'b0110110000100111101: color_data = Z;
		19'b0110110000100111110: color_data = Z;
		19'b0110110000100111111: color_data = Z;
		19'b0110110000101000000: color_data = Z;
		19'b0110110000101000001: color_data = Z;
		19'b0110110000101000010: color_data = Z;
		19'b0110110000101000011: color_data = Z;
		19'b0110110000101000100: color_data = Z;
		19'b0110110000101000101: color_data = Z;
		19'b0110110000101000110: color_data = Z;
		19'b0110110000101000111: color_data = Z;
		19'b0110110000101001000: color_data = Z;
		19'b0110110010100111000: color_data = Z;
		19'b0110110010100111001: color_data = Z;
		19'b0110110010100111010: color_data = Z;
		19'b0110110010100111011: color_data = Z;
		19'b0110110010100111100: color_data = Z;
		19'b0110110010100111101: color_data = Z;
		19'b0110110010100111110: color_data = Z;
		19'b0110110010100111111: color_data = Z;
		19'b0110110010101000000: color_data = Z;
		19'b0110110010101000001: color_data = Z;
		19'b0110110010101000010: color_data = Z;
		19'b0110110010101000011: color_data = Z;
		19'b0110110010101000100: color_data = Z;
		19'b0110110010101000101: color_data = Z;
		19'b0110110010101000110: color_data = Z;
		19'b0110110010101000111: color_data = Z;
		19'b0110110010101001000: color_data = Z;
		19'b0110110010101001001: color_data = Z;
		19'b0110110100100110111: color_data = Z;
		19'b0110110100100111000: color_data = Z;
		19'b0110110100100111001: color_data = Z;
		19'b0110110100100111010: color_data = Z;
		19'b0110110100100111011: color_data = Z;
		19'b0110110100100111100: color_data = Z;
		19'b0110110100100111101: color_data = Z;
		19'b0110110100100111110: color_data = Z;
		19'b0110110100100111111: color_data = Z;
		19'b0110110100101000000: color_data = Z;
		19'b0110110100101000001: color_data = Z;
		19'b0110110100101000010: color_data = Z;
		19'b0110110100101000011: color_data = Z;
		19'b0110110100101000100: color_data = Z;
		19'b0110110100101000101: color_data = Z;
		19'b0110110100101000110: color_data = Z;
		19'b0110110100101000111: color_data = Z;
		19'b0110110100101001000: color_data = Z;
		19'b0110110100101001001: color_data = Z;
		19'b0110110100101001010: color_data = Z;
		19'b0110110110100110110: color_data = Z;
		19'b0110110110100110111: color_data = Z;
		19'b0110110110100111000: color_data = Z;
		19'b0110110110100111001: color_data = Z;
		19'b0110110110100111010: color_data = Z;
		19'b0110110110100111011: color_data = Z;
		19'b0110110110100111100: color_data = Z;
		19'b0110110110100111101: color_data = Z;
		19'b0110110110100111110: color_data = Z;
		19'b0110110110100111111: color_data = Z;
		19'b0110110110101000000: color_data = Z;
		19'b0110110110101000001: color_data = Z;
		19'b0110110110101000010: color_data = Z;
		19'b0110110110101000011: color_data = Z;
		19'b0110110110101000100: color_data = Z;
		19'b0110110110101000101: color_data = Z;
		19'b0110110110101000110: color_data = Z;
		19'b0110110110101000111: color_data = Z;
		19'b0110110110101001000: color_data = Z;
		19'b0110110110101001001: color_data = Z;
		19'b0110110110101001010: color_data = Z;
		19'b0110110110101001011: color_data = Z;
		19'b0110111000100110101: color_data = Z;
		19'b0110111000100110110: color_data = Z;
		19'b0110111000100110111: color_data = Z;
		19'b0110111000100111000: color_data = Z;
		19'b0110111000100111001: color_data = Z;
		19'b0110111000100111010: color_data = Z;
		19'b0110111000100111011: color_data = Z;
		19'b0110111000100111100: color_data = Z;
		19'b0110111000100111101: color_data = Z;
		19'b0110111000100111110: color_data = Z;
		19'b0110111000100111111: color_data = Z;
		19'b0110111000101000000: color_data = Z;
		19'b0110111000101000001: color_data = Z;
		19'b0110111000101000010: color_data = Z;
		19'b0110111000101000011: color_data = Z;
		19'b0110111000101000100: color_data = Z;
		19'b0110111000101000101: color_data = Z;
		19'b0110111000101000110: color_data = Z;
		19'b0110111000101000111: color_data = Z;
		19'b0110111000101001000: color_data = Z;
		19'b0110111000101001001: color_data = Z;
		19'b0110111000101001010: color_data = Z;
		19'b0110111000101001011: color_data = Z;
		19'b0110111000101001100: color_data = Z;
		19'b0110111000101001101: color_data = Z;
		19'b0110111010100110100: color_data = Z;
		19'b0110111010100110101: color_data = Z;
		19'b0110111010100110110: color_data = Z;
		19'b0110111010100110111: color_data = Z;
		19'b0110111010100111000: color_data = Z;
		19'b0110111010100111001: color_data = Z;
		19'b0110111010100111010: color_data = Z;
		19'b0110111010100111011: color_data = Z;
		19'b0110111010100111100: color_data = Z;
		19'b0110111010100111101: color_data = Z;
		19'b0110111010100111110: color_data = Z;
		19'b0110111010100111111: color_data = Z;
		19'b0110111010101000000: color_data = Z;
		19'b0110111010101000001: color_data = Z;
		19'b0110111010101000010: color_data = Z;
		19'b0110111010101000011: color_data = Z;
		19'b0110111010101000100: color_data = Z;
		19'b0110111010101000101: color_data = Z;
		19'b0110111010101000110: color_data = Z;
		19'b0110111010101000111: color_data = Z;
		19'b0110111010101001000: color_data = Z;
		19'b0110111010101001001: color_data = Z;
		19'b0110111010101001010: color_data = Z;
		19'b0110111010101001011: color_data = Z;
		19'b0110111010101001100: color_data = Z;
		19'b0110111010101001101: color_data = Z;
		19'b0110111010101001110: color_data = Z;
		19'b0110111100100110010: color_data = Z;
		19'b0110111100100110011: color_data = Z;
		19'b0110111100100110100: color_data = Z;
		19'b0110111100100110101: color_data = Z;
		19'b0110111100100110110: color_data = Z;
		19'b0110111100100110111: color_data = Z;
		19'b0110111100100111000: color_data = Z;
		19'b0110111100100111001: color_data = Z;
		19'b0110111100100111010: color_data = Z;
		19'b0110111100100111011: color_data = Z;
		19'b0110111100100111100: color_data = Z;
		19'b0110111100100111101: color_data = Z;
		19'b0110111100100111110: color_data = Z;
		19'b0110111100100111111: color_data = Z;
		19'b0110111100101000000: color_data = Z;
		19'b0110111100101000001: color_data = Z;
		19'b0110111100101000010: color_data = Z;
		19'b0110111100101000011: color_data = Z;
		19'b0110111100101000100: color_data = Z;
		19'b0110111100101000101: color_data = Z;
		19'b0110111100101000110: color_data = Z;
		19'b0110111100101000111: color_data = Z;
		19'b0110111100101001000: color_data = Z;
		19'b0110111100101001001: color_data = Z;
		19'b0110111100101001010: color_data = Z;
		19'b0110111100101001011: color_data = Z;
		19'b0110111100101001100: color_data = Z;
		19'b0110111100101001101: color_data = Z;
		19'b0110111100101001110: color_data = Z;
		19'b0110111100101001111: color_data = Z;
		19'b0110111110100110000: color_data = Z;
		19'b0110111110100110001: color_data = Z;
		19'b0110111110100110010: color_data = Z;
		19'b0110111110100110011: color_data = Z;
		19'b0110111110100110100: color_data = Z;
		19'b0110111110100110101: color_data = Z;
		19'b0110111110100110110: color_data = Z;
		19'b0110111110100110111: color_data = Z;
		19'b0110111110100111000: color_data = Z;
		19'b0110111110100111001: color_data = Z;
		19'b0110111110100111010: color_data = Z;
		19'b0110111110100111011: color_data = Z;
		19'b0110111110100111100: color_data = Z;
		19'b0110111110100111101: color_data = Z;
		19'b0110111110100111110: color_data = Z;
		19'b0110111110100111111: color_data = Z;
		19'b0110111110101000000: color_data = Z;
		19'b0110111110101000001: color_data = Z;
		19'b0110111110101000010: color_data = Z;
		19'b0110111110101000011: color_data = Z;
		19'b0110111110101000100: color_data = Z;
		19'b0110111110101000101: color_data = Z;
		19'b0110111110101000110: color_data = Z;
		19'b0110111110101000111: color_data = Z;
		19'b0110111110101001000: color_data = Z;
		19'b0110111110101001001: color_data = Z;
		19'b0110111110101001010: color_data = Z;
		19'b0110111110101001011: color_data = Z;
		19'b0110111110101001100: color_data = Z;
		19'b0110111110101001101: color_data = Z;
		19'b0110111110101001110: color_data = Z;
		19'b0110111110101001111: color_data = Z;
		19'b0111000000100101111: color_data = Z;
		19'b0111000000100110000: color_data = Z;
		19'b0111000000100110001: color_data = Z;
		19'b0111000000100110010: color_data = Z;
		19'b0111000000100110011: color_data = Z;
		19'b0111000000100110100: color_data = Z;
		19'b0111000000100110101: color_data = Z;
		19'b0111000000100110110: color_data = Z;
		19'b0111000000100110111: color_data = Z;
		19'b0111000000100111000: color_data = Z;
		19'b0111000000100111001: color_data = Z;
		19'b0111000000100111010: color_data = Z;
		19'b0111000000100111011: color_data = Z;
		19'b0111000000100111100: color_data = Z;
		19'b0111000000100111101: color_data = Z;
		19'b0111000000100111110: color_data = Z;
		19'b0111000000100111111: color_data = Z;
		19'b0111000000101000000: color_data = Z;
		19'b0111000000101000001: color_data = Z;
		19'b0111000000101000010: color_data = Z;
		19'b0111000000101000011: color_data = Z;
		19'b0111000000101000100: color_data = Z;
		19'b0111000000101000101: color_data = Z;
		19'b0111000000101000110: color_data = Z;
		19'b0111000000101000111: color_data = Z;
		19'b0111000000101001000: color_data = Z;
		19'b0111000000101001001: color_data = Z;
		19'b0111000000101001010: color_data = Z;
		19'b0111000000101001011: color_data = Z;
		19'b0111000000101001100: color_data = Z;
		19'b0111000000101001101: color_data = Z;
		19'b0111000000101001110: color_data = Z;
		19'b0111000000101001111: color_data = Z;
		19'b0111000010100101111: color_data = Z;
		19'b0111000010100110000: color_data = Z;
		19'b0111000010100110001: color_data = Z;
		19'b0111000010100110010: color_data = Z;
		19'b0111000010100110011: color_data = Z;
		19'b0111000010100110100: color_data = Z;
		19'b0111000010100110101: color_data = Z;
		19'b0111000010100110110: color_data = Z;
		19'b0111000010100110111: color_data = Z;
		19'b0111000010100111000: color_data = Z;
		19'b0111000010100111001: color_data = Z;
		19'b0111000010100111010: color_data = Z;
		19'b0111000010100111011: color_data = Z;
		19'b0111000010100111100: color_data = Z;
		19'b0111000010100111101: color_data = Z;
		19'b0111000010100111110: color_data = Z;
		19'b0111000010100111111: color_data = Z;
		19'b0111000010101000000: color_data = Z;
		19'b0111000010101000001: color_data = Z;
		19'b0111000010101000010: color_data = Z;
		19'b0111000010101000011: color_data = Z;
		19'b0111000010101000100: color_data = Z;
		19'b0111000010101000101: color_data = Z;
		19'b0111000010101000110: color_data = Z;
		19'b0111000010101000111: color_data = Z;
		19'b0111000010101001000: color_data = Z;
		19'b0111000010101001001: color_data = Z;
		19'b0111000010101001010: color_data = Z;
		19'b0111000010101001011: color_data = Z;
		19'b0111000010101001100: color_data = Z;
		19'b0111000010101001101: color_data = Z;
		19'b0111000010101001110: color_data = Z;
		19'b0111000010101001111: color_data = Z;
		19'b0111000100100101110: color_data = Z;
		19'b0111000100100101111: color_data = Z;
		19'b0111000100100110000: color_data = Z;
		19'b0111000100100110001: color_data = Z;
		19'b0111000100100110010: color_data = Z;
		19'b0111000100100110011: color_data = Z;
		19'b0111000100100110100: color_data = Z;
		19'b0111000100100110101: color_data = Z;
		19'b0111000100100110110: color_data = Z;
		19'b0111000100100110111: color_data = Z;
		19'b0111000100100111000: color_data = Z;
		19'b0111000100100111001: color_data = Z;
		19'b0111000100100111010: color_data = Z;
		19'b0111000100100111011: color_data = Z;
		19'b0111000100100111100: color_data = Z;
		19'b0111000100100111101: color_data = Z;
		19'b0111000100100111110: color_data = Z;
		19'b0111000100100111111: color_data = Z;
		19'b0111000100101000000: color_data = Z;
		19'b0111000100101000001: color_data = Z;
		19'b0111000100101000010: color_data = Z;
		19'b0111000100101000011: color_data = Z;
		19'b0111000100101000100: color_data = Z;
		19'b0111000100101000101: color_data = Z;
		19'b0111000100101000110: color_data = Z;
		19'b0111000100101000111: color_data = Z;
		19'b0111000100101001100: color_data = Z;
		19'b0111000100101001101: color_data = Z;
		19'b0111000100101001110: color_data = Z;
		19'b0111000100101001111: color_data = Z;
		19'b0111000100101010000: color_data = Z;
		19'b0111000110100101110: color_data = Z;
		19'b0111000110100101111: color_data = Z;
		19'b0111000110100110000: color_data = Z;
		19'b0111000110100110001: color_data = Z;
		19'b0111000110100110010: color_data = Z;
		19'b0111000110100110011: color_data = Z;
		19'b0111000110100110100: color_data = Z;
		19'b0111000110100111000: color_data = Z;
		19'b0111000110100111001: color_data = Z;
		19'b0111000110100111010: color_data = Z;
		19'b0111000110100111011: color_data = Z;
		19'b0111000110100111100: color_data = Z;
		19'b0111000110100111101: color_data = Z;
		19'b0111000110100111110: color_data = Z;
		19'b0111000110100111111: color_data = Z;
		19'b0111000110101000000: color_data = Z;
		19'b0111000110101000001: color_data = Z;
		19'b0111000110101000010: color_data = Z;
		19'b0111000110101000011: color_data = Z;
		19'b0111000110101000100: color_data = Z;
		19'b0111000110101000101: color_data = Z;
		19'b0111000110101000110: color_data = Z;
		19'b0111000110101001101: color_data = Z;
		19'b0111000110101001110: color_data = Z;
		19'b0111000110101001111: color_data = Z;
		19'b0111000110101010000: color_data = Z;
		19'b0111001000100101110: color_data = Z;
		19'b0111001000100101111: color_data = Z;
		19'b0111001000100110000: color_data = Z;
		19'b0111001000100110001: color_data = Z;
		19'b0111001000100110010: color_data = Z;
		19'b0111001000100111001: color_data = Z;
		19'b0111001000100111010: color_data = Z;
		19'b0111001000100111011: color_data = Z;
		19'b0111001000100111100: color_data = Z;
		19'b0111001000100111101: color_data = Z;
		19'b0111001000100111110: color_data = Z;
		19'b0111001000100111111: color_data = Z;
		19'b0111001000101000000: color_data = Z;
		19'b0111001000101000001: color_data = Z;
		19'b0111001000101000010: color_data = Z;
		19'b0111001000101000011: color_data = Z;
		19'b0111001000101000100: color_data = Z;
		19'b0111001000101000101: color_data = Z;
		19'b0111001000101001110: color_data = Z;
		19'b0111001000101001111: color_data = Z;
		19'b0111001000101010000: color_data = Z;
		19'b0111001010100101110: color_data = Z;
		19'b0111001010100101111: color_data = Z;
		19'b0111001010100110000: color_data = Z;
		19'b0111001010100110001: color_data = Z;
		19'b0111001010100111011: color_data = Z;
		19'b0111001010100111100: color_data = Z;
		19'b0111001010100111101: color_data = Z;
		19'b0111001010100111110: color_data = Z;
		19'b0111001010100111111: color_data = Z;
		19'b0111001010101000000: color_data = Z;
		19'b0111001010101000001: color_data = Z;
		19'b0111001010101000010: color_data = Z;
		19'b0111001010101000011: color_data = Z;
		19'b0111001010101000100: color_data = Z;
		19'b0111001010101000101: color_data = Z;
		19'b0111001010101001110: color_data = Z;
		19'b0111001010101001111: color_data = Z;
		19'b0111001010101010000: color_data = Z;
		19'b0111001100100101110: color_data = Z;
		19'b0111001100100101111: color_data = Z;
		19'b0111001100100110000: color_data = Z;
		19'b0111001100100110001: color_data = Z;
		19'b0111001100100111011: color_data = Z;
		19'b0111001100100111100: color_data = Z;
		19'b0111001100100111101: color_data = Z;
		19'b0111001100100111110: color_data = Z;
		19'b0111001100100111111: color_data = Z;
		19'b0111001100101000000: color_data = Z;
		19'b0111001100101000001: color_data = Z;
		19'b0111001100101000010: color_data = Z;
		19'b0111001100101000011: color_data = Z;
		19'b0111001100101000100: color_data = Z;
		19'b0111001100101000101: color_data = Z;
		19'b0111001100101001110: color_data = Z;
		19'b0111001100101001111: color_data = Z;
		19'b0111001100101010000: color_data = Z;
		19'b0111001110100101110: color_data = Z;
		19'b0111001110100101111: color_data = Z;
		19'b0111001110100110000: color_data = Z;
		19'b0111001110100111011: color_data = Z;
		19'b0111001110100111100: color_data = Z;
		19'b0111001110100111101: color_data = Z;
		19'b0111001110100111110: color_data = Z;
		19'b0111001110100111111: color_data = Z;
		19'b0111001110101000000: color_data = Z;
		19'b0111001110101000001: color_data = Z;
		19'b0111001110101000010: color_data = Z;
		19'b0111001110101000011: color_data = Z;
		19'b0111001110101000100: color_data = Z;
		19'b0111001110101000101: color_data = Z;
		19'b0111001110101001110: color_data = Z;
		19'b0111001110101001111: color_data = Z;
		19'b0111001110101010000: color_data = Z;
		19'b0111010000100101110: color_data = Z;
		19'b0111010000100101111: color_data = Z;
		19'b0111010000100110000: color_data = Z;
		19'b0111010000100111011: color_data = Z;
		19'b0111010000100111100: color_data = Z;
		19'b0111010000100111101: color_data = Z;
		19'b0111010000100111110: color_data = Z;
		19'b0111010000100111111: color_data = Z;
		19'b0111010000101000000: color_data = Z;
		19'b0111010000101000001: color_data = Z;
		19'b0111010000101000010: color_data = Z;
		19'b0111010000101000011: color_data = Z;
		19'b0111010000101000100: color_data = Z;
		19'b0111010000101000101: color_data = Z;
		19'b0111010000101001110: color_data = Z;
		19'b0111010000101001111: color_data = Z;
		19'b0111010000101010000: color_data = Z;
		19'b0111010010100101110: color_data = Z;
		19'b0111010010100101111: color_data = Z;
		19'b0111010010100110000: color_data = Z;
		19'b0111010010100111011: color_data = Z;
		19'b0111010010100111100: color_data = Z;
		19'b0111010010100111101: color_data = Z;
		19'b0111010010100111110: color_data = Z;
		19'b0111010010100111111: color_data = Z;
		19'b0111010010101000000: color_data = Z;
		19'b0111010010101000001: color_data = Z;
		19'b0111010010101000010: color_data = Z;
		19'b0111010010101000011: color_data = Z;
		19'b0111010010101000100: color_data = Z;
		19'b0111010010101000101: color_data = Z;
		19'b0111010010101000110: color_data = Z;
		19'b0111010010101001110: color_data = Z;
		19'b0111010010101001111: color_data = Z;
		19'b0111010010101010000: color_data = Z;
		19'b0111010100100101110: color_data = Z;
		19'b0111010100100101111: color_data = Z;
		19'b0111010100100110000: color_data = Z;
		19'b0111010100100110001: color_data = Z;
		19'b0111010100100111010: color_data = Z;
		19'b0111010100100111011: color_data = Z;
		19'b0111010100100111100: color_data = Z;
		19'b0111010100100111101: color_data = Z;
		19'b0111010100100111110: color_data = Z;
		19'b0111010100100111111: color_data = Z;
		19'b0111010100101000000: color_data = Z;
		19'b0111010100101000001: color_data = Z;
		19'b0111010100101000010: color_data = Z;
		19'b0111010100101000011: color_data = Z;
		19'b0111010100101000100: color_data = Z;
		19'b0111010100101000101: color_data = Z;
		19'b0111010100101000110: color_data = Z;
		19'b0111010100101000111: color_data = Z;
		19'b0111010100101001101: color_data = Z;
		19'b0111010100101001110: color_data = Z;
		19'b0111010100101001111: color_data = Z;
		19'b0111010100101010000: color_data = Z;
		19'b0111010110100101110: color_data = Z;
		19'b0111010110100101111: color_data = Z;
		19'b0111010110100110000: color_data = Z;
		19'b0111010110100110001: color_data = Z;
		19'b0111010110100111010: color_data = Z;
		19'b0111010110100111011: color_data = Z;
		19'b0111010110100111100: color_data = Z;
		19'b0111010110100111101: color_data = Z;
		19'b0111010110100111110: color_data = Z;
		19'b0111010110100111111: color_data = Z;
		19'b0111010110101000000: color_data = Z;
		19'b0111010110101000001: color_data = Z;
		19'b0111010110101000010: color_data = Z;
		19'b0111010110101000011: color_data = Z;
		19'b0111010110101000100: color_data = Z;
		19'b0111010110101000101: color_data = Z;
		19'b0111010110101000110: color_data = Z;
		19'b0111010110101000111: color_data = Z;
		19'b0111010110101001110: color_data = Z;
		19'b0111010110101001111: color_data = Z;
		19'b0111010110101010000: color_data = Z;
		19'b0111011000100101110: color_data = Z;
		19'b0111011000100101111: color_data = Z;
		19'b0111011000100110000: color_data = Z;
		19'b0111011000100110001: color_data = Z;
		19'b0111011000100111001: color_data = Z;
		19'b0111011000100111010: color_data = Z;
		19'b0111011000100111011: color_data = Z;
		19'b0111011000100111100: color_data = Z;
		19'b0111011000100111101: color_data = Z;
		19'b0111011000100111110: color_data = Z;
		19'b0111011000100111111: color_data = Z;
		19'b0111011000101000000: color_data = Z;
		19'b0111011000101000001: color_data = Z;
		19'b0111011000101000010: color_data = Z;
		19'b0111011000101000011: color_data = Z;
		19'b0111011000101000100: color_data = Z;
		19'b0111011000101000101: color_data = Z;
		19'b0111011000101000110: color_data = Z;
		19'b0111011000101000111: color_data = Z;
		19'b0111011000101001000: color_data = Z;
		19'b0111011000101001001: color_data = Z;
		19'b0111011000101001011: color_data = Z;
		19'b0111011000101001100: color_data = Z;
		19'b0111011000101001111: color_data = Z;
		19'b0111011000101010000: color_data = Z;
		19'b0111011010100101111: color_data = Z;
		19'b0111011010100110000: color_data = Z;
		19'b0111011010100110001: color_data = Z;
		19'b0111011010100110010: color_data = Z;
		19'b0111011010100111010: color_data = Z;
		19'b0111011010100111011: color_data = Z;
		19'b0111011010100111100: color_data = Z;
		19'b0111011010100111101: color_data = Z;
		19'b0111011010100111110: color_data = Z;
		19'b0111011010100111111: color_data = Z;
		19'b0111011010101000000: color_data = Z;
		19'b0111011010101000001: color_data = Z;
		19'b0111011010101000010: color_data = Z;
		19'b0111011010101000011: color_data = Z;
		19'b0111011010101000100: color_data = Z;
		19'b0111011010101000101: color_data = Z;
		19'b0111011010101000110: color_data = Z;
		19'b0111011010101000111: color_data = Z;
		19'b0111011010101001000: color_data = Z;
		19'b0111011010101001001: color_data = Z;
		19'b0111011010101001010: color_data = Z;
		19'b0111011010101001011: color_data = Z;
		19'b0111011010101001100: color_data = Z;
		19'b0111011010101001111: color_data = Z;
		19'b0111011100100101111: color_data = Z;
		19'b0111011100100110000: color_data = Z;
		19'b0111011100100110001: color_data = Z;
		19'b0111011100100110010: color_data = Z;
		19'b0111011100100110011: color_data = Z;
		19'b0111011100100110100: color_data = Z;
		19'b0111011100100111001: color_data = Z;
		19'b0111011100100111010: color_data = Z;
		19'b0111011100100111011: color_data = Z;
		19'b0111011100100111100: color_data = Z;
		19'b0111011100100111101: color_data = Z;
		19'b0111011100100111110: color_data = Z;
		19'b0111011100100111111: color_data = Z;
		19'b0111011100101000000: color_data = Z;
		19'b0111011100101000001: color_data = Z;
		19'b0111011100101000010: color_data = Z;
		19'b0111011100101000011: color_data = Z;
		19'b0111011100101000100: color_data = Z;
		19'b0111011100101000101: color_data = Z;
		19'b0111011100101000110: color_data = Z;
		19'b0111011100101000111: color_data = Z;
		19'b0111011100101001000: color_data = Z;
		19'b0111011100101001001: color_data = Z;
		19'b0111011100101001010: color_data = Z;
		19'b0111011100101001011: color_data = Z;
		19'b0111011100101001100: color_data = Z;
		19'b0111011100101001101: color_data = Z;
		19'b0111011100101001111: color_data = Z;
		19'b0111011110100101111: color_data = Z;
		19'b0111011110100110000: color_data = Z;
		19'b0111011110100110001: color_data = Z;
		19'b0111011110100110010: color_data = Z;
		19'b0111011110100110011: color_data = Z;
		19'b0111011110100110100: color_data = Z;
		19'b0111011110100110101: color_data = Z;
		19'b0111011110100110110: color_data = Z;
		19'b0111011110100110111: color_data = Z;
		19'b0111011110100111000: color_data = Z;
		19'b0111011110100111001: color_data = Z;
		19'b0111011110100111010: color_data = Z;
		19'b0111011110100111011: color_data = Z;
		19'b0111011110100111100: color_data = Z;
		19'b0111011110100111101: color_data = Z;
		19'b0111011110100111110: color_data = Z;
		19'b0111011110100111111: color_data = Z;
		19'b0111011110101000000: color_data = Z;
		19'b0111011110101000001: color_data = Z;
		19'b0111011110101000010: color_data = Z;
		19'b0111011110101000011: color_data = Z;
		19'b0111011110101000100: color_data = Z;
		19'b0111011110101000101: color_data = Z;
		19'b0111011110101000110: color_data = Z;
		19'b0111011110101000111: color_data = Z;
		19'b0111011110101001000: color_data = Z;
		19'b0111011110101001001: color_data = Z;
		19'b0111011110101001010: color_data = Z;
		19'b0111011110101001011: color_data = Z;
		19'b0111011110101001100: color_data = Z;
		19'b0111011110101001101: color_data = Z;
		19'b0111100000100101111: color_data = Z;
		19'b0111100000100110000: color_data = Z;
		19'b0111100000100110001: color_data = Z;
		19'b0111100000100110010: color_data = Z;
		19'b0111100000100110011: color_data = Z;
		19'b0111100000100110100: color_data = Z;
		19'b0111100000100110101: color_data = Z;
		19'b0111100000100110110: color_data = Z;
		19'b0111100000100110111: color_data = Z;
		19'b0111100000100111000: color_data = Z;
		19'b0111100000100111001: color_data = Z;
		19'b0111100000100111010: color_data = Z;
		19'b0111100000100111011: color_data = Z;
		19'b0111100000100111100: color_data = Z;
		19'b0111100000100111101: color_data = Z;
		19'b0111100000100111110: color_data = Z;
		19'b0111100000100111111: color_data = Z;
		19'b0111100000101000000: color_data = Z;
		19'b0111100000101000001: color_data = Z;
		19'b0111100000101000010: color_data = Z;
		19'b0111100000101000011: color_data = Z;
		19'b0111100000101000100: color_data = Z;
		19'b0111100000101000101: color_data = Z;
		19'b0111100000101000110: color_data = Z;
		19'b0111100000101000111: color_data = Z;
		19'b0111100000101001000: color_data = Z;
		19'b0111100000101001001: color_data = Z;
		19'b0111100000101001010: color_data = Z;
		19'b0111100000101001011: color_data = Z;
		19'b0111100000101001100: color_data = Z;
		19'b0111100000101001101: color_data = Z;
		19'b0111100010100101111: color_data = Z;
		19'b0111100010100110000: color_data = Z;
		19'b0111100010100110001: color_data = Z;
		19'b0111100010100110010: color_data = Z;
		19'b0111100010100110011: color_data = Z;
		19'b0111100010100110100: color_data = Z;
		19'b0111100010100110101: color_data = Z;
		19'b0111100010100110110: color_data = Z;
		19'b0111100010100110111: color_data = Z;
		19'b0111100010100111000: color_data = Z;
		19'b0111100010100111001: color_data = Z;
		19'b0111100010100111010: color_data = Z;
		19'b0111100010100111011: color_data = Z;
		19'b0111100010100111100: color_data = Z;
		19'b0111100010100111101: color_data = Z;
		19'b0111100010100111110: color_data = Z;
		19'b0111100010100111111: color_data = Z;
		19'b0111100010101000001: color_data = Z;
		19'b0111100010101000010: color_data = Z;
		19'b0111100010101000011: color_data = Z;
		19'b0111100010101000101: color_data = Z;
		19'b0111100010101000110: color_data = Z;
		19'b0111100010101000111: color_data = Z;
		19'b0111100010101001000: color_data = Z;
		19'b0111100010101001001: color_data = Z;
		19'b0111100010101001010: color_data = Z;
		19'b0111100010101001011: color_data = Z;
		19'b0111100010101001100: color_data = Z;
		19'b0111100010101001101: color_data = Z;
		19'b0111100010101001110: color_data = Z;
		19'b0111100100100110000: color_data = Z;
		19'b0111100100100110001: color_data = Z;
		19'b0111100100100110010: color_data = Z;
		19'b0111100100100110011: color_data = Z;
		19'b0111100100100110100: color_data = Z;
		19'b0111100100100110101: color_data = Z;
		19'b0111100100100110110: color_data = Z;
		19'b0111100100100110111: color_data = Z;
		19'b0111100100100111000: color_data = Z;
		19'b0111100100100111001: color_data = Z;
		19'b0111100100100111010: color_data = Z;
		19'b0111100100100111011: color_data = Z;
		19'b0111100100100111100: color_data = Z;
		19'b0111100100100111101: color_data = Z;
		19'b0111100100100111110: color_data = Z;
		19'b0111100100100111111: color_data = Z;
		19'b0111100100101000000: color_data = Z;
		19'b0111100100101000010: color_data = Z;
		19'b0111100100101000011: color_data = Z;
		19'b0111100100101000100: color_data = Z;
		19'b0111100100101000101: color_data = Z;
		19'b0111100100101000110: color_data = Z;
		19'b0111100100101000111: color_data = Z;
		19'b0111100100101001000: color_data = Z;
		19'b0111100100101001001: color_data = Z;
		19'b0111100100101001010: color_data = Z;
		19'b0111100100101001011: color_data = Z;
		19'b0111100100101001100: color_data = Z;
		19'b0111100100101001101: color_data = Z;
		19'b0111100100101001110: color_data = Z;
		19'b0111100110100110000: color_data = Z;
		19'b0111100110100110001: color_data = Z;
		19'b0111100110100110010: color_data = Z;
		19'b0111100110100110011: color_data = Z;
		19'b0111100110100110100: color_data = Z;
		19'b0111100110100110101: color_data = Z;
		19'b0111100110100110110: color_data = Z;
		19'b0111100110100110111: color_data = Z;
		19'b0111100110100111000: color_data = Z;
		19'b0111100110100111001: color_data = Z;
		19'b0111100110100111010: color_data = Z;
		19'b0111100110100111011: color_data = Z;
		19'b0111100110100111100: color_data = Z;
		19'b0111100110100111101: color_data = Z;
		19'b0111100110100111110: color_data = Z;
		19'b0111100110100111111: color_data = Z;
		19'b0111100110101000000: color_data = Z;
		19'b0111100110101000001: color_data = Z;
		19'b0111100110101000010: color_data = Z;
		19'b0111100110101000011: color_data = Z;
		19'b0111100110101000100: color_data = Z;
		19'b0111100110101000101: color_data = Z;
		19'b0111100110101000110: color_data = Z;
		19'b0111100110101000111: color_data = Z;
		19'b0111100110101001011: color_data = Z;
		19'b0111100110101001100: color_data = Z;
		19'b0111100110101001101: color_data = Z;
		19'b0111100110101001110: color_data = Z;
		19'b0111101000100110001: color_data = Z;
		19'b0111101000100110010: color_data = Z;
		19'b0111101000100110011: color_data = Z;
		19'b0111101000100110100: color_data = Z;
		19'b0111101000100110101: color_data = Z;
		19'b0111101000100110110: color_data = Z;
		19'b0111101000100110111: color_data = Z;
		19'b0111101000100111100: color_data = Z;
		19'b0111101000100111101: color_data = Z;
		19'b0111101000100111110: color_data = Z;
		19'b0111101000100111111: color_data = Z;
		19'b0111101000101000000: color_data = Z;
		19'b0111101000101000001: color_data = Z;
		19'b0111101000101000010: color_data = Z;
		19'b0111101000101000011: color_data = Z;
		19'b0111101000101000100: color_data = Z;
		19'b0111101000101000101: color_data = Z;
		19'b0111101000101001100: color_data = Z;
		19'b0111101000101001101: color_data = Z;
		19'b0111101000101001110: color_data = Z;
		19'b0111101010100110010: color_data = Z;
		19'b0111101010100110011: color_data = Z;
		19'b0111101010100110100: color_data = Z;
		19'b0111101010100110101: color_data = Z;
		19'b0111101010100110110: color_data = Z;
		19'b0111101010100111010: color_data = Z;
		19'b0111101010100111011: color_data = Z;
		19'b0111101010100111111: color_data = Z;
		19'b0111101010101000000: color_data = Z;
		19'b0111101010101000111: color_data = Z;
		19'b0111101010101001100: color_data = Z;
		19'b0111101010101001101: color_data = Z;
		19'b0111101010101001110: color_data = Z;
		19'b0111101100100110010: color_data = Z;
		19'b0111101100100110011: color_data = Z;
		19'b0111101100100110100: color_data = Z;
		19'b0111101100100110101: color_data = Z;
		19'b0111101100100110110: color_data = Z;
		19'b0111101100100111101: color_data = Z;
		19'b0111101100100111110: color_data = Z;
		19'b0111101100101000001: color_data = Z;
		19'b0111101100101000010: color_data = Z;
		19'b0111101100101000100: color_data = Z;
		19'b0111101100101000101: color_data = Z;
		19'b0111101100101001100: color_data = Z;
		19'b0111101100101001101: color_data = Z;
		19'b0111101110100110011: color_data = Z;
		19'b0111101110100110100: color_data = Z;
		19'b0111101110100110101: color_data = Z;
		19'b0111101110100110110: color_data = Z;
		19'b0111101110100111111: color_data = Z;
		19'b0111101110101000000: color_data = Z;
		19'b0111101110101001100: color_data = Z;
		19'b0111101110101001101: color_data = Z;
		19'b0111110000100110100: color_data = Z;
		19'b0111110000100110101: color_data = Z;
		19'b0111110000100110110: color_data = Z;
		19'b0111110000100110111: color_data = Z;
		19'b0111110000101001011: color_data = Z;
		19'b0111110000101001100: color_data = Z;
		19'b0111110000101001101: color_data = Z;
		19'b0111110010100110101: color_data = Z;
		19'b0111110010100110110: color_data = Z;
		19'b0111110010100110111: color_data = Z;
		19'b0111110010100111000: color_data = Z;
		19'b0111110010100111001: color_data = Z;
		19'b0111110010101000110: color_data = Z;
		19'b0111110010101001000: color_data = Z;
		19'b0111110010101001010: color_data = Z;
		19'b0111110010101001011: color_data = Z;
		19'b0111110010101001100: color_data = Z;
		19'b0111110100100110101: color_data = Z;
		19'b0111110100100110110: color_data = Z;
		19'b0111110100100110111: color_data = Z;
		19'b0111110100100111000: color_data = Z;
		19'b0111110100100111001: color_data = Z;
		19'b0111110100100111010: color_data = Z;
		19'b0111110100100111011: color_data = Z;
		19'b0111110100100111111: color_data = Z;
		19'b0111110100101000100: color_data = Z;
		19'b0111110100101000101: color_data = Z;
		19'b0111110100101001010: color_data = Z;
		19'b0111110100101001011: color_data = Z;
		19'b0111110110100110110: color_data = Z;
		19'b0111110110100110111: color_data = Z;
		19'b0111110110100111000: color_data = Z;
		19'b0111110110100111001: color_data = Z;
		19'b0111110110100111010: color_data = Z;
		19'b0111110110100111011: color_data = Z;
		19'b0111110110100111100: color_data = Z;
		19'b0111110110100111101: color_data = Z;
		19'b0111110110101000000: color_data = Z;
		19'b0111110110101000010: color_data = Z;
		19'b0111110110101000011: color_data = Z;
		19'b0111110110101001000: color_data = Z;
		19'b0111110110101001001: color_data = Z;
		19'b0111111000100111000: color_data = Z;
		19'b0111111000100111001: color_data = Z;
		19'b0111111000100111010: color_data = Z;
		19'b0111111000100111011: color_data = Z;
		19'b0111111000100111100: color_data = Z;
		19'b0111111000100111101: color_data = Z;
		19'b0111111000100111110: color_data = Z;
		19'b0111111000100111111: color_data = Z;
		19'b0111111000101000101: color_data = Z;
		19'b0111111000101000110: color_data = Z;
		19'b0111111000101000111: color_data = Z;
		19'b0111111000101001000: color_data = Z;
		19'b0111111010100111001: color_data = Z;
		19'b0111111010100111010: color_data = Z;
		19'b0111111010100111011: color_data = Z;
		19'b0111111010100111100: color_data = Z;
		19'b0111111010100111101: color_data = Z;
		19'b0111111010100111110: color_data = Z;
		19'b0111111010100111111: color_data = Z;
		19'b0111111010101000000: color_data = Z;
		19'b0111111010101000001: color_data = Z;
		19'b0111111010101000010: color_data = Z;
		19'b0111111010101000011: color_data = Z;
		19'b0111111010101000100: color_data = Z;
		19'b0111111010101000101: color_data = Z;
		19'b0111111010101000110: color_data = Z;
		19'b0111111010101000111: color_data = Z;
		19'b0111111100100111011: color_data = Z;
		19'b0111111100100111100: color_data = Z;
		19'b0111111100100111101: color_data = Z;
		19'b0111111100100111110: color_data = Z;
		19'b0111111100100111111: color_data = Z;
		19'b0111111100101000000: color_data = Z;
		19'b0111111100101000001: color_data = Z;
		19'b0111111100101000010: color_data = Z;
		19'b0111111100101000011: color_data = Z;
		19'b0111111100101000100: color_data = Z;
		19'b0111111100101000101: color_data = Z;
		19'b0111111100101000110: color_data = Z;
		19'b0111111110100111110: color_data = Z;
		19'b0111111110100111111: color_data = Z;
		19'b0111111110101000000: color_data = Z;
		19'b0111111110101000001: color_data = Z;
		19'b0111111110101000010: color_data = Z;
		19'b0111111110101000011: color_data = Z;
		19'b0111111110101000100: color_data = Z;
		19'b1000000000101000000: color_data = Z;
		19'b1000000000101000001: color_data = Z;
		19'b1000000000101000010: color_data = Z;
		19'b1000000000101000011: color_data = Z;
		19'b1000000010100111011: color_data = Z;
		19'b1000000010100111100: color_data = Z;
		19'b1000000010100111101: color_data = Z;
		19'b1000000010101000110: color_data = Z;
		19'b1000000100100111011: color_data = Z;
		19'b1000000100100111100: color_data = Z;
		19'b1000000100100111101: color_data = Z;
		19'b1000000100100111110: color_data = Z;
		19'b1000000100101000010: color_data = Z;
		19'b1000000100101000011: color_data = Z;
		19'b1000000100101000100: color_data = Z;
		19'b1000000100101000101: color_data = Z;
		19'b1000000100101000110: color_data = Z;
		19'b1000000110100111100: color_data = Z;
		19'b1000000110100111101: color_data = Z;
		19'b1000000110100111110: color_data = Z;
		19'b1000000110100111111: color_data = Z;
		19'b1000000110101000000: color_data = Z;
		19'b1000000110101000001: color_data = Z;
		19'b1000000110101000010: color_data = Z;
		19'b1000000110101000011: color_data = Z;
		19'b1000000110101000100: color_data = Z;
		19'b1000000110101000101: color_data = Z;
		19'b1000000110101000110: color_data = Z;
		19'b1000001000100111100: color_data = Z;
		19'b1000001000100111101: color_data = Z;
		19'b1000001000100111110: color_data = Z;
		19'b1000001000100111111: color_data = Z;
		19'b1000001000101000000: color_data = Z;
		19'b1000001000101000001: color_data = Z;
		19'b1000001000101000010: color_data = Z;
		19'b1000001000101000011: color_data = Z;
		19'b1000001000101000100: color_data = Z;
		19'b1000001000101000101: color_data = Z;
		19'b1000001000101000110: color_data = Z;
		19'b1000001010100111100: color_data = Z;
		19'b1000001010100111101: color_data = Z;
		19'b1000001010100111110: color_data = Z;
		19'b1000001010100111111: color_data = Z;
		19'b1000001010101000000: color_data = Z;
		19'b1000001010101000001: color_data = Z;
		19'b1000001010101000010: color_data = Z;
		19'b1000001010101000011: color_data = Z;
		19'b1000001010101000100: color_data = Z;
		19'b1000001010101000101: color_data = Z;
		19'b1000001010101000110: color_data = Z;
		19'b1000001100100111101: color_data = Z;
		19'b1000001100100111110: color_data = Z;
		19'b1000001100100111111: color_data = Z;
		19'b1000001100101000000: color_data = Z;
		19'b1000001100101000001: color_data = Z;
		19'b1000001100101000010: color_data = Z;
		19'b1000001100101000011: color_data = Z;
		19'b1000001100101000100: color_data = Z;
		19'b1000001100101000101: color_data = Z;
		19'b1000001100101000110: color_data = Z;
		19'b1000001110100111110: color_data = Z;
		19'b1000001110100111111: color_data = Z;
		19'b1000001110101000000: color_data = Z;
		19'b1000001110101000001: color_data = Z;
		19'b1000001110101000010: color_data = Z;
		19'b1000001110101000011: color_data = Z;
		19'b1000001110101000100: color_data = Z;
		19'b1000001110101000101: color_data = Z;
		19'b1000010000101000000: color_data = Z;
		19'b1000010000101000001: color_data = Z;
		19'b1000010000101000010: color_data = Z;
		19'b1000010000101000011: color_data = Z;
		19'b1000010000101000100: color_data = Z;
		default: color_data = 12'b000000000000;
	endcase
endmodule
