module death_3_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);
    parameter Z = 12'b111111111111; 
	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		19'b0000001000100110010: color_data = Z;
		19'b0000001000100110011: color_data = Z;
		19'b0000001000100110100: color_data = Z;
		19'b0000001000100110101: color_data = Z;
		19'b0000001000100110110: color_data = Z;
		19'b0000001000100110111: color_data = Z;
		19'b0000001000100111000: color_data = Z;
		19'b0000001000100111001: color_data = Z;
		19'b0000001000100111010: color_data = Z;
		19'b0000001000100111011: color_data = Z;
		19'b0000001000100111100: color_data = Z;
		19'b0000001000100111101: color_data = Z;
		19'b0000001000101010000: color_data = Z;
		19'b0000001000101010001: color_data = Z;
		19'b0000001000101010010: color_data = Z;
		19'b0000001000101010011: color_data = Z;
		19'b0000001000101010100: color_data = Z;
		19'b0000001000101010101: color_data = Z;
		19'b0000001000101010110: color_data = Z;
		19'b0000001010100101111: color_data = Z;
		19'b0000001010100110000: color_data = Z;
		19'b0000001010100110001: color_data = Z;
		19'b0000001010100110010: color_data = Z;
		19'b0000001010100110011: color_data = Z;
		19'b0000001010100110100: color_data = Z;
		19'b0000001010100110101: color_data = Z;
		19'b0000001010100110110: color_data = Z;
		19'b0000001010100110111: color_data = Z;
		19'b0000001010100111000: color_data = Z;
		19'b0000001010100111001: color_data = Z;
		19'b0000001010100111010: color_data = Z;
		19'b0000001010100111011: color_data = Z;
		19'b0000001010100111100: color_data = Z;
		19'b0000001010100111101: color_data = Z;
		19'b0000001010100111110: color_data = Z;
		19'b0000001010100111111: color_data = Z;
		19'b0000001010101000000: color_data = Z;
		19'b0000001010101000001: color_data = Z;
		19'b0000001010101000010: color_data = Z;
		19'b0000001010101000011: color_data = Z;
		19'b0000001010101000100: color_data = Z;
		19'b0000001010101000101: color_data = Z;
		19'b0000001010101000110: color_data = Z;
		19'b0000001010101000111: color_data = Z;
		19'b0000001010101001000: color_data = Z;
		19'b0000001010101001001: color_data = Z;
		19'b0000001010101001010: color_data = Z;
		19'b0000001010101001011: color_data = Z;
		19'b0000001010101001100: color_data = Z;
		19'b0000001010101001101: color_data = Z;
		19'b0000001010101001110: color_data = Z;
		19'b0000001010101001111: color_data = Z;
		19'b0000001010101010000: color_data = Z;
		19'b0000001010101010001: color_data = Z;
		19'b0000001010101010010: color_data = Z;
		19'b0000001010101010011: color_data = Z;
		19'b0000001010101010100: color_data = Z;
		19'b0000001010101010101: color_data = Z;
		19'b0000001010101010110: color_data = Z;
		19'b0000001010101010111: color_data = Z;
		19'b0000001010101011000: color_data = Z;
		19'b0000001010101011001: color_data = Z;
		19'b0000001010101011010: color_data = Z;
		19'b0000001100100101100: color_data = Z;
		19'b0000001100100101101: color_data = Z;
		19'b0000001100100101110: color_data = Z;
		19'b0000001100100101111: color_data = Z;
		19'b0000001100100110000: color_data = Z;
		19'b0000001100100110001: color_data = Z;
		19'b0000001100100110010: color_data = Z;
		19'b0000001100100110011: color_data = Z;
		19'b0000001100100110100: color_data = Z;
		19'b0000001100100110101: color_data = Z;
		19'b0000001100100110110: color_data = Z;
		19'b0000001100100110111: color_data = Z;
		19'b0000001100100111000: color_data = Z;
		19'b0000001100100111001: color_data = Z;
		19'b0000001100100111010: color_data = Z;
		19'b0000001100100111011: color_data = Z;
		19'b0000001100100111100: color_data = Z;
		19'b0000001100100111101: color_data = Z;
		19'b0000001100100111110: color_data = Z;
		19'b0000001100100111111: color_data = Z;
		19'b0000001100101000000: color_data = Z;
		19'b0000001100101000001: color_data = Z;
		19'b0000001100101000010: color_data = Z;
		19'b0000001100101000011: color_data = Z;
		19'b0000001100101000100: color_data = Z;
		19'b0000001100101000101: color_data = Z;
		19'b0000001100101000110: color_data = Z;
		19'b0000001100101000111: color_data = Z;
		19'b0000001100101001000: color_data = Z;
		19'b0000001100101001001: color_data = Z;
		19'b0000001100101001010: color_data = Z;
		19'b0000001100101001011: color_data = Z;
		19'b0000001100101001100: color_data = Z;
		19'b0000001100101001101: color_data = Z;
		19'b0000001100101001110: color_data = Z;
		19'b0000001100101001111: color_data = Z;
		19'b0000001100101010000: color_data = Z;
		19'b0000001100101010001: color_data = Z;
		19'b0000001100101010010: color_data = Z;
		19'b0000001100101010011: color_data = Z;
		19'b0000001100101010100: color_data = Z;
		19'b0000001100101010101: color_data = Z;
		19'b0000001100101010110: color_data = Z;
		19'b0000001100101010111: color_data = Z;
		19'b0000001100101011000: color_data = Z;
		19'b0000001100101011001: color_data = Z;
		19'b0000001100101011010: color_data = Z;
		19'b0000001100101011011: color_data = Z;
		19'b0000001100101011100: color_data = Z;
		19'b0000001100101011101: color_data = Z;
		19'b0000001110100101001: color_data = Z;
		19'b0000001110100101010: color_data = Z;
		19'b0000001110100101011: color_data = Z;
		19'b0000001110100101100: color_data = Z;
		19'b0000001110100101101: color_data = Z;
		19'b0000001110100101110: color_data = Z;
		19'b0000001110100101111: color_data = Z;
		19'b0000001110100110000: color_data = Z;
		19'b0000001110100110001: color_data = Z;
		19'b0000001110100110010: color_data = Z;
		19'b0000001110100110011: color_data = Z;
		19'b0000001110100110100: color_data = Z;
		19'b0000001110100110101: color_data = Z;
		19'b0000001110100110110: color_data = Z;
		19'b0000001110100110111: color_data = Z;
		19'b0000001110100111000: color_data = Z;
		19'b0000001110100111001: color_data = Z;
		19'b0000001110100111010: color_data = Z;
		19'b0000001110100111011: color_data = Z;
		19'b0000001110100111100: color_data = Z;
		19'b0000001110100111101: color_data = Z;
		19'b0000001110100111110: color_data = Z;
		19'b0000001110100111111: color_data = Z;
		19'b0000001110101000000: color_data = Z;
		19'b0000001110101000001: color_data = Z;
		19'b0000001110101000010: color_data = Z;
		19'b0000001110101000011: color_data = Z;
		19'b0000001110101000100: color_data = Z;
		19'b0000001110101000101: color_data = Z;
		19'b0000001110101000110: color_data = Z;
		19'b0000001110101000111: color_data = Z;
		19'b0000001110101001000: color_data = Z;
		19'b0000001110101001001: color_data = Z;
		19'b0000001110101001010: color_data = Z;
		19'b0000001110101001011: color_data = Z;
		19'b0000001110101001100: color_data = Z;
		19'b0000001110101001101: color_data = Z;
		19'b0000001110101001110: color_data = Z;
		19'b0000001110101001111: color_data = Z;
		19'b0000001110101010000: color_data = Z;
		19'b0000001110101010001: color_data = Z;
		19'b0000001110101010010: color_data = Z;
		19'b0000001110101010011: color_data = Z;
		19'b0000001110101010100: color_data = Z;
		19'b0000001110101010101: color_data = Z;
		19'b0000001110101010110: color_data = Z;
		19'b0000001110101010111: color_data = Z;
		19'b0000001110101011000: color_data = Z;
		19'b0000001110101011001: color_data = Z;
		19'b0000001110101011010: color_data = Z;
		19'b0000001110101011011: color_data = Z;
		19'b0000001110101011100: color_data = Z;
		19'b0000001110101011101: color_data = Z;
		19'b0000001110101011110: color_data = Z;
		19'b0000001110101011111: color_data = Z;
		19'b0000001110101100000: color_data = Z;
		19'b0000010000100100100: color_data = Z;
		19'b0000010000100100101: color_data = Z;
		19'b0000010000100100110: color_data = Z;
		19'b0000010000100100111: color_data = Z;
		19'b0000010000100101000: color_data = Z;
		19'b0000010000100101001: color_data = Z;
		19'b0000010000100101010: color_data = Z;
		19'b0000010000100101011: color_data = Z;
		19'b0000010000100101100: color_data = Z;
		19'b0000010000100101101: color_data = Z;
		19'b0000010000100101110: color_data = Z;
		19'b0000010000100101111: color_data = Z;
		19'b0000010000100110000: color_data = Z;
		19'b0000010000100111100: color_data = Z;
		19'b0000010000100111101: color_data = Z;
		19'b0000010000100111110: color_data = Z;
		19'b0000010000100111111: color_data = Z;
		19'b0000010000101000000: color_data = Z;
		19'b0000010000101000001: color_data = Z;
		19'b0000010000101000010: color_data = Z;
		19'b0000010000101000011: color_data = Z;
		19'b0000010000101000100: color_data = Z;
		19'b0000010000101000101: color_data = Z;
		19'b0000010000101000110: color_data = Z;
		19'b0000010000101000111: color_data = Z;
		19'b0000010000101001000: color_data = Z;
		19'b0000010000101001001: color_data = Z;
		19'b0000010000101001010: color_data = Z;
		19'b0000010000101001011: color_data = Z;
		19'b0000010000101001100: color_data = Z;
		19'b0000010000101001101: color_data = Z;
		19'b0000010000101001110: color_data = Z;
		19'b0000010000101001111: color_data = Z;
		19'b0000010000101010000: color_data = Z;
		19'b0000010000101010001: color_data = Z;
		19'b0000010000101010010: color_data = Z;
		19'b0000010000101010011: color_data = Z;
		19'b0000010000101010100: color_data = Z;
		19'b0000010000101010101: color_data = Z;
		19'b0000010000101010110: color_data = Z;
		19'b0000010000101010111: color_data = Z;
		19'b0000010000101011000: color_data = Z;
		19'b0000010000101011001: color_data = Z;
		19'b0000010000101011010: color_data = Z;
		19'b0000010000101011011: color_data = Z;
		19'b0000010000101011100: color_data = Z;
		19'b0000010000101011101: color_data = Z;
		19'b0000010000101011110: color_data = Z;
		19'b0000010000101011111: color_data = Z;
		19'b0000010000101100000: color_data = Z;
		19'b0000010000101100001: color_data = Z;
		19'b0000010000101100010: color_data = Z;
		19'b0000010000101100011: color_data = Z;
		19'b0000010010100100010: color_data = Z;
		19'b0000010010100100011: color_data = Z;
		19'b0000010010100100100: color_data = Z;
		19'b0000010010100100101: color_data = Z;
		19'b0000010010100100110: color_data = Z;
		19'b0000010010100100111: color_data = Z;
		19'b0000010010100101000: color_data = Z;
		19'b0000010010100101001: color_data = Z;
		19'b0000010010100101010: color_data = Z;
		19'b0000010010100101011: color_data = Z;
		19'b0000010010100111010: color_data = Z;
		19'b0000010010100111011: color_data = Z;
		19'b0000010010100111100: color_data = Z;
		19'b0000010010100111101: color_data = Z;
		19'b0000010010100111110: color_data = Z;
		19'b0000010010100111111: color_data = Z;
		19'b0000010010101000000: color_data = Z;
		19'b0000010010101000001: color_data = Z;
		19'b0000010010101000010: color_data = Z;
		19'b0000010010101000011: color_data = Z;
		19'b0000010010101000100: color_data = Z;
		19'b0000010010101000101: color_data = Z;
		19'b0000010010101000110: color_data = Z;
		19'b0000010010101000111: color_data = Z;
		19'b0000010010101001000: color_data = Z;
		19'b0000010010101001001: color_data = Z;
		19'b0000010010101001010: color_data = Z;
		19'b0000010010101001011: color_data = Z;
		19'b0000010010101001100: color_data = Z;
		19'b0000010010101001101: color_data = Z;
		19'b0000010010101001110: color_data = Z;
		19'b0000010010101001111: color_data = Z;
		19'b0000010010101010000: color_data = Z;
		19'b0000010010101010001: color_data = Z;
		19'b0000010010101010010: color_data = Z;
		19'b0000010010101010011: color_data = Z;
		19'b0000010010101010100: color_data = Z;
		19'b0000010010101010101: color_data = Z;
		19'b0000010010101010110: color_data = Z;
		19'b0000010010101010111: color_data = Z;
		19'b0000010010101011000: color_data = Z;
		19'b0000010010101011001: color_data = Z;
		19'b0000010010101011010: color_data = Z;
		19'b0000010010101011011: color_data = Z;
		19'b0000010010101011100: color_data = Z;
		19'b0000010010101011101: color_data = Z;
		19'b0000010010101011110: color_data = Z;
		19'b0000010010101011111: color_data = Z;
		19'b0000010010101100000: color_data = Z;
		19'b0000010010101100001: color_data = Z;
		19'b0000010010101100010: color_data = Z;
		19'b0000010010101100011: color_data = Z;
		19'b0000010010101100100: color_data = Z;
		19'b0000010010101100101: color_data = Z;
		19'b0000010010101100110: color_data = Z;
		19'b0000010100100110111: color_data = Z;
		19'b0000010100100111000: color_data = Z;
		19'b0000010100100111001: color_data = Z;
		19'b0000010100100111010: color_data = Z;
		19'b0000010100100111011: color_data = Z;
		19'b0000010100100111100: color_data = Z;
		19'b0000010100100111101: color_data = Z;
		19'b0000010100100111110: color_data = Z;
		19'b0000010100100111111: color_data = Z;
		19'b0000010100101000000: color_data = Z;
		19'b0000010100101000001: color_data = Z;
		19'b0000010100101000010: color_data = Z;
		19'b0000010100101000011: color_data = Z;
		19'b0000010100101000100: color_data = Z;
		19'b0000010100101000101: color_data = Z;
		19'b0000010100101000110: color_data = Z;
		19'b0000010100101000111: color_data = Z;
		19'b0000010100101001000: color_data = Z;
		19'b0000010100101001001: color_data = Z;
		19'b0000010100101001010: color_data = Z;
		19'b0000010100101001011: color_data = Z;
		19'b0000010100101001100: color_data = Z;
		19'b0000010100101001101: color_data = Z;
		19'b0000010100101001110: color_data = Z;
		19'b0000010100101001111: color_data = Z;
		19'b0000010100101010000: color_data = Z;
		19'b0000010100101010001: color_data = Z;
		19'b0000010100101010010: color_data = Z;
		19'b0000010100101010011: color_data = Z;
		19'b0000010100101010100: color_data = Z;
		19'b0000010100101010101: color_data = Z;
		19'b0000010100101010110: color_data = Z;
		19'b0000010100101010111: color_data = Z;
		19'b0000010100101011000: color_data = Z;
		19'b0000010100101011001: color_data = Z;
		19'b0000010100101011010: color_data = Z;
		19'b0000010100101011011: color_data = Z;
		19'b0000010100101011100: color_data = Z;
		19'b0000010100101011101: color_data = Z;
		19'b0000010100101011110: color_data = Z;
		19'b0000010100101011111: color_data = Z;
		19'b0000010100101100000: color_data = Z;
		19'b0000010100101100001: color_data = Z;
		19'b0000010100101100010: color_data = Z;
		19'b0000010100101100011: color_data = Z;
		19'b0000010100101100100: color_data = Z;
		19'b0000010100101100101: color_data = Z;
		19'b0000010100101100110: color_data = Z;
		19'b0000010100101100111: color_data = Z;
		19'b0000010100101101000: color_data = Z;
		19'b0000010100101101001: color_data = Z;
		19'b0000010110100110010: color_data = Z;
		19'b0000010110100110011: color_data = Z;
		19'b0000010110100110100: color_data = Z;
		19'b0000010110100110101: color_data = Z;
		19'b0000010110100110110: color_data = Z;
		19'b0000010110100110111: color_data = Z;
		19'b0000010110100111000: color_data = Z;
		19'b0000010110100111001: color_data = Z;
		19'b0000010110100111010: color_data = Z;
		19'b0000010110100111011: color_data = Z;
		19'b0000010110100111100: color_data = Z;
		19'b0000010110100111101: color_data = Z;
		19'b0000010110100111110: color_data = Z;
		19'b0000010110100111111: color_data = Z;
		19'b0000010110101000000: color_data = Z;
		19'b0000010110101000001: color_data = Z;
		19'b0000010110101000010: color_data = Z;
		19'b0000010110101000011: color_data = Z;
		19'b0000010110101000100: color_data = Z;
		19'b0000010110101000101: color_data = Z;
		19'b0000010110101000110: color_data = Z;
		19'b0000010110101000111: color_data = Z;
		19'b0000010110101001000: color_data = Z;
		19'b0000010110101001001: color_data = Z;
		19'b0000010110101001010: color_data = Z;
		19'b0000010110101001011: color_data = Z;
		19'b0000010110101001100: color_data = Z;
		19'b0000010110101001101: color_data = Z;
		19'b0000010110101001110: color_data = Z;
		19'b0000010110101001111: color_data = Z;
		19'b0000010110101010000: color_data = Z;
		19'b0000010110101010001: color_data = Z;
		19'b0000010110101010010: color_data = Z;
		19'b0000010110101010011: color_data = Z;
		19'b0000010110101010100: color_data = Z;
		19'b0000010110101010101: color_data = Z;
		19'b0000010110101010110: color_data = Z;
		19'b0000010110101010111: color_data = Z;
		19'b0000010110101011000: color_data = Z;
		19'b0000010110101011001: color_data = Z;
		19'b0000010110101011010: color_data = Z;
		19'b0000010110101011011: color_data = Z;
		19'b0000010110101011100: color_data = Z;
		19'b0000010110101011101: color_data = Z;
		19'b0000010110101011110: color_data = Z;
		19'b0000010110101011111: color_data = Z;
		19'b0000010110101100000: color_data = Z;
		19'b0000010110101100001: color_data = Z;
		19'b0000010110101100010: color_data = Z;
		19'b0000010110101100011: color_data = Z;
		19'b0000010110101100100: color_data = Z;
		19'b0000010110101100101: color_data = Z;
		19'b0000010110101100110: color_data = Z;
		19'b0000010110101100111: color_data = Z;
		19'b0000010110101101000: color_data = Z;
		19'b0000010110101101001: color_data = Z;
		19'b0000010110101101010: color_data = Z;
		19'b0000010110101101011: color_data = Z;
		19'b0000010110101101100: color_data = Z;
		19'b0000011000100011101: color_data = Z;
		19'b0000011000100101101: color_data = Z;
		19'b0000011000100101110: color_data = Z;
		19'b0000011000100101111: color_data = Z;
		19'b0000011000100110000: color_data = Z;
		19'b0000011000100110001: color_data = Z;
		19'b0000011000100110010: color_data = Z;
		19'b0000011000100110011: color_data = Z;
		19'b0000011000100110100: color_data = Z;
		19'b0000011000100110101: color_data = Z;
		19'b0000011000100110110: color_data = Z;
		19'b0000011000100110111: color_data = Z;
		19'b0000011000100111000: color_data = Z;
		19'b0000011000100111001: color_data = Z;
		19'b0000011000100111010: color_data = Z;
		19'b0000011000100111011: color_data = Z;
		19'b0000011000100111100: color_data = Z;
		19'b0000011000100111101: color_data = Z;
		19'b0000011000100111110: color_data = Z;
		19'b0000011000100111111: color_data = Z;
		19'b0000011000101000000: color_data = Z;
		19'b0000011000101000001: color_data = Z;
		19'b0000011000101000010: color_data = Z;
		19'b0000011000101000011: color_data = Z;
		19'b0000011000101000100: color_data = Z;
		19'b0000011000101000101: color_data = Z;
		19'b0000011000101000110: color_data = Z;
		19'b0000011000101000111: color_data = Z;
		19'b0000011000101001000: color_data = Z;
		19'b0000011000101001001: color_data = Z;
		19'b0000011000101001010: color_data = Z;
		19'b0000011000101001011: color_data = Z;
		19'b0000011000101001100: color_data = Z;
		19'b0000011000101001101: color_data = Z;
		19'b0000011000101001110: color_data = Z;
		19'b0000011000101001111: color_data = Z;
		19'b0000011000101010000: color_data = Z;
		19'b0000011000101010001: color_data = Z;
		19'b0000011000101010010: color_data = Z;
		19'b0000011000101010011: color_data = Z;
		19'b0000011000101010100: color_data = Z;
		19'b0000011000101010101: color_data = Z;
		19'b0000011000101010110: color_data = Z;
		19'b0000011000101010111: color_data = Z;
		19'b0000011000101011000: color_data = Z;
		19'b0000011000101011001: color_data = Z;
		19'b0000011000101011010: color_data = Z;
		19'b0000011000101011011: color_data = Z;
		19'b0000011000101011100: color_data = Z;
		19'b0000011000101011101: color_data = Z;
		19'b0000011000101011110: color_data = Z;
		19'b0000011000101011111: color_data = Z;
		19'b0000011000101100000: color_data = Z;
		19'b0000011000101100001: color_data = Z;
		19'b0000011000101100010: color_data = Z;
		19'b0000011000101100011: color_data = Z;
		19'b0000011000101100100: color_data = Z;
		19'b0000011000101100101: color_data = Z;
		19'b0000011000101100110: color_data = Z;
		19'b0000011000101100111: color_data = Z;
		19'b0000011000101101000: color_data = Z;
		19'b0000011000101101001: color_data = Z;
		19'b0000011000101101010: color_data = Z;
		19'b0000011000101101011: color_data = Z;
		19'b0000011000101101100: color_data = Z;
		19'b0000011000101101101: color_data = Z;
		19'b0000011000101101110: color_data = Z;
		19'b0000011000101101111: color_data = Z;
		19'b0000011010100011100: color_data = Z;
		19'b0000011010100011101: color_data = Z;
		19'b0000011010100011110: color_data = Z;
		19'b0000011010100011111: color_data = Z;
		19'b0000011010100100000: color_data = Z;
		19'b0000011010100100001: color_data = Z;
		19'b0000011010100100010: color_data = Z;
		19'b0000011010100100011: color_data = Z;
		19'b0000011010100100100: color_data = Z;
		19'b0000011010100100101: color_data = Z;
		19'b0000011010100100110: color_data = Z;
		19'b0000011010100100111: color_data = Z;
		19'b0000011010100101000: color_data = Z;
		19'b0000011010100101001: color_data = Z;
		19'b0000011010100101010: color_data = Z;
		19'b0000011010100101011: color_data = Z;
		19'b0000011010100101100: color_data = Z;
		19'b0000011010100101101: color_data = Z;
		19'b0000011010100101110: color_data = Z;
		19'b0000011010100101111: color_data = Z;
		19'b0000011010100110000: color_data = Z;
		19'b0000011010100110001: color_data = Z;
		19'b0000011010100110010: color_data = Z;
		19'b0000011010100110011: color_data = Z;
		19'b0000011010100110100: color_data = Z;
		19'b0000011010100110101: color_data = Z;
		19'b0000011010100110110: color_data = Z;
		19'b0000011010100110111: color_data = Z;
		19'b0000011010100111000: color_data = Z;
		19'b0000011010100111001: color_data = Z;
		19'b0000011010100111010: color_data = Z;
		19'b0000011010100111011: color_data = Z;
		19'b0000011010100111100: color_data = Z;
		19'b0000011010100111101: color_data = Z;
		19'b0000011010100111110: color_data = Z;
		19'b0000011010100111111: color_data = Z;
		19'b0000011010101000000: color_data = Z;
		19'b0000011010101000001: color_data = Z;
		19'b0000011010101000010: color_data = Z;
		19'b0000011010101000011: color_data = Z;
		19'b0000011010101000100: color_data = Z;
		19'b0000011010101000101: color_data = Z;
		19'b0000011010101000110: color_data = Z;
		19'b0000011010101000111: color_data = Z;
		19'b0000011010101001000: color_data = Z;
		19'b0000011010101001001: color_data = Z;
		19'b0000011010101001010: color_data = Z;
		19'b0000011010101001011: color_data = Z;
		19'b0000011010101001100: color_data = Z;
		19'b0000011010101001101: color_data = Z;
		19'b0000011010101001110: color_data = Z;
		19'b0000011010101001111: color_data = Z;
		19'b0000011010101010000: color_data = Z;
		19'b0000011010101010001: color_data = Z;
		19'b0000011010101010010: color_data = Z;
		19'b0000011010101010011: color_data = Z;
		19'b0000011010101010100: color_data = Z;
		19'b0000011010101010101: color_data = Z;
		19'b0000011010101010110: color_data = Z;
		19'b0000011010101010111: color_data = Z;
		19'b0000011010101011000: color_data = Z;
		19'b0000011010101011001: color_data = Z;
		19'b0000011010101011010: color_data = Z;
		19'b0000011010101011011: color_data = Z;
		19'b0000011010101011100: color_data = Z;
		19'b0000011010101011101: color_data = Z;
		19'b0000011010101011110: color_data = Z;
		19'b0000011010101011111: color_data = Z;
		19'b0000011010101100000: color_data = Z;
		19'b0000011010101100001: color_data = Z;
		19'b0000011010101100010: color_data = Z;
		19'b0000011010101100011: color_data = Z;
		19'b0000011010101100100: color_data = Z;
		19'b0000011010101100101: color_data = Z;
		19'b0000011010101100110: color_data = Z;
		19'b0000011010101100111: color_data = Z;
		19'b0000011010101101000: color_data = Z;
		19'b0000011010101101001: color_data = Z;
		19'b0000011010101101010: color_data = Z;
		19'b0000011010101101011: color_data = Z;
		19'b0000011010101101100: color_data = Z;
		19'b0000011010101101101: color_data = Z;
		19'b0000011010101101110: color_data = Z;
		19'b0000011010101101111: color_data = Z;
		19'b0000011010101110000: color_data = Z;
		19'b0000011010101110001: color_data = Z;
		19'b0000011010101110010: color_data = Z;
		19'b0000011100100011011: color_data = Z;
		19'b0000011100100011100: color_data = Z;
		19'b0000011100100011101: color_data = Z;
		19'b0000011100100011110: color_data = Z;
		19'b0000011100100011111: color_data = Z;
		19'b0000011100100100000: color_data = Z;
		19'b0000011100100100001: color_data = Z;
		19'b0000011100100100010: color_data = Z;
		19'b0000011100100100011: color_data = Z;
		19'b0000011100100100100: color_data = Z;
		19'b0000011100100100101: color_data = Z;
		19'b0000011100100100110: color_data = Z;
		19'b0000011100100100111: color_data = Z;
		19'b0000011100100101000: color_data = Z;
		19'b0000011100100101001: color_data = Z;
		19'b0000011100100101010: color_data = Z;
		19'b0000011100100101011: color_data = Z;
		19'b0000011100100101100: color_data = Z;
		19'b0000011100100101101: color_data = Z;
		19'b0000011100100101110: color_data = Z;
		19'b0000011100100101111: color_data = Z;
		19'b0000011100100110000: color_data = Z;
		19'b0000011100100110001: color_data = Z;
		19'b0000011100100110010: color_data = Z;
		19'b0000011100100110011: color_data = Z;
		19'b0000011100100110100: color_data = Z;
		19'b0000011100100110101: color_data = Z;
		19'b0000011100100110110: color_data = Z;
		19'b0000011100100110111: color_data = Z;
		19'b0000011100100111000: color_data = Z;
		19'b0000011100100111001: color_data = Z;
		19'b0000011100100111010: color_data = Z;
		19'b0000011100100111011: color_data = Z;
		19'b0000011100100111100: color_data = Z;
		19'b0000011100100111101: color_data = Z;
		19'b0000011100100111110: color_data = Z;
		19'b0000011100100111111: color_data = Z;
		19'b0000011100101000000: color_data = Z;
		19'b0000011100101000001: color_data = Z;
		19'b0000011100101000010: color_data = Z;
		19'b0000011100101000011: color_data = Z;
		19'b0000011100101000100: color_data = Z;
		19'b0000011100101000101: color_data = Z;
		19'b0000011100101000110: color_data = Z;
		19'b0000011100101000111: color_data = Z;
		19'b0000011100101001000: color_data = Z;
		19'b0000011100101001001: color_data = Z;
		19'b0000011100101001010: color_data = Z;
		19'b0000011100101001011: color_data = Z;
		19'b0000011100101001100: color_data = Z;
		19'b0000011100101001101: color_data = Z;
		19'b0000011100101001110: color_data = Z;
		19'b0000011100101001111: color_data = Z;
		19'b0000011100101010000: color_data = Z;
		19'b0000011100101010001: color_data = Z;
		19'b0000011100101010010: color_data = Z;
		19'b0000011100101010011: color_data = Z;
		19'b0000011100101010100: color_data = Z;
		19'b0000011100101010101: color_data = Z;
		19'b0000011100101010110: color_data = Z;
		19'b0000011100101010111: color_data = Z;
		19'b0000011100101011000: color_data = Z;
		19'b0000011100101011001: color_data = Z;
		19'b0000011100101011010: color_data = Z;
		19'b0000011100101011011: color_data = Z;
		19'b0000011100101011100: color_data = Z;
		19'b0000011100101011101: color_data = Z;
		19'b0000011100101011110: color_data = Z;
		19'b0000011100101011111: color_data = Z;
		19'b0000011100101100000: color_data = Z;
		19'b0000011100101100001: color_data = Z;
		19'b0000011100101100010: color_data = Z;
		19'b0000011100101100011: color_data = Z;
		19'b0000011100101100100: color_data = Z;
		19'b0000011100101100101: color_data = Z;
		19'b0000011100101100110: color_data = Z;
		19'b0000011100101100111: color_data = Z;
		19'b0000011100101101000: color_data = Z;
		19'b0000011100101101001: color_data = Z;
		19'b0000011100101101010: color_data = Z;
		19'b0000011100101101011: color_data = Z;
		19'b0000011100101101100: color_data = Z;
		19'b0000011100101101101: color_data = Z;
		19'b0000011100101101110: color_data = Z;
		19'b0000011100101101111: color_data = Z;
		19'b0000011100101110000: color_data = Z;
		19'b0000011100101110001: color_data = Z;
		19'b0000011100101110010: color_data = Z;
		19'b0000011100101110011: color_data = Z;
		19'b0000011100101110100: color_data = Z;
		19'b0000011100101110101: color_data = Z;
		19'b0000011100101110110: color_data = Z;
		19'b0000011110100011010: color_data = Z;
		19'b0000011110100011011: color_data = Z;
		19'b0000011110100011100: color_data = Z;
		19'b0000011110100011101: color_data = Z;
		19'b0000011110100011110: color_data = Z;
		19'b0000011110100011111: color_data = Z;
		19'b0000011110100100000: color_data = Z;
		19'b0000011110100100001: color_data = Z;
		19'b0000011110100100010: color_data = Z;
		19'b0000011110100100011: color_data = Z;
		19'b0000011110100100100: color_data = Z;
		19'b0000011110100100101: color_data = Z;
		19'b0000011110100100110: color_data = Z;
		19'b0000011110100100111: color_data = Z;
		19'b0000011110100101000: color_data = Z;
		19'b0000011110100101001: color_data = Z;
		19'b0000011110100101010: color_data = Z;
		19'b0000011110100101011: color_data = Z;
		19'b0000011110100101100: color_data = Z;
		19'b0000011110100101101: color_data = Z;
		19'b0000011110100101110: color_data = Z;
		19'b0000011110100101111: color_data = Z;
		19'b0000011110100110000: color_data = Z;
		19'b0000011110100110001: color_data = Z;
		19'b0000011110100110010: color_data = Z;
		19'b0000011110100110011: color_data = Z;
		19'b0000011110100110100: color_data = Z;
		19'b0000011110100110101: color_data = Z;
		19'b0000011110100110110: color_data = Z;
		19'b0000011110100110111: color_data = Z;
		19'b0000011110100111000: color_data = Z;
		19'b0000011110100111001: color_data = Z;
		19'b0000011110100111010: color_data = Z;
		19'b0000011110100111011: color_data = Z;
		19'b0000011110100111100: color_data = Z;
		19'b0000011110100111101: color_data = Z;
		19'b0000011110100111110: color_data = Z;
		19'b0000011110100111111: color_data = Z;
		19'b0000011110101000000: color_data = Z;
		19'b0000011110101000001: color_data = Z;
		19'b0000011110101000010: color_data = Z;
		19'b0000011110101000011: color_data = Z;
		19'b0000011110101000100: color_data = Z;
		19'b0000011110101000101: color_data = Z;
		19'b0000011110101000110: color_data = Z;
		19'b0000011110101000111: color_data = Z;
		19'b0000011110101001000: color_data = Z;
		19'b0000011110101001001: color_data = Z;
		19'b0000011110101001010: color_data = Z;
		19'b0000011110101001011: color_data = Z;
		19'b0000011110101001100: color_data = Z;
		19'b0000011110101001101: color_data = Z;
		19'b0000011110101001110: color_data = Z;
		19'b0000011110101001111: color_data = Z;
		19'b0000011110101010000: color_data = Z;
		19'b0000011110101010001: color_data = Z;
		19'b0000011110101010010: color_data = Z;
		19'b0000011110101010011: color_data = Z;
		19'b0000011110101010100: color_data = Z;
		19'b0000011110101010101: color_data = Z;
		19'b0000011110101010110: color_data = Z;
		19'b0000011110101010111: color_data = Z;
		19'b0000011110101011000: color_data = Z;
		19'b0000011110101011001: color_data = Z;
		19'b0000011110101011010: color_data = Z;
		19'b0000011110101011011: color_data = Z;
		19'b0000011110101011100: color_data = Z;
		19'b0000011110101011101: color_data = Z;
		19'b0000011110101011110: color_data = Z;
		19'b0000011110101011111: color_data = Z;
		19'b0000011110101100000: color_data = Z;
		19'b0000011110101100001: color_data = Z;
		19'b0000011110101100010: color_data = Z;
		19'b0000011110101100011: color_data = Z;
		19'b0000011110101100100: color_data = Z;
		19'b0000011110101100101: color_data = Z;
		19'b0000011110101100110: color_data = Z;
		19'b0000011110101100111: color_data = Z;
		19'b0000011110101101000: color_data = Z;
		19'b0000011110101101001: color_data = Z;
		19'b0000011110101101010: color_data = Z;
		19'b0000011110101101011: color_data = Z;
		19'b0000011110101101100: color_data = Z;
		19'b0000011110101101101: color_data = Z;
		19'b0000011110101101110: color_data = Z;
		19'b0000011110101101111: color_data = Z;
		19'b0000011110101110000: color_data = Z;
		19'b0000011110101110001: color_data = Z;
		19'b0000011110101110010: color_data = Z;
		19'b0000011110101110011: color_data = Z;
		19'b0000011110101110100: color_data = Z;
		19'b0000011110101110101: color_data = Z;
		19'b0000011110101110110: color_data = Z;
		19'b0000011110101110111: color_data = Z;
		19'b0000011110101111000: color_data = Z;
		19'b0000011110101111001: color_data = Z;
		19'b0000100000100010111: color_data = Z;
		19'b0000100000100011000: color_data = Z;
		19'b0000100000100011001: color_data = Z;
		19'b0000100000100011010: color_data = Z;
		19'b0000100000100011011: color_data = Z;
		19'b0000100000100011100: color_data = Z;
		19'b0000100000100011101: color_data = Z;
		19'b0000100000100011110: color_data = Z;
		19'b0000100000100011111: color_data = Z;
		19'b0000100000100100000: color_data = Z;
		19'b0000100000100100001: color_data = Z;
		19'b0000100000100100010: color_data = Z;
		19'b0000100000100100011: color_data = Z;
		19'b0000100000100100100: color_data = Z;
		19'b0000100000100100101: color_data = Z;
		19'b0000100000100100110: color_data = Z;
		19'b0000100000100100111: color_data = Z;
		19'b0000100000100101000: color_data = Z;
		19'b0000100000100101001: color_data = Z;
		19'b0000100000100101010: color_data = Z;
		19'b0000100000100101011: color_data = Z;
		19'b0000100000100101100: color_data = Z;
		19'b0000100000100101101: color_data = Z;
		19'b0000100000100101110: color_data = Z;
		19'b0000100000100101111: color_data = Z;
		19'b0000100000100110000: color_data = Z;
		19'b0000100000100110001: color_data = Z;
		19'b0000100000100110010: color_data = Z;
		19'b0000100000100110011: color_data = Z;
		19'b0000100000100110100: color_data = Z;
		19'b0000100000100110101: color_data = Z;
		19'b0000100000100110110: color_data = Z;
		19'b0000100000100110111: color_data = Z;
		19'b0000100000100111000: color_data = Z;
		19'b0000100000100111001: color_data = Z;
		19'b0000100000100111010: color_data = Z;
		19'b0000100000100111011: color_data = Z;
		19'b0000100000100111100: color_data = Z;
		19'b0000100000100111101: color_data = Z;
		19'b0000100000100111110: color_data = Z;
		19'b0000100000100111111: color_data = Z;
		19'b0000100000101000000: color_data = Z;
		19'b0000100000101000001: color_data = Z;
		19'b0000100000101000010: color_data = Z;
		19'b0000100000101000011: color_data = Z;
		19'b0000100000101000100: color_data = Z;
		19'b0000100000101000101: color_data = Z;
		19'b0000100000101000110: color_data = Z;
		19'b0000100000101000111: color_data = Z;
		19'b0000100000101001000: color_data = Z;
		19'b0000100000101001001: color_data = Z;
		19'b0000100000101001010: color_data = Z;
		19'b0000100000101001011: color_data = Z;
		19'b0000100000101001100: color_data = Z;
		19'b0000100000101001101: color_data = Z;
		19'b0000100000101001110: color_data = Z;
		19'b0000100000101001111: color_data = Z;
		19'b0000100000101010000: color_data = Z;
		19'b0000100000101010001: color_data = Z;
		19'b0000100000101010010: color_data = Z;
		19'b0000100000101010011: color_data = Z;
		19'b0000100000101010100: color_data = Z;
		19'b0000100000101010101: color_data = Z;
		19'b0000100000101010110: color_data = Z;
		19'b0000100000101010111: color_data = Z;
		19'b0000100000101011000: color_data = Z;
		19'b0000100000101011001: color_data = Z;
		19'b0000100000101011010: color_data = Z;
		19'b0000100000101011011: color_data = Z;
		19'b0000100000101011100: color_data = Z;
		19'b0000100000101011101: color_data = Z;
		19'b0000100000101011110: color_data = Z;
		19'b0000100000101011111: color_data = Z;
		19'b0000100000101100000: color_data = Z;
		19'b0000100000101100001: color_data = Z;
		19'b0000100000101100010: color_data = Z;
		19'b0000100000101100011: color_data = Z;
		19'b0000100000101100100: color_data = Z;
		19'b0000100000101100101: color_data = Z;
		19'b0000100000101100110: color_data = Z;
		19'b0000100000101100111: color_data = Z;
		19'b0000100000101101000: color_data = Z;
		19'b0000100000101101001: color_data = Z;
		19'b0000100000101101010: color_data = Z;
		19'b0000100000101101011: color_data = Z;
		19'b0000100000101101100: color_data = Z;
		19'b0000100000101101101: color_data = Z;
		19'b0000100000101101110: color_data = Z;
		19'b0000100000101101111: color_data = Z;
		19'b0000100000101110000: color_data = Z;
		19'b0000100000101110001: color_data = Z;
		19'b0000100000101110010: color_data = Z;
		19'b0000100000101110011: color_data = Z;
		19'b0000100000101110100: color_data = Z;
		19'b0000100000101110101: color_data = Z;
		19'b0000100000101110110: color_data = Z;
		19'b0000100000101110111: color_data = Z;
		19'b0000100000101111000: color_data = Z;
		19'b0000100000101111001: color_data = Z;
		19'b0000100000101111010: color_data = Z;
		19'b0000100000101111011: color_data = Z;
		19'b0000100000101111100: color_data = Z;
		19'b0000100010100010101: color_data = Z;
		19'b0000100010100010110: color_data = Z;
		19'b0000100010100010111: color_data = Z;
		19'b0000100010100011000: color_data = Z;
		19'b0000100010100011001: color_data = Z;
		19'b0000100010100011010: color_data = Z;
		19'b0000100010100011011: color_data = Z;
		19'b0000100010100011100: color_data = Z;
		19'b0000100010100011101: color_data = Z;
		19'b0000100010100011110: color_data = Z;
		19'b0000100010100011111: color_data = Z;
		19'b0000100010100100000: color_data = Z;
		19'b0000100010100100001: color_data = Z;
		19'b0000100010100100010: color_data = Z;
		19'b0000100010100100011: color_data = Z;
		19'b0000100010100100100: color_data = Z;
		19'b0000100010100100101: color_data = Z;
		19'b0000100010100100110: color_data = Z;
		19'b0000100010100100111: color_data = Z;
		19'b0000100010100101000: color_data = Z;
		19'b0000100010100101001: color_data = Z;
		19'b0000100010100101010: color_data = Z;
		19'b0000100010100101011: color_data = Z;
		19'b0000100010100101100: color_data = Z;
		19'b0000100010100101101: color_data = Z;
		19'b0000100010100101110: color_data = Z;
		19'b0000100010100101111: color_data = Z;
		19'b0000100010100110000: color_data = Z;
		19'b0000100010100110001: color_data = Z;
		19'b0000100010100110010: color_data = Z;
		19'b0000100010100110011: color_data = Z;
		19'b0000100010100110100: color_data = Z;
		19'b0000100010100110101: color_data = Z;
		19'b0000100010100110110: color_data = Z;
		19'b0000100010100110111: color_data = Z;
		19'b0000100010100111000: color_data = Z;
		19'b0000100010100111001: color_data = Z;
		19'b0000100010100111010: color_data = Z;
		19'b0000100010100111011: color_data = Z;
		19'b0000100010100111100: color_data = Z;
		19'b0000100010100111101: color_data = Z;
		19'b0000100010100111110: color_data = Z;
		19'b0000100010100111111: color_data = Z;
		19'b0000100010101000000: color_data = Z;
		19'b0000100010101000001: color_data = Z;
		19'b0000100010101000010: color_data = Z;
		19'b0000100010101000011: color_data = Z;
		19'b0000100010101000100: color_data = Z;
		19'b0000100010101000101: color_data = Z;
		19'b0000100010101000110: color_data = Z;
		19'b0000100010101000111: color_data = Z;
		19'b0000100010101001000: color_data = Z;
		19'b0000100010101001001: color_data = Z;
		19'b0000100010101001010: color_data = Z;
		19'b0000100010101001011: color_data = Z;
		19'b0000100010101001100: color_data = Z;
		19'b0000100010101001101: color_data = Z;
		19'b0000100010101001110: color_data = Z;
		19'b0000100010101001111: color_data = Z;
		19'b0000100010101010000: color_data = Z;
		19'b0000100010101010001: color_data = Z;
		19'b0000100010101010010: color_data = Z;
		19'b0000100010101010011: color_data = Z;
		19'b0000100010101010100: color_data = Z;
		19'b0000100010101010101: color_data = Z;
		19'b0000100010101010110: color_data = Z;
		19'b0000100010101010111: color_data = Z;
		19'b0000100010101011000: color_data = Z;
		19'b0000100010101011001: color_data = Z;
		19'b0000100010101011010: color_data = Z;
		19'b0000100010101011011: color_data = Z;
		19'b0000100010101011100: color_data = Z;
		19'b0000100010101011101: color_data = Z;
		19'b0000100010101011110: color_data = Z;
		19'b0000100010101011111: color_data = Z;
		19'b0000100010101100000: color_data = Z;
		19'b0000100010101100001: color_data = Z;
		19'b0000100010101100010: color_data = Z;
		19'b0000100010101100011: color_data = Z;
		19'b0000100010101100100: color_data = Z;
		19'b0000100010101100101: color_data = Z;
		19'b0000100010101100110: color_data = Z;
		19'b0000100010101100111: color_data = Z;
		19'b0000100010101101000: color_data = Z;
		19'b0000100010101101001: color_data = Z;
		19'b0000100010101101010: color_data = Z;
		19'b0000100010101101011: color_data = Z;
		19'b0000100010101101100: color_data = Z;
		19'b0000100010101101101: color_data = Z;
		19'b0000100010101101110: color_data = Z;
		19'b0000100010101101111: color_data = Z;
		19'b0000100010101110000: color_data = Z;
		19'b0000100010101110001: color_data = Z;
		19'b0000100010101110010: color_data = Z;
		19'b0000100010101110011: color_data = Z;
		19'b0000100010101110100: color_data = Z;
		19'b0000100010101110101: color_data = Z;
		19'b0000100010101110110: color_data = Z;
		19'b0000100010101110111: color_data = Z;
		19'b0000100010101111000: color_data = Z;
		19'b0000100010101111001: color_data = Z;
		19'b0000100010101111010: color_data = Z;
		19'b0000100010101111011: color_data = Z;
		19'b0000100010101111100: color_data = Z;
		19'b0000100010101111101: color_data = Z;
		19'b0000100010101111110: color_data = Z;
		19'b0000100100100010010: color_data = Z;
		19'b0000100100100010011: color_data = Z;
		19'b0000100100100010100: color_data = Z;
		19'b0000100100100010101: color_data = Z;
		19'b0000100100100010110: color_data = Z;
		19'b0000100100100010111: color_data = Z;
		19'b0000100100100011000: color_data = Z;
		19'b0000100100100011001: color_data = Z;
		19'b0000100100100011010: color_data = Z;
		19'b0000100100100011011: color_data = Z;
		19'b0000100100100011100: color_data = Z;
		19'b0000100100100011101: color_data = Z;
		19'b0000100100100011110: color_data = Z;
		19'b0000100100100011111: color_data = Z;
		19'b0000100100100100000: color_data = Z;
		19'b0000100100100100001: color_data = Z;
		19'b0000100100100100010: color_data = Z;
		19'b0000100100100100011: color_data = Z;
		19'b0000100100100100100: color_data = Z;
		19'b0000100100100100101: color_data = Z;
		19'b0000100100100100110: color_data = Z;
		19'b0000100100100100111: color_data = Z;
		19'b0000100100100101000: color_data = Z;
		19'b0000100100100101001: color_data = Z;
		19'b0000100100100101010: color_data = Z;
		19'b0000100100100101011: color_data = Z;
		19'b0000100100100101100: color_data = Z;
		19'b0000100100100101101: color_data = Z;
		19'b0000100100100101110: color_data = Z;
		19'b0000100100100101111: color_data = Z;
		19'b0000100100100110000: color_data = Z;
		19'b0000100100100110001: color_data = Z;
		19'b0000100100100110010: color_data = Z;
		19'b0000100100100110011: color_data = Z;
		19'b0000100100100110100: color_data = Z;
		19'b0000100100100110101: color_data = Z;
		19'b0000100100100110110: color_data = Z;
		19'b0000100100100110111: color_data = Z;
		19'b0000100100100111000: color_data = Z;
		19'b0000100100100111001: color_data = Z;
		19'b0000100100100111010: color_data = Z;
		19'b0000100100100111011: color_data = Z;
		19'b0000100100100111100: color_data = Z;
		19'b0000100100100111101: color_data = Z;
		19'b0000100100100111110: color_data = Z;
		19'b0000100100100111111: color_data = Z;
		19'b0000100100101000000: color_data = Z;
		19'b0000100100101000001: color_data = Z;
		19'b0000100100101000010: color_data = Z;
		19'b0000100100101000011: color_data = Z;
		19'b0000100100101000100: color_data = Z;
		19'b0000100100101000101: color_data = Z;
		19'b0000100100101000110: color_data = Z;
		19'b0000100100101000111: color_data = Z;
		19'b0000100100101001000: color_data = Z;
		19'b0000100100101001001: color_data = Z;
		19'b0000100100101001010: color_data = Z;
		19'b0000100100101001011: color_data = Z;
		19'b0000100100101001100: color_data = Z;
		19'b0000100100101001101: color_data = Z;
		19'b0000100100101001110: color_data = Z;
		19'b0000100100101001111: color_data = Z;
		19'b0000100100101010000: color_data = Z;
		19'b0000100100101010001: color_data = Z;
		19'b0000100100101010010: color_data = Z;
		19'b0000100100101010011: color_data = Z;
		19'b0000100100101010100: color_data = Z;
		19'b0000100100101010101: color_data = Z;
		19'b0000100100101010110: color_data = Z;
		19'b0000100100101010111: color_data = Z;
		19'b0000100100101011000: color_data = Z;
		19'b0000100100101011001: color_data = Z;
		19'b0000100100101011010: color_data = Z;
		19'b0000100100101011011: color_data = Z;
		19'b0000100100101011100: color_data = Z;
		19'b0000100100101011101: color_data = Z;
		19'b0000100100101011110: color_data = Z;
		19'b0000100100101011111: color_data = Z;
		19'b0000100100101100000: color_data = Z;
		19'b0000100100101100001: color_data = Z;
		19'b0000100100101100010: color_data = Z;
		19'b0000100100101100011: color_data = Z;
		19'b0000100100101100100: color_data = Z;
		19'b0000100100101100101: color_data = Z;
		19'b0000100100101100110: color_data = Z;
		19'b0000100100101100111: color_data = Z;
		19'b0000100100101101000: color_data = Z;
		19'b0000100100101101001: color_data = Z;
		19'b0000100100101101010: color_data = Z;
		19'b0000100100101101011: color_data = Z;
		19'b0000100100101101100: color_data = Z;
		19'b0000100100101101101: color_data = Z;
		19'b0000100100101101110: color_data = Z;
		19'b0000100100101101111: color_data = Z;
		19'b0000100100101110000: color_data = Z;
		19'b0000100100101110001: color_data = Z;
		19'b0000100100101110010: color_data = Z;
		19'b0000100100101110011: color_data = Z;
		19'b0000100100101110100: color_data = Z;
		19'b0000100100101110101: color_data = Z;
		19'b0000100100101110110: color_data = Z;
		19'b0000100100101110111: color_data = Z;
		19'b0000100100101111000: color_data = Z;
		19'b0000100100101111001: color_data = Z;
		19'b0000100100101111010: color_data = Z;
		19'b0000100100101111011: color_data = Z;
		19'b0000100100101111100: color_data = Z;
		19'b0000100100101111101: color_data = Z;
		19'b0000100100101111110: color_data = Z;
		19'b0000100100101111111: color_data = Z;
		19'b0000100100110000000: color_data = Z;
		19'b0000100110100010000: color_data = Z;
		19'b0000100110100010001: color_data = Z;
		19'b0000100110100010010: color_data = Z;
		19'b0000100110100010011: color_data = Z;
		19'b0000100110100010100: color_data = Z;
		19'b0000100110100010101: color_data = Z;
		19'b0000100110100010110: color_data = Z;
		19'b0000100110100010111: color_data = Z;
		19'b0000100110100011000: color_data = Z;
		19'b0000100110100011001: color_data = Z;
		19'b0000100110100011010: color_data = Z;
		19'b0000100110100011011: color_data = Z;
		19'b0000100110100011100: color_data = Z;
		19'b0000100110100011101: color_data = Z;
		19'b0000100110100011110: color_data = Z;
		19'b0000100110100011111: color_data = Z;
		19'b0000100110100100000: color_data = Z;
		19'b0000100110100100001: color_data = Z;
		19'b0000100110100100010: color_data = Z;
		19'b0000100110100100011: color_data = Z;
		19'b0000100110100100100: color_data = Z;
		19'b0000100110100100101: color_data = Z;
		19'b0000100110100100110: color_data = Z;
		19'b0000100110100100111: color_data = Z;
		19'b0000100110100101000: color_data = Z;
		19'b0000100110100101001: color_data = Z;
		19'b0000100110100101010: color_data = Z;
		19'b0000100110100101011: color_data = Z;
		19'b0000100110100101100: color_data = Z;
		19'b0000100110100101101: color_data = Z;
		19'b0000100110100101110: color_data = Z;
		19'b0000100110100101111: color_data = Z;
		19'b0000100110100110000: color_data = Z;
		19'b0000100110100110001: color_data = Z;
		19'b0000100110100110010: color_data = Z;
		19'b0000100110100110011: color_data = Z;
		19'b0000100110100110100: color_data = Z;
		19'b0000100110100110101: color_data = Z;
		19'b0000100110100110110: color_data = Z;
		19'b0000100110100110111: color_data = Z;
		19'b0000100110100111000: color_data = Z;
		19'b0000100110100111001: color_data = Z;
		19'b0000100110100111010: color_data = Z;
		19'b0000100110100111011: color_data = Z;
		19'b0000100110100111100: color_data = Z;
		19'b0000100110100111101: color_data = Z;
		19'b0000100110100111110: color_data = Z;
		19'b0000100110100111111: color_data = Z;
		19'b0000100110101000000: color_data = Z;
		19'b0000100110101000001: color_data = Z;
		19'b0000100110101000010: color_data = Z;
		19'b0000100110101000011: color_data = Z;
		19'b0000100110101000100: color_data = Z;
		19'b0000100110101000101: color_data = Z;
		19'b0000100110101000110: color_data = Z;
		19'b0000100110101000111: color_data = Z;
		19'b0000100110101001000: color_data = Z;
		19'b0000100110101001001: color_data = Z;
		19'b0000100110101001010: color_data = Z;
		19'b0000100110101001011: color_data = Z;
		19'b0000100110101001100: color_data = Z;
		19'b0000100110101001101: color_data = Z;
		19'b0000100110101001110: color_data = Z;
		19'b0000100110101001111: color_data = Z;
		19'b0000100110101010000: color_data = Z;
		19'b0000100110101010001: color_data = Z;
		19'b0000100110101010010: color_data = Z;
		19'b0000100110101010011: color_data = Z;
		19'b0000100110101010100: color_data = Z;
		19'b0000100110101010101: color_data = Z;
		19'b0000100110101010110: color_data = Z;
		19'b0000100110101010111: color_data = Z;
		19'b0000100110101011000: color_data = Z;
		19'b0000100110101011001: color_data = Z;
		19'b0000100110101011010: color_data = Z;
		19'b0000100110101011011: color_data = Z;
		19'b0000100110101011100: color_data = Z;
		19'b0000100110101011101: color_data = Z;
		19'b0000100110101011110: color_data = Z;
		19'b0000100110101011111: color_data = Z;
		19'b0000100110101100000: color_data = Z;
		19'b0000100110101100001: color_data = Z;
		19'b0000100110101100010: color_data = Z;
		19'b0000100110101100011: color_data = Z;
		19'b0000100110101100100: color_data = Z;
		19'b0000100110101100101: color_data = Z;
		19'b0000100110101100110: color_data = Z;
		19'b0000100110101100111: color_data = Z;
		19'b0000100110101101000: color_data = Z;
		19'b0000100110101101001: color_data = Z;
		19'b0000100110101101010: color_data = Z;
		19'b0000100110101101011: color_data = Z;
		19'b0000100110101101100: color_data = Z;
		19'b0000100110101101101: color_data = Z;
		19'b0000100110101101110: color_data = Z;
		19'b0000100110101101111: color_data = Z;
		19'b0000100110101110000: color_data = Z;
		19'b0000100110101110001: color_data = Z;
		19'b0000100110101110010: color_data = Z;
		19'b0000100110101110011: color_data = Z;
		19'b0000100110101110100: color_data = Z;
		19'b0000100110101110101: color_data = Z;
		19'b0000100110101110110: color_data = Z;
		19'b0000100110101110111: color_data = Z;
		19'b0000100110101111000: color_data = Z;
		19'b0000100110101111001: color_data = Z;
		19'b0000100110101111010: color_data = Z;
		19'b0000100110101111011: color_data = Z;
		19'b0000100110101111100: color_data = Z;
		19'b0000100110101111101: color_data = Z;
		19'b0000100110101111110: color_data = Z;
		19'b0000100110101111111: color_data = Z;
		19'b0000100110110000000: color_data = Z;
		19'b0000100110110000001: color_data = Z;
		19'b0000100110110000010: color_data = Z;
		19'b0000100110110000011: color_data = Z;
		19'b0000101000100001101: color_data = Z;
		19'b0000101000100001110: color_data = Z;
		19'b0000101000100001111: color_data = Z;
		19'b0000101000100010000: color_data = Z;
		19'b0000101000100010001: color_data = Z;
		19'b0000101000100010010: color_data = Z;
		19'b0000101000100010011: color_data = Z;
		19'b0000101000100010100: color_data = Z;
		19'b0000101000100010101: color_data = Z;
		19'b0000101000100010110: color_data = Z;
		19'b0000101000100010111: color_data = Z;
		19'b0000101000100011000: color_data = Z;
		19'b0000101000100011001: color_data = Z;
		19'b0000101000100011010: color_data = Z;
		19'b0000101000100011011: color_data = Z;
		19'b0000101000100011100: color_data = Z;
		19'b0000101000100011101: color_data = Z;
		19'b0000101000100011110: color_data = Z;
		19'b0000101000100011111: color_data = Z;
		19'b0000101000100100000: color_data = Z;
		19'b0000101000100100001: color_data = Z;
		19'b0000101000100100010: color_data = Z;
		19'b0000101000100100011: color_data = Z;
		19'b0000101000100100100: color_data = Z;
		19'b0000101000100100101: color_data = Z;
		19'b0000101000100100110: color_data = Z;
		19'b0000101000100100111: color_data = Z;
		19'b0000101000100101000: color_data = Z;
		19'b0000101000100101001: color_data = Z;
		19'b0000101000100101010: color_data = Z;
		19'b0000101000100101011: color_data = Z;
		19'b0000101000100101100: color_data = Z;
		19'b0000101000100101101: color_data = Z;
		19'b0000101000100101110: color_data = Z;
		19'b0000101000100101111: color_data = Z;
		19'b0000101000100110000: color_data = Z;
		19'b0000101000100110001: color_data = Z;
		19'b0000101000100110010: color_data = Z;
		19'b0000101000100110011: color_data = Z;
		19'b0000101000100110100: color_data = Z;
		19'b0000101000100110101: color_data = Z;
		19'b0000101000100110110: color_data = Z;
		19'b0000101000100110111: color_data = Z;
		19'b0000101000100111000: color_data = Z;
		19'b0000101000100111001: color_data = Z;
		19'b0000101000100111010: color_data = Z;
		19'b0000101000100111011: color_data = Z;
		19'b0000101000100111100: color_data = Z;
		19'b0000101000100111101: color_data = Z;
		19'b0000101000100111110: color_data = Z;
		19'b0000101000100111111: color_data = Z;
		19'b0000101000101000000: color_data = Z;
		19'b0000101000101000001: color_data = Z;
		19'b0000101000101000010: color_data = Z;
		19'b0000101000101000011: color_data = Z;
		19'b0000101000101000100: color_data = Z;
		19'b0000101000101000101: color_data = Z;
		19'b0000101000101000110: color_data = Z;
		19'b0000101000101000111: color_data = Z;
		19'b0000101000101001000: color_data = Z;
		19'b0000101000101001001: color_data = Z;
		19'b0000101000101001010: color_data = Z;
		19'b0000101000101001011: color_data = Z;
		19'b0000101000101001100: color_data = Z;
		19'b0000101000101001101: color_data = Z;
		19'b0000101000101001110: color_data = Z;
		19'b0000101000101001111: color_data = Z;
		19'b0000101000101010000: color_data = Z;
		19'b0000101000101010001: color_data = Z;
		19'b0000101000101010010: color_data = Z;
		19'b0000101000101010011: color_data = Z;
		19'b0000101000101010100: color_data = Z;
		19'b0000101000101010101: color_data = Z;
		19'b0000101000101010110: color_data = Z;
		19'b0000101000101010111: color_data = Z;
		19'b0000101000101011000: color_data = Z;
		19'b0000101000101011001: color_data = Z;
		19'b0000101000101011010: color_data = Z;
		19'b0000101000101011011: color_data = Z;
		19'b0000101000101011100: color_data = Z;
		19'b0000101000101011101: color_data = Z;
		19'b0000101000101011110: color_data = Z;
		19'b0000101000101011111: color_data = Z;
		19'b0000101000101100000: color_data = Z;
		19'b0000101000101100001: color_data = Z;
		19'b0000101000101100010: color_data = Z;
		19'b0000101000101100011: color_data = Z;
		19'b0000101000101100100: color_data = Z;
		19'b0000101000101100101: color_data = Z;
		19'b0000101000101100110: color_data = Z;
		19'b0000101000101100111: color_data = Z;
		19'b0000101000101101000: color_data = Z;
		19'b0000101000101101001: color_data = Z;
		19'b0000101000101101010: color_data = Z;
		19'b0000101000101101011: color_data = Z;
		19'b0000101000101101100: color_data = Z;
		19'b0000101000101101101: color_data = Z;
		19'b0000101000101101110: color_data = Z;
		19'b0000101000101101111: color_data = Z;
		19'b0000101000101110000: color_data = Z;
		19'b0000101000101110001: color_data = Z;
		19'b0000101000101110010: color_data = Z;
		19'b0000101000101110011: color_data = Z;
		19'b0000101000101110100: color_data = Z;
		19'b0000101000101110101: color_data = Z;
		19'b0000101000101110110: color_data = Z;
		19'b0000101000101110111: color_data = Z;
		19'b0000101000101111000: color_data = Z;
		19'b0000101000101111001: color_data = Z;
		19'b0000101000101111010: color_data = Z;
		19'b0000101000101111011: color_data = Z;
		19'b0000101000101111100: color_data = Z;
		19'b0000101000101111101: color_data = Z;
		19'b0000101000101111110: color_data = Z;
		19'b0000101000101111111: color_data = Z;
		19'b0000101000110000000: color_data = Z;
		19'b0000101000110000001: color_data = Z;
		19'b0000101000110000010: color_data = Z;
		19'b0000101000110000011: color_data = Z;
		19'b0000101000110000100: color_data = Z;
		19'b0000101000110000101: color_data = Z;
		19'b0000101000110000110: color_data = Z;
		19'b0000101010100001100: color_data = Z;
		19'b0000101010100001101: color_data = Z;
		19'b0000101010100001110: color_data = Z;
		19'b0000101010100001111: color_data = Z;
		19'b0000101010100010000: color_data = Z;
		19'b0000101010100010001: color_data = Z;
		19'b0000101010100010010: color_data = Z;
		19'b0000101010100010011: color_data = Z;
		19'b0000101010100010100: color_data = Z;
		19'b0000101010100010101: color_data = Z;
		19'b0000101010100010110: color_data = Z;
		19'b0000101010100010111: color_data = Z;
		19'b0000101010100011000: color_data = Z;
		19'b0000101010100011001: color_data = Z;
		19'b0000101010100011010: color_data = Z;
		19'b0000101010100011011: color_data = Z;
		19'b0000101010100011100: color_data = Z;
		19'b0000101010100011101: color_data = Z;
		19'b0000101010100011110: color_data = Z;
		19'b0000101010100011111: color_data = Z;
		19'b0000101010100100000: color_data = Z;
		19'b0000101010100100001: color_data = Z;
		19'b0000101010100100010: color_data = Z;
		19'b0000101010100100011: color_data = Z;
		19'b0000101010100100100: color_data = Z;
		19'b0000101010100100101: color_data = Z;
		19'b0000101010100100110: color_data = Z;
		19'b0000101010100100111: color_data = Z;
		19'b0000101010100101000: color_data = Z;
		19'b0000101010100101001: color_data = Z;
		19'b0000101010100101010: color_data = Z;
		19'b0000101010100101011: color_data = Z;
		19'b0000101010100101100: color_data = Z;
		19'b0000101010100101101: color_data = Z;
		19'b0000101010100101110: color_data = Z;
		19'b0000101010100101111: color_data = Z;
		19'b0000101010100110000: color_data = Z;
		19'b0000101010100110001: color_data = Z;
		19'b0000101010100110010: color_data = Z;
		19'b0000101010100110011: color_data = Z;
		19'b0000101010100110100: color_data = Z;
		19'b0000101010100110101: color_data = Z;
		19'b0000101010100110110: color_data = Z;
		19'b0000101010100110111: color_data = Z;
		19'b0000101010100111000: color_data = Z;
		19'b0000101010100111001: color_data = Z;
		19'b0000101010100111010: color_data = Z;
		19'b0000101010100111011: color_data = Z;
		19'b0000101010100111100: color_data = Z;
		19'b0000101010100111101: color_data = Z;
		19'b0000101010100111110: color_data = Z;
		19'b0000101010100111111: color_data = Z;
		19'b0000101010101000000: color_data = Z;
		19'b0000101010101000001: color_data = Z;
		19'b0000101010101000010: color_data = Z;
		19'b0000101010101000011: color_data = Z;
		19'b0000101010101000100: color_data = Z;
		19'b0000101010101000101: color_data = Z;
		19'b0000101010101000110: color_data = Z;
		19'b0000101010101000111: color_data = Z;
		19'b0000101010101001000: color_data = Z;
		19'b0000101010101001001: color_data = Z;
		19'b0000101010101001010: color_data = Z;
		19'b0000101010101001011: color_data = Z;
		19'b0000101010101001100: color_data = Z;
		19'b0000101010101001101: color_data = Z;
		19'b0000101010101001110: color_data = Z;
		19'b0000101010101001111: color_data = Z;
		19'b0000101010101010000: color_data = Z;
		19'b0000101010101010001: color_data = Z;
		19'b0000101010101010010: color_data = Z;
		19'b0000101010101010011: color_data = Z;
		19'b0000101010101010100: color_data = Z;
		19'b0000101010101010101: color_data = Z;
		19'b0000101010101010110: color_data = Z;
		19'b0000101010101010111: color_data = Z;
		19'b0000101010101011000: color_data = Z;
		19'b0000101010101011001: color_data = Z;
		19'b0000101010101011010: color_data = Z;
		19'b0000101010101011011: color_data = Z;
		19'b0000101010101011100: color_data = Z;
		19'b0000101010101011101: color_data = Z;
		19'b0000101010101011110: color_data = Z;
		19'b0000101010101011111: color_data = Z;
		19'b0000101010101100000: color_data = Z;
		19'b0000101010101100001: color_data = Z;
		19'b0000101010101100010: color_data = Z;
		19'b0000101010101100011: color_data = Z;
		19'b0000101010101100100: color_data = Z;
		19'b0000101010101100101: color_data = Z;
		19'b0000101010101100110: color_data = Z;
		19'b0000101010101100111: color_data = Z;
		19'b0000101010101101000: color_data = Z;
		19'b0000101010101101001: color_data = Z;
		19'b0000101010101101010: color_data = Z;
		19'b0000101010101101011: color_data = Z;
		19'b0000101010101101100: color_data = Z;
		19'b0000101010101101101: color_data = Z;
		19'b0000101010101101110: color_data = Z;
		19'b0000101010101101111: color_data = Z;
		19'b0000101010101110000: color_data = Z;
		19'b0000101010101110001: color_data = Z;
		19'b0000101010101110010: color_data = Z;
		19'b0000101010101110011: color_data = Z;
		19'b0000101010101110100: color_data = Z;
		19'b0000101010101110101: color_data = Z;
		19'b0000101010101110110: color_data = Z;
		19'b0000101010101110111: color_data = Z;
		19'b0000101010101111000: color_data = Z;
		19'b0000101010101111001: color_data = Z;
		19'b0000101010101111010: color_data = Z;
		19'b0000101010101111011: color_data = Z;
		19'b0000101010101111100: color_data = Z;
		19'b0000101010101111101: color_data = Z;
		19'b0000101010101111110: color_data = Z;
		19'b0000101010101111111: color_data = Z;
		19'b0000101010110000000: color_data = Z;
		19'b0000101010110000001: color_data = Z;
		19'b0000101010110000010: color_data = Z;
		19'b0000101010110000011: color_data = Z;
		19'b0000101010110000100: color_data = Z;
		19'b0000101010110000101: color_data = Z;
		19'b0000101010110000110: color_data = Z;
		19'b0000101010110000111: color_data = Z;
		19'b0000101010110001000: color_data = Z;
		19'b0000101100100001010: color_data = Z;
		19'b0000101100100001011: color_data = Z;
		19'b0000101100100001100: color_data = Z;
		19'b0000101100100001101: color_data = Z;
		19'b0000101100100001110: color_data = Z;
		19'b0000101100100001111: color_data = Z;
		19'b0000101100100010000: color_data = Z;
		19'b0000101100100010001: color_data = Z;
		19'b0000101100100010010: color_data = Z;
		19'b0000101100100010011: color_data = Z;
		19'b0000101100100010100: color_data = Z;
		19'b0000101100100010101: color_data = Z;
		19'b0000101100100010110: color_data = Z;
		19'b0000101100100010111: color_data = Z;
		19'b0000101100100011000: color_data = Z;
		19'b0000101100100011001: color_data = Z;
		19'b0000101100100011010: color_data = Z;
		19'b0000101100100011011: color_data = Z;
		19'b0000101100100011100: color_data = Z;
		19'b0000101100100011101: color_data = Z;
		19'b0000101100100011110: color_data = Z;
		19'b0000101100100011111: color_data = Z;
		19'b0000101100100100000: color_data = Z;
		19'b0000101100100100001: color_data = Z;
		19'b0000101100100100010: color_data = Z;
		19'b0000101100100100011: color_data = Z;
		19'b0000101100100100100: color_data = Z;
		19'b0000101100100100101: color_data = Z;
		19'b0000101100100100110: color_data = Z;
		19'b0000101100100100111: color_data = Z;
		19'b0000101100100101000: color_data = Z;
		19'b0000101100100101001: color_data = Z;
		19'b0000101100100101010: color_data = Z;
		19'b0000101100100101011: color_data = Z;
		19'b0000101100100101100: color_data = Z;
		19'b0000101100100101101: color_data = Z;
		19'b0000101100100101110: color_data = Z;
		19'b0000101100100101111: color_data = Z;
		19'b0000101100100110000: color_data = Z;
		19'b0000101100100110001: color_data = Z;
		19'b0000101100100110010: color_data = Z;
		19'b0000101100100110011: color_data = Z;
		19'b0000101100100110100: color_data = Z;
		19'b0000101100100110101: color_data = Z;
		19'b0000101100100110110: color_data = Z;
		19'b0000101100100110111: color_data = Z;
		19'b0000101100100111000: color_data = Z;
		19'b0000101100100111001: color_data = Z;
		19'b0000101100100111010: color_data = Z;
		19'b0000101100100111011: color_data = Z;
		19'b0000101100100111100: color_data = Z;
		19'b0000101100100111101: color_data = Z;
		19'b0000101100100111110: color_data = Z;
		19'b0000101100100111111: color_data = Z;
		19'b0000101100101000000: color_data = Z;
		19'b0000101100101000001: color_data = Z;
		19'b0000101100101000010: color_data = Z;
		19'b0000101100101000011: color_data = Z;
		19'b0000101100101000100: color_data = Z;
		19'b0000101100101000101: color_data = Z;
		19'b0000101100101000110: color_data = Z;
		19'b0000101100101000111: color_data = Z;
		19'b0000101100101001000: color_data = Z;
		19'b0000101100101001001: color_data = Z;
		19'b0000101100101001010: color_data = Z;
		19'b0000101100101001011: color_data = Z;
		19'b0000101100101001100: color_data = Z;
		19'b0000101100101001101: color_data = Z;
		19'b0000101100101001110: color_data = Z;
		19'b0000101100101001111: color_data = Z;
		19'b0000101100101010000: color_data = Z;
		19'b0000101100101010001: color_data = Z;
		19'b0000101100101010010: color_data = Z;
		19'b0000101100101010011: color_data = Z;
		19'b0000101100101010100: color_data = Z;
		19'b0000101100101010101: color_data = Z;
		19'b0000101100101010110: color_data = Z;
		19'b0000101100101010111: color_data = Z;
		19'b0000101100101011000: color_data = Z;
		19'b0000101100101011001: color_data = Z;
		19'b0000101100101011010: color_data = Z;
		19'b0000101100101011011: color_data = Z;
		19'b0000101100101011100: color_data = Z;
		19'b0000101100101011101: color_data = Z;
		19'b0000101100101011110: color_data = Z;
		19'b0000101100101011111: color_data = Z;
		19'b0000101100101100000: color_data = Z;
		19'b0000101100101100001: color_data = Z;
		19'b0000101100101100010: color_data = Z;
		19'b0000101100101100011: color_data = Z;
		19'b0000101100101100100: color_data = Z;
		19'b0000101100101100101: color_data = Z;
		19'b0000101100101100110: color_data = Z;
		19'b0000101100101100111: color_data = Z;
		19'b0000101100101101000: color_data = Z;
		19'b0000101100101101001: color_data = Z;
		19'b0000101100101101010: color_data = Z;
		19'b0000101100101101011: color_data = Z;
		19'b0000101100101101100: color_data = Z;
		19'b0000101100101101101: color_data = Z;
		19'b0000101100101101110: color_data = Z;
		19'b0000101100101101111: color_data = Z;
		19'b0000101100101110000: color_data = Z;
		19'b0000101100101110001: color_data = Z;
		19'b0000101100101110010: color_data = Z;
		19'b0000101100101110011: color_data = Z;
		19'b0000101100101110100: color_data = Z;
		19'b0000101100101110101: color_data = Z;
		19'b0000101100101110110: color_data = Z;
		19'b0000101100101110111: color_data = Z;
		19'b0000101100101111000: color_data = Z;
		19'b0000101100101111001: color_data = Z;
		19'b0000101100101111010: color_data = Z;
		19'b0000101100101111011: color_data = Z;
		19'b0000101100101111100: color_data = Z;
		19'b0000101100101111101: color_data = Z;
		19'b0000101100101111110: color_data = Z;
		19'b0000101100101111111: color_data = Z;
		19'b0000101100110000000: color_data = Z;
		19'b0000101100110000001: color_data = Z;
		19'b0000101100110000010: color_data = Z;
		19'b0000101100110000011: color_data = Z;
		19'b0000101100110000100: color_data = Z;
		19'b0000101100110000101: color_data = Z;
		19'b0000101100110000110: color_data = Z;
		19'b0000101100110000111: color_data = Z;
		19'b0000101100110001000: color_data = Z;
		19'b0000101100110001001: color_data = Z;
		19'b0000101100110001010: color_data = Z;
		19'b0000101110100000110: color_data = Z;
		19'b0000101110100001000: color_data = Z;
		19'b0000101110100001001: color_data = Z;
		19'b0000101110100001010: color_data = Z;
		19'b0000101110100001011: color_data = Z;
		19'b0000101110100001100: color_data = Z;
		19'b0000101110100001101: color_data = Z;
		19'b0000101110100001110: color_data = Z;
		19'b0000101110100001111: color_data = Z;
		19'b0000101110100010000: color_data = Z;
		19'b0000101110100010001: color_data = Z;
		19'b0000101110100010010: color_data = Z;
		19'b0000101110100010011: color_data = Z;
		19'b0000101110100010100: color_data = Z;
		19'b0000101110100010101: color_data = Z;
		19'b0000101110100010110: color_data = Z;
		19'b0000101110100010111: color_data = Z;
		19'b0000101110100011000: color_data = Z;
		19'b0000101110100011001: color_data = Z;
		19'b0000101110100011010: color_data = Z;
		19'b0000101110100011011: color_data = Z;
		19'b0000101110100011100: color_data = Z;
		19'b0000101110100011101: color_data = Z;
		19'b0000101110100011110: color_data = Z;
		19'b0000101110100011111: color_data = Z;
		19'b0000101110100100000: color_data = Z;
		19'b0000101110100100001: color_data = Z;
		19'b0000101110100100010: color_data = Z;
		19'b0000101110100100011: color_data = Z;
		19'b0000101110100100100: color_data = Z;
		19'b0000101110100100101: color_data = Z;
		19'b0000101110100100110: color_data = Z;
		19'b0000101110100100111: color_data = Z;
		19'b0000101110100101000: color_data = Z;
		19'b0000101110100101001: color_data = Z;
		19'b0000101110100101010: color_data = Z;
		19'b0000101110100101011: color_data = Z;
		19'b0000101110100101100: color_data = Z;
		19'b0000101110100101101: color_data = Z;
		19'b0000101110100101110: color_data = Z;
		19'b0000101110100101111: color_data = Z;
		19'b0000101110100110000: color_data = Z;
		19'b0000101110100110001: color_data = Z;
		19'b0000101110100110010: color_data = Z;
		19'b0000101110100110011: color_data = Z;
		19'b0000101110100110100: color_data = Z;
		19'b0000101110100110101: color_data = Z;
		19'b0000101110100110110: color_data = Z;
		19'b0000101110100110111: color_data = Z;
		19'b0000101110100111000: color_data = Z;
		19'b0000101110100111001: color_data = Z;
		19'b0000101110100111010: color_data = Z;
		19'b0000101110100111011: color_data = Z;
		19'b0000101110100111100: color_data = Z;
		19'b0000101110100111101: color_data = Z;
		19'b0000101110100111110: color_data = Z;
		19'b0000101110100111111: color_data = Z;
		19'b0000101110101000000: color_data = Z;
		19'b0000101110101000001: color_data = Z;
		19'b0000101110101000010: color_data = Z;
		19'b0000101110101000011: color_data = Z;
		19'b0000101110101000100: color_data = Z;
		19'b0000101110101000101: color_data = Z;
		19'b0000101110101000110: color_data = Z;
		19'b0000101110101000111: color_data = Z;
		19'b0000101110101001000: color_data = Z;
		19'b0000101110101001001: color_data = Z;
		19'b0000101110101001010: color_data = Z;
		19'b0000101110101001011: color_data = Z;
		19'b0000101110101001100: color_data = Z;
		19'b0000101110101001101: color_data = Z;
		19'b0000101110101001110: color_data = Z;
		19'b0000101110101001111: color_data = Z;
		19'b0000101110101010000: color_data = Z;
		19'b0000101110101010001: color_data = Z;
		19'b0000101110101010010: color_data = Z;
		19'b0000101110101010011: color_data = Z;
		19'b0000101110101010100: color_data = Z;
		19'b0000101110101010101: color_data = Z;
		19'b0000101110101010110: color_data = Z;
		19'b0000101110101010111: color_data = Z;
		19'b0000101110101011000: color_data = Z;
		19'b0000101110101011001: color_data = Z;
		19'b0000101110101011010: color_data = Z;
		19'b0000101110101011011: color_data = Z;
		19'b0000101110101011100: color_data = Z;
		19'b0000101110101011101: color_data = Z;
		19'b0000101110101011110: color_data = Z;
		19'b0000101110101011111: color_data = Z;
		19'b0000101110101100000: color_data = Z;
		19'b0000101110101100001: color_data = Z;
		19'b0000101110101100010: color_data = Z;
		19'b0000101110101100011: color_data = Z;
		19'b0000101110101100100: color_data = Z;
		19'b0000101110101100101: color_data = Z;
		19'b0000101110101100110: color_data = Z;
		19'b0000101110101100111: color_data = Z;
		19'b0000101110101101000: color_data = Z;
		19'b0000101110101101001: color_data = Z;
		19'b0000101110101101010: color_data = Z;
		19'b0000101110101101011: color_data = Z;
		19'b0000101110101101100: color_data = Z;
		19'b0000101110101101101: color_data = Z;
		19'b0000101110101101110: color_data = Z;
		19'b0000101110101101111: color_data = Z;
		19'b0000101110101110000: color_data = Z;
		19'b0000101110101110001: color_data = Z;
		19'b0000101110101110010: color_data = Z;
		19'b0000101110101110011: color_data = Z;
		19'b0000101110101110100: color_data = Z;
		19'b0000101110101110101: color_data = Z;
		19'b0000101110101110110: color_data = Z;
		19'b0000101110101110111: color_data = Z;
		19'b0000101110101111000: color_data = Z;
		19'b0000101110101111001: color_data = Z;
		19'b0000101110101111010: color_data = Z;
		19'b0000101110101111011: color_data = Z;
		19'b0000101110101111100: color_data = Z;
		19'b0000101110101111101: color_data = Z;
		19'b0000101110101111110: color_data = Z;
		19'b0000101110101111111: color_data = Z;
		19'b0000101110110000000: color_data = Z;
		19'b0000101110110000001: color_data = Z;
		19'b0000101110110000010: color_data = Z;
		19'b0000101110110000011: color_data = Z;
		19'b0000101110110000100: color_data = Z;
		19'b0000101110110000101: color_data = Z;
		19'b0000101110110000110: color_data = Z;
		19'b0000101110110000111: color_data = Z;
		19'b0000101110110001000: color_data = Z;
		19'b0000101110110001001: color_data = Z;
		19'b0000101110110001010: color_data = Z;
		19'b0000101110110001011: color_data = Z;
		19'b0000110000100000110: color_data = Z;
		19'b0000110000100000111: color_data = Z;
		19'b0000110000100001000: color_data = Z;
		19'b0000110000100001001: color_data = Z;
		19'b0000110000100001010: color_data = Z;
		19'b0000110000100001011: color_data = Z;
		19'b0000110000100001100: color_data = Z;
		19'b0000110000100001101: color_data = Z;
		19'b0000110000100001110: color_data = Z;
		19'b0000110000100001111: color_data = Z;
		19'b0000110000100010000: color_data = Z;
		19'b0000110000100010001: color_data = Z;
		19'b0000110000100010010: color_data = Z;
		19'b0000110000100010011: color_data = Z;
		19'b0000110000100010100: color_data = Z;
		19'b0000110000100010101: color_data = Z;
		19'b0000110000100010110: color_data = Z;
		19'b0000110000100010111: color_data = Z;
		19'b0000110000100011000: color_data = Z;
		19'b0000110000100011001: color_data = Z;
		19'b0000110000100011010: color_data = Z;
		19'b0000110000100011011: color_data = Z;
		19'b0000110000100011100: color_data = Z;
		19'b0000110000100011101: color_data = Z;
		19'b0000110000100011110: color_data = Z;
		19'b0000110000100011111: color_data = Z;
		19'b0000110000100100000: color_data = Z;
		19'b0000110000100100001: color_data = Z;
		19'b0000110000100100010: color_data = Z;
		19'b0000110000100100011: color_data = Z;
		19'b0000110000100100100: color_data = Z;
		19'b0000110000100100101: color_data = Z;
		19'b0000110000100100110: color_data = Z;
		19'b0000110000100100111: color_data = Z;
		19'b0000110000100101000: color_data = Z;
		19'b0000110000100101001: color_data = Z;
		19'b0000110000100101010: color_data = Z;
		19'b0000110000100101011: color_data = Z;
		19'b0000110000100101100: color_data = Z;
		19'b0000110000100101101: color_data = Z;
		19'b0000110000100101110: color_data = Z;
		19'b0000110000100101111: color_data = Z;
		19'b0000110000100110000: color_data = Z;
		19'b0000110000100110001: color_data = Z;
		19'b0000110000100110010: color_data = Z;
		19'b0000110000100110011: color_data = Z;
		19'b0000110000100110100: color_data = Z;
		19'b0000110000100110101: color_data = Z;
		19'b0000110000100110110: color_data = Z;
		19'b0000110000100110111: color_data = Z;
		19'b0000110000100111000: color_data = Z;
		19'b0000110000100111001: color_data = Z;
		19'b0000110000100111010: color_data = Z;
		19'b0000110000100111011: color_data = Z;
		19'b0000110000100111100: color_data = Z;
		19'b0000110000100111101: color_data = Z;
		19'b0000110000100111110: color_data = Z;
		19'b0000110000100111111: color_data = Z;
		19'b0000110000101000000: color_data = Z;
		19'b0000110000101000001: color_data = Z;
		19'b0000110000101000010: color_data = Z;
		19'b0000110000101000011: color_data = Z;
		19'b0000110000101000100: color_data = Z;
		19'b0000110000101000101: color_data = Z;
		19'b0000110000101000110: color_data = Z;
		19'b0000110000101000111: color_data = Z;
		19'b0000110000101001000: color_data = Z;
		19'b0000110000101001001: color_data = Z;
		19'b0000110000101001010: color_data = Z;
		19'b0000110000101001011: color_data = Z;
		19'b0000110000101001100: color_data = Z;
		19'b0000110000101001101: color_data = Z;
		19'b0000110000101001110: color_data = Z;
		19'b0000110000101001111: color_data = Z;
		19'b0000110000101010000: color_data = Z;
		19'b0000110000101010001: color_data = Z;
		19'b0000110000101010010: color_data = Z;
		19'b0000110000101010011: color_data = Z;
		19'b0000110000101010100: color_data = Z;
		19'b0000110000101010101: color_data = Z;
		19'b0000110000101010110: color_data = Z;
		19'b0000110000101010111: color_data = Z;
		19'b0000110000101011000: color_data = Z;
		19'b0000110000101011001: color_data = Z;
		19'b0000110000101011010: color_data = Z;
		19'b0000110000101011011: color_data = Z;
		19'b0000110000101011100: color_data = Z;
		19'b0000110000101011101: color_data = Z;
		19'b0000110000101011110: color_data = Z;
		19'b0000110000101011111: color_data = Z;
		19'b0000110000101100000: color_data = Z;
		19'b0000110000101100001: color_data = Z;
		19'b0000110000101100010: color_data = Z;
		19'b0000110000101100011: color_data = Z;
		19'b0000110000101100100: color_data = Z;
		19'b0000110000101100101: color_data = Z;
		19'b0000110000101100110: color_data = Z;
		19'b0000110000101100111: color_data = Z;
		19'b0000110000101101000: color_data = Z;
		19'b0000110000101101001: color_data = Z;
		19'b0000110000101101010: color_data = Z;
		19'b0000110000101101011: color_data = Z;
		19'b0000110000101101100: color_data = Z;
		19'b0000110000101101101: color_data = Z;
		19'b0000110000101101110: color_data = Z;
		19'b0000110000101101111: color_data = Z;
		19'b0000110000101110000: color_data = Z;
		19'b0000110000101110001: color_data = Z;
		19'b0000110000101110010: color_data = Z;
		19'b0000110000101110011: color_data = Z;
		19'b0000110000101110100: color_data = Z;
		19'b0000110000101110101: color_data = Z;
		19'b0000110000101110110: color_data = Z;
		19'b0000110000101110111: color_data = Z;
		19'b0000110000101111000: color_data = Z;
		19'b0000110000101111001: color_data = Z;
		19'b0000110000101111010: color_data = Z;
		19'b0000110000101111011: color_data = Z;
		19'b0000110000101111100: color_data = Z;
		19'b0000110000101111101: color_data = Z;
		19'b0000110000101111110: color_data = Z;
		19'b0000110000101111111: color_data = Z;
		19'b0000110000110000000: color_data = Z;
		19'b0000110000110000001: color_data = Z;
		19'b0000110000110000010: color_data = Z;
		19'b0000110000110000011: color_data = Z;
		19'b0000110000110000100: color_data = Z;
		19'b0000110000110000101: color_data = Z;
		19'b0000110000110000110: color_data = Z;
		19'b0000110000110000111: color_data = Z;
		19'b0000110000110001000: color_data = Z;
		19'b0000110000110001001: color_data = Z;
		19'b0000110000110001010: color_data = Z;
		19'b0000110000110001011: color_data = Z;
		19'b0000110000110001100: color_data = Z;
		19'b0000110000110001101: color_data = Z;
		19'b0000110010100000100: color_data = Z;
		19'b0000110010100000101: color_data = Z;
		19'b0000110010100000110: color_data = Z;
		19'b0000110010100000111: color_data = Z;
		19'b0000110010100001000: color_data = Z;
		19'b0000110010100001001: color_data = Z;
		19'b0000110010100001010: color_data = Z;
		19'b0000110010100001011: color_data = Z;
		19'b0000110010100001100: color_data = Z;
		19'b0000110010100001101: color_data = Z;
		19'b0000110010100001110: color_data = Z;
		19'b0000110010100001111: color_data = Z;
		19'b0000110010100010000: color_data = Z;
		19'b0000110010100010001: color_data = Z;
		19'b0000110010100010010: color_data = Z;
		19'b0000110010100010011: color_data = Z;
		19'b0000110010100010100: color_data = Z;
		19'b0000110010100010101: color_data = Z;
		19'b0000110010100010110: color_data = Z;
		19'b0000110010100010111: color_data = Z;
		19'b0000110010100011000: color_data = Z;
		19'b0000110010100011001: color_data = Z;
		19'b0000110010100011010: color_data = Z;
		19'b0000110010100011011: color_data = Z;
		19'b0000110010100011100: color_data = Z;
		19'b0000110010100011101: color_data = Z;
		19'b0000110010100011110: color_data = Z;
		19'b0000110010100011111: color_data = Z;
		19'b0000110010100100000: color_data = Z;
		19'b0000110010100100001: color_data = Z;
		19'b0000110010100100010: color_data = Z;
		19'b0000110010100100011: color_data = Z;
		19'b0000110010100100100: color_data = Z;
		19'b0000110010100100101: color_data = Z;
		19'b0000110010100100110: color_data = Z;
		19'b0000110010100100111: color_data = Z;
		19'b0000110010100101000: color_data = Z;
		19'b0000110010100101001: color_data = Z;
		19'b0000110010100101010: color_data = Z;
		19'b0000110010100101011: color_data = Z;
		19'b0000110010100101100: color_data = Z;
		19'b0000110010100101101: color_data = Z;
		19'b0000110010100101110: color_data = Z;
		19'b0000110010100101111: color_data = Z;
		19'b0000110010100110000: color_data = Z;
		19'b0000110010100110001: color_data = Z;
		19'b0000110010100110010: color_data = Z;
		19'b0000110010100110011: color_data = Z;
		19'b0000110010100110100: color_data = Z;
		19'b0000110010100110101: color_data = Z;
		19'b0000110010100110110: color_data = Z;
		19'b0000110010100110111: color_data = Z;
		19'b0000110010100111000: color_data = Z;
		19'b0000110010100111001: color_data = Z;
		19'b0000110010100111010: color_data = Z;
		19'b0000110010100111011: color_data = Z;
		19'b0000110010100111100: color_data = Z;
		19'b0000110010100111101: color_data = Z;
		19'b0000110010100111110: color_data = Z;
		19'b0000110010100111111: color_data = Z;
		19'b0000110010101000000: color_data = Z;
		19'b0000110010101000001: color_data = Z;
		19'b0000110010101000010: color_data = Z;
		19'b0000110010101000011: color_data = Z;
		19'b0000110010101000100: color_data = Z;
		19'b0000110010101000101: color_data = Z;
		19'b0000110010101000110: color_data = Z;
		19'b0000110010101000111: color_data = Z;
		19'b0000110010101001000: color_data = Z;
		19'b0000110010101001001: color_data = Z;
		19'b0000110010101001010: color_data = Z;
		19'b0000110010101001011: color_data = Z;
		19'b0000110010101001100: color_data = Z;
		19'b0000110010101001101: color_data = Z;
		19'b0000110010101001110: color_data = Z;
		19'b0000110010101001111: color_data = Z;
		19'b0000110010101010000: color_data = Z;
		19'b0000110010101010001: color_data = Z;
		19'b0000110010101010010: color_data = Z;
		19'b0000110010101010011: color_data = Z;
		19'b0000110010101010100: color_data = Z;
		19'b0000110010101010101: color_data = Z;
		19'b0000110010101010110: color_data = Z;
		19'b0000110010101010111: color_data = Z;
		19'b0000110010101011000: color_data = Z;
		19'b0000110010101011001: color_data = Z;
		19'b0000110010101011010: color_data = Z;
		19'b0000110010101011011: color_data = Z;
		19'b0000110010101011100: color_data = Z;
		19'b0000110010101011101: color_data = Z;
		19'b0000110010101011110: color_data = Z;
		19'b0000110010101011111: color_data = Z;
		19'b0000110010101100000: color_data = Z;
		19'b0000110010101100001: color_data = Z;
		19'b0000110010101100010: color_data = Z;
		19'b0000110010101100011: color_data = Z;
		19'b0000110010101100100: color_data = Z;
		19'b0000110010101100101: color_data = Z;
		19'b0000110010101100110: color_data = Z;
		19'b0000110010101100111: color_data = Z;
		19'b0000110010101101000: color_data = Z;
		19'b0000110010101101001: color_data = Z;
		19'b0000110010101101010: color_data = Z;
		19'b0000110010101101011: color_data = Z;
		19'b0000110010101101100: color_data = Z;
		19'b0000110010101101101: color_data = Z;
		19'b0000110010101101110: color_data = Z;
		19'b0000110010101101111: color_data = Z;
		19'b0000110010101110000: color_data = Z;
		19'b0000110010101110001: color_data = Z;
		19'b0000110010101110010: color_data = Z;
		19'b0000110010101110011: color_data = Z;
		19'b0000110010101110100: color_data = Z;
		19'b0000110010101110101: color_data = Z;
		19'b0000110010101110110: color_data = Z;
		19'b0000110010101110111: color_data = Z;
		19'b0000110010101111000: color_data = Z;
		19'b0000110010101111001: color_data = Z;
		19'b0000110010101111010: color_data = Z;
		19'b0000110010101111011: color_data = Z;
		19'b0000110010101111100: color_data = Z;
		19'b0000110010101111101: color_data = Z;
		19'b0000110010101111110: color_data = Z;
		19'b0000110010101111111: color_data = Z;
		19'b0000110010110000000: color_data = Z;
		19'b0000110010110000001: color_data = Z;
		19'b0000110010110000010: color_data = Z;
		19'b0000110010110000011: color_data = Z;
		19'b0000110010110000100: color_data = Z;
		19'b0000110010110000101: color_data = Z;
		19'b0000110010110000110: color_data = Z;
		19'b0000110010110000111: color_data = Z;
		19'b0000110010110001000: color_data = Z;
		19'b0000110010110001001: color_data = Z;
		19'b0000110010110001010: color_data = Z;
		19'b0000110010110001011: color_data = Z;
		19'b0000110010110001100: color_data = Z;
		19'b0000110010110001101: color_data = Z;
		19'b0000110010110001110: color_data = Z;
		19'b0000110100100000010: color_data = Z;
		19'b0000110100100000011: color_data = Z;
		19'b0000110100100000100: color_data = Z;
		19'b0000110100100000101: color_data = Z;
		19'b0000110100100000110: color_data = Z;
		19'b0000110100100000111: color_data = Z;
		19'b0000110100100001000: color_data = Z;
		19'b0000110100100001001: color_data = Z;
		19'b0000110100100001010: color_data = Z;
		19'b0000110100100001011: color_data = Z;
		19'b0000110100100001100: color_data = Z;
		19'b0000110100100001101: color_data = Z;
		19'b0000110100100001110: color_data = Z;
		19'b0000110100100001111: color_data = Z;
		19'b0000110100100010000: color_data = Z;
		19'b0000110100100010001: color_data = Z;
		19'b0000110100100010010: color_data = Z;
		19'b0000110100100010011: color_data = Z;
		19'b0000110100100010100: color_data = Z;
		19'b0000110100100010101: color_data = Z;
		19'b0000110100100010110: color_data = Z;
		19'b0000110100100010111: color_data = Z;
		19'b0000110100100011000: color_data = Z;
		19'b0000110100100011001: color_data = Z;
		19'b0000110100100011010: color_data = Z;
		19'b0000110100100011011: color_data = Z;
		19'b0000110100100011100: color_data = Z;
		19'b0000110100100011101: color_data = Z;
		19'b0000110100100011110: color_data = Z;
		19'b0000110100100011111: color_data = Z;
		19'b0000110100100100000: color_data = Z;
		19'b0000110100100100001: color_data = Z;
		19'b0000110100100100010: color_data = Z;
		19'b0000110100100100011: color_data = Z;
		19'b0000110100100100100: color_data = Z;
		19'b0000110100100100101: color_data = Z;
		19'b0000110100100100110: color_data = Z;
		19'b0000110100100100111: color_data = Z;
		19'b0000110100100101000: color_data = Z;
		19'b0000110100100101001: color_data = Z;
		19'b0000110100100101010: color_data = Z;
		19'b0000110100100101011: color_data = Z;
		19'b0000110100100101100: color_data = Z;
		19'b0000110100100101101: color_data = Z;
		19'b0000110100100101110: color_data = Z;
		19'b0000110100100101111: color_data = Z;
		19'b0000110100100110000: color_data = Z;
		19'b0000110100100110001: color_data = Z;
		19'b0000110100100110010: color_data = Z;
		19'b0000110100100110011: color_data = Z;
		19'b0000110100100110100: color_data = Z;
		19'b0000110100100110101: color_data = Z;
		19'b0000110100100110110: color_data = Z;
		19'b0000110100100110111: color_data = Z;
		19'b0000110100100111000: color_data = Z;
		19'b0000110100100111001: color_data = Z;
		19'b0000110100100111010: color_data = Z;
		19'b0000110100100111011: color_data = Z;
		19'b0000110100100111100: color_data = Z;
		19'b0000110100100111101: color_data = Z;
		19'b0000110100100111110: color_data = Z;
		19'b0000110100100111111: color_data = Z;
		19'b0000110100101000000: color_data = Z;
		19'b0000110100101000001: color_data = Z;
		19'b0000110100101000010: color_data = Z;
		19'b0000110100101000011: color_data = Z;
		19'b0000110100101000100: color_data = Z;
		19'b0000110100101000101: color_data = Z;
		19'b0000110100101000110: color_data = Z;
		19'b0000110100101000111: color_data = Z;
		19'b0000110100101001000: color_data = Z;
		19'b0000110100101001001: color_data = Z;
		19'b0000110100101001010: color_data = Z;
		19'b0000110100101001011: color_data = Z;
		19'b0000110100101001100: color_data = Z;
		19'b0000110100101001101: color_data = Z;
		19'b0000110100101001110: color_data = Z;
		19'b0000110100101001111: color_data = Z;
		19'b0000110100101010000: color_data = Z;
		19'b0000110100101010001: color_data = Z;
		19'b0000110100101010010: color_data = Z;
		19'b0000110100101010011: color_data = Z;
		19'b0000110100101010100: color_data = Z;
		19'b0000110100101010101: color_data = Z;
		19'b0000110100101010110: color_data = Z;
		19'b0000110100101010111: color_data = Z;
		19'b0000110100101011000: color_data = Z;
		19'b0000110100101011001: color_data = Z;
		19'b0000110100101011010: color_data = Z;
		19'b0000110100101011011: color_data = Z;
		19'b0000110100101011100: color_data = Z;
		19'b0000110100101011101: color_data = Z;
		19'b0000110100101011110: color_data = Z;
		19'b0000110100101011111: color_data = Z;
		19'b0000110100101100000: color_data = Z;
		19'b0000110100101100001: color_data = Z;
		19'b0000110100101100010: color_data = Z;
		19'b0000110100101100011: color_data = Z;
		19'b0000110100101100100: color_data = Z;
		19'b0000110100101100101: color_data = Z;
		19'b0000110100101100110: color_data = Z;
		19'b0000110100101100111: color_data = Z;
		19'b0000110100101101000: color_data = Z;
		19'b0000110100101101001: color_data = Z;
		19'b0000110100101101010: color_data = Z;
		19'b0000110100101101011: color_data = Z;
		19'b0000110100101101100: color_data = Z;
		19'b0000110100101101101: color_data = Z;
		19'b0000110100101101110: color_data = Z;
		19'b0000110100101101111: color_data = Z;
		19'b0000110100101110000: color_data = Z;
		19'b0000110100101110001: color_data = Z;
		19'b0000110100101110010: color_data = Z;
		19'b0000110100101110011: color_data = Z;
		19'b0000110100101110100: color_data = Z;
		19'b0000110100101110101: color_data = Z;
		19'b0000110100101110110: color_data = Z;
		19'b0000110100101110111: color_data = Z;
		19'b0000110100101111000: color_data = Z;
		19'b0000110100101111001: color_data = Z;
		19'b0000110100101111010: color_data = Z;
		19'b0000110100101111011: color_data = Z;
		19'b0000110100101111100: color_data = Z;
		19'b0000110100101111101: color_data = Z;
		19'b0000110100101111110: color_data = Z;
		19'b0000110100101111111: color_data = Z;
		19'b0000110100110000000: color_data = Z;
		19'b0000110100110000001: color_data = Z;
		19'b0000110100110000010: color_data = Z;
		19'b0000110100110000011: color_data = Z;
		19'b0000110100110000100: color_data = Z;
		19'b0000110100110000101: color_data = Z;
		19'b0000110100110000110: color_data = Z;
		19'b0000110100110000111: color_data = Z;
		19'b0000110100110001000: color_data = Z;
		19'b0000110100110001001: color_data = Z;
		19'b0000110100110001010: color_data = Z;
		19'b0000110100110001011: color_data = Z;
		19'b0000110100110001100: color_data = Z;
		19'b0000110100110001101: color_data = Z;
		19'b0000110100110001110: color_data = Z;
		19'b0000110100110001111: color_data = Z;
		19'b0000110110011111000: color_data = Z;
		19'b0000110110011111001: color_data = Z;
		19'b0000110110100000000: color_data = Z;
		19'b0000110110100000001: color_data = Z;
		19'b0000110110100000010: color_data = Z;
		19'b0000110110100000011: color_data = Z;
		19'b0000110110100000100: color_data = Z;
		19'b0000110110100000101: color_data = Z;
		19'b0000110110100000110: color_data = Z;
		19'b0000110110100000111: color_data = Z;
		19'b0000110110100001000: color_data = Z;
		19'b0000110110100001001: color_data = Z;
		19'b0000110110100001010: color_data = Z;
		19'b0000110110100001011: color_data = Z;
		19'b0000110110100001100: color_data = Z;
		19'b0000110110100001101: color_data = Z;
		19'b0000110110100001110: color_data = Z;
		19'b0000110110100001111: color_data = Z;
		19'b0000110110100010000: color_data = Z;
		19'b0000110110100010001: color_data = Z;
		19'b0000110110100010010: color_data = Z;
		19'b0000110110100010011: color_data = Z;
		19'b0000110110100010100: color_data = Z;
		19'b0000110110100010101: color_data = Z;
		19'b0000110110100010110: color_data = Z;
		19'b0000110110100010111: color_data = Z;
		19'b0000110110100011000: color_data = Z;
		19'b0000110110100011001: color_data = Z;
		19'b0000110110100011010: color_data = Z;
		19'b0000110110100011011: color_data = Z;
		19'b0000110110100011100: color_data = Z;
		19'b0000110110100011101: color_data = Z;
		19'b0000110110100011110: color_data = Z;
		19'b0000110110100011111: color_data = Z;
		19'b0000110110100100000: color_data = Z;
		19'b0000110110100100001: color_data = Z;
		19'b0000110110100100010: color_data = Z;
		19'b0000110110100100011: color_data = Z;
		19'b0000110110100100100: color_data = Z;
		19'b0000110110100100101: color_data = Z;
		19'b0000110110100100110: color_data = Z;
		19'b0000110110100100111: color_data = Z;
		19'b0000110110100101000: color_data = Z;
		19'b0000110110100101001: color_data = Z;
		19'b0000110110100101010: color_data = Z;
		19'b0000110110100101011: color_data = Z;
		19'b0000110110100101100: color_data = Z;
		19'b0000110110100101101: color_data = Z;
		19'b0000110110100101110: color_data = Z;
		19'b0000110110100101111: color_data = Z;
		19'b0000110110100110000: color_data = Z;
		19'b0000110110100110001: color_data = Z;
		19'b0000110110100110010: color_data = Z;
		19'b0000110110100110011: color_data = Z;
		19'b0000110110100110100: color_data = Z;
		19'b0000110110100110101: color_data = Z;
		19'b0000110110100110110: color_data = Z;
		19'b0000110110100110111: color_data = Z;
		19'b0000110110100111000: color_data = Z;
		19'b0000110110100111001: color_data = Z;
		19'b0000110110100111010: color_data = Z;
		19'b0000110110100111011: color_data = Z;
		19'b0000110110100111100: color_data = Z;
		19'b0000110110100111101: color_data = Z;
		19'b0000110110100111110: color_data = Z;
		19'b0000110110100111111: color_data = Z;
		19'b0000110110101000000: color_data = Z;
		19'b0000110110101000001: color_data = Z;
		19'b0000110110101000010: color_data = Z;
		19'b0000110110101000011: color_data = Z;
		19'b0000110110101000100: color_data = Z;
		19'b0000110110101000101: color_data = Z;
		19'b0000110110101000110: color_data = Z;
		19'b0000110110101000111: color_data = Z;
		19'b0000110110101001000: color_data = Z;
		19'b0000110110101001001: color_data = Z;
		19'b0000110110101001010: color_data = Z;
		19'b0000110110101001011: color_data = Z;
		19'b0000110110101001100: color_data = Z;
		19'b0000110110101001101: color_data = Z;
		19'b0000110110101001110: color_data = Z;
		19'b0000110110101001111: color_data = Z;
		19'b0000110110101010000: color_data = Z;
		19'b0000110110101010001: color_data = Z;
		19'b0000110110101010010: color_data = Z;
		19'b0000110110101010011: color_data = Z;
		19'b0000110110101010100: color_data = Z;
		19'b0000110110101010101: color_data = Z;
		19'b0000110110101010110: color_data = Z;
		19'b0000110110101010111: color_data = Z;
		19'b0000110110101011000: color_data = Z;
		19'b0000110110101011001: color_data = Z;
		19'b0000110110101011010: color_data = Z;
		19'b0000110110101011011: color_data = Z;
		19'b0000110110101011100: color_data = Z;
		19'b0000110110101011101: color_data = Z;
		19'b0000110110101011110: color_data = Z;
		19'b0000110110101011111: color_data = Z;
		19'b0000110110101100000: color_data = Z;
		19'b0000110110101100001: color_data = Z;
		19'b0000110110101100010: color_data = Z;
		19'b0000110110101100011: color_data = Z;
		19'b0000110110101100100: color_data = Z;
		19'b0000110110101100101: color_data = Z;
		19'b0000110110101100110: color_data = Z;
		19'b0000110110101100111: color_data = Z;
		19'b0000110110101101000: color_data = Z;
		19'b0000110110101101001: color_data = Z;
		19'b0000110110101101010: color_data = Z;
		19'b0000110110101101011: color_data = Z;
		19'b0000110110101101100: color_data = Z;
		19'b0000110110101101101: color_data = Z;
		19'b0000110110101101110: color_data = Z;
		19'b0000110110101101111: color_data = Z;
		19'b0000110110101110000: color_data = Z;
		19'b0000110110101110001: color_data = Z;
		19'b0000110110101110010: color_data = Z;
		19'b0000110110101110011: color_data = Z;
		19'b0000110110101110100: color_data = Z;
		19'b0000110110101110101: color_data = Z;
		19'b0000110110101110110: color_data = Z;
		19'b0000110110101110111: color_data = Z;
		19'b0000110110101111000: color_data = Z;
		19'b0000110110101111001: color_data = Z;
		19'b0000110110101111010: color_data = Z;
		19'b0000110110101111011: color_data = Z;
		19'b0000110110101111100: color_data = Z;
		19'b0000110110101111101: color_data = Z;
		19'b0000110110101111110: color_data = Z;
		19'b0000110110101111111: color_data = Z;
		19'b0000110110110000000: color_data = Z;
		19'b0000110110110000001: color_data = Z;
		19'b0000110110110000010: color_data = Z;
		19'b0000110110110000011: color_data = Z;
		19'b0000110110110000100: color_data = Z;
		19'b0000110110110000101: color_data = Z;
		19'b0000110110110000110: color_data = Z;
		19'b0000110110110000111: color_data = Z;
		19'b0000110110110001000: color_data = Z;
		19'b0000110110110001001: color_data = Z;
		19'b0000110110110001010: color_data = Z;
		19'b0000110110110001011: color_data = Z;
		19'b0000110110110001100: color_data = Z;
		19'b0000110110110001101: color_data = Z;
		19'b0000110110110001110: color_data = Z;
		19'b0000110110110001111: color_data = Z;
		19'b0000110110110010000: color_data = Z;
		19'b0000111000011110110: color_data = Z;
		19'b0000111000011110111: color_data = Z;
		19'b0000111000011111000: color_data = Z;
		19'b0000111000011111110: color_data = Z;
		19'b0000111000011111111: color_data = Z;
		19'b0000111000100000000: color_data = Z;
		19'b0000111000100000001: color_data = Z;
		19'b0000111000100000010: color_data = Z;
		19'b0000111000100000011: color_data = Z;
		19'b0000111000100000100: color_data = Z;
		19'b0000111000100000101: color_data = Z;
		19'b0000111000100000110: color_data = Z;
		19'b0000111000100000111: color_data = Z;
		19'b0000111000100001000: color_data = Z;
		19'b0000111000100001001: color_data = Z;
		19'b0000111000100001010: color_data = Z;
		19'b0000111000100001011: color_data = Z;
		19'b0000111000100001100: color_data = Z;
		19'b0000111000100001101: color_data = Z;
		19'b0000111000100001110: color_data = Z;
		19'b0000111000100001111: color_data = Z;
		19'b0000111000100010000: color_data = Z;
		19'b0000111000100010001: color_data = Z;
		19'b0000111000100010010: color_data = Z;
		19'b0000111000100010011: color_data = Z;
		19'b0000111000100010100: color_data = Z;
		19'b0000111000100010101: color_data = Z;
		19'b0000111000100010110: color_data = Z;
		19'b0000111000100010111: color_data = Z;
		19'b0000111000100011000: color_data = Z;
		19'b0000111000100011001: color_data = Z;
		19'b0000111000100011010: color_data = Z;
		19'b0000111000100011011: color_data = Z;
		19'b0000111000100011100: color_data = Z;
		19'b0000111000100011101: color_data = Z;
		19'b0000111000100011110: color_data = Z;
		19'b0000111000100011111: color_data = Z;
		19'b0000111000100100000: color_data = Z;
		19'b0000111000100100001: color_data = Z;
		19'b0000111000100100010: color_data = Z;
		19'b0000111000100100011: color_data = Z;
		19'b0000111000100100100: color_data = Z;
		19'b0000111000100100101: color_data = Z;
		19'b0000111000100100110: color_data = Z;
		19'b0000111000100100111: color_data = Z;
		19'b0000111000100101000: color_data = Z;
		19'b0000111000100101001: color_data = Z;
		19'b0000111000100101010: color_data = Z;
		19'b0000111000100101011: color_data = Z;
		19'b0000111000100101100: color_data = Z;
		19'b0000111000100101101: color_data = Z;
		19'b0000111000100101110: color_data = Z;
		19'b0000111000100101111: color_data = Z;
		19'b0000111000100110000: color_data = Z;
		19'b0000111000100110001: color_data = Z;
		19'b0000111000100110010: color_data = Z;
		19'b0000111000100110011: color_data = Z;
		19'b0000111000100110100: color_data = Z;
		19'b0000111000100110101: color_data = Z;
		19'b0000111000100110110: color_data = Z;
		19'b0000111000100110111: color_data = Z;
		19'b0000111000100111000: color_data = Z;
		19'b0000111000100111001: color_data = Z;
		19'b0000111000100111010: color_data = Z;
		19'b0000111000100111011: color_data = Z;
		19'b0000111000100111100: color_data = Z;
		19'b0000111000100111101: color_data = Z;
		19'b0000111000100111110: color_data = Z;
		19'b0000111000100111111: color_data = Z;
		19'b0000111000101000000: color_data = Z;
		19'b0000111000101000001: color_data = Z;
		19'b0000111000101000010: color_data = Z;
		19'b0000111000101000011: color_data = Z;
		19'b0000111000101000100: color_data = Z;
		19'b0000111000101000101: color_data = Z;
		19'b0000111000101000110: color_data = Z;
		19'b0000111000101000111: color_data = Z;
		19'b0000111000101001000: color_data = Z;
		19'b0000111000101001001: color_data = Z;
		19'b0000111000101001010: color_data = Z;
		19'b0000111000101001011: color_data = Z;
		19'b0000111000101001100: color_data = Z;
		19'b0000111000101001101: color_data = Z;
		19'b0000111000101001110: color_data = Z;
		19'b0000111000101001111: color_data = Z;
		19'b0000111000101010000: color_data = Z;
		19'b0000111000101010001: color_data = Z;
		19'b0000111000101010010: color_data = Z;
		19'b0000111000101010011: color_data = Z;
		19'b0000111000101010100: color_data = Z;
		19'b0000111000101010101: color_data = Z;
		19'b0000111000101010110: color_data = Z;
		19'b0000111000101010111: color_data = Z;
		19'b0000111000101011000: color_data = Z;
		19'b0000111000101011001: color_data = Z;
		19'b0000111000101011010: color_data = Z;
		19'b0000111000101011011: color_data = Z;
		19'b0000111000101011100: color_data = Z;
		19'b0000111000101011101: color_data = Z;
		19'b0000111000101011110: color_data = Z;
		19'b0000111000101011111: color_data = Z;
		19'b0000111000101100000: color_data = Z;
		19'b0000111000101100001: color_data = Z;
		19'b0000111000101100010: color_data = Z;
		19'b0000111000101100011: color_data = Z;
		19'b0000111000101100100: color_data = Z;
		19'b0000111000101100101: color_data = Z;
		19'b0000111000101100110: color_data = Z;
		19'b0000111000101100111: color_data = Z;
		19'b0000111000101101000: color_data = Z;
		19'b0000111000101101001: color_data = Z;
		19'b0000111000101101010: color_data = Z;
		19'b0000111000101101011: color_data = Z;
		19'b0000111000101101100: color_data = Z;
		19'b0000111000101101101: color_data = Z;
		19'b0000111000101101110: color_data = Z;
		19'b0000111000101101111: color_data = Z;
		19'b0000111000101110000: color_data = Z;
		19'b0000111000101110001: color_data = Z;
		19'b0000111000101110010: color_data = Z;
		19'b0000111000101110011: color_data = Z;
		19'b0000111000101110100: color_data = Z;
		19'b0000111000101110101: color_data = Z;
		19'b0000111000101110110: color_data = Z;
		19'b0000111000101110111: color_data = Z;
		19'b0000111000101111000: color_data = Z;
		19'b0000111000101111001: color_data = Z;
		19'b0000111000101111010: color_data = Z;
		19'b0000111000101111011: color_data = Z;
		19'b0000111000101111100: color_data = Z;
		19'b0000111000101111101: color_data = Z;
		19'b0000111000101111110: color_data = Z;
		19'b0000111000101111111: color_data = Z;
		19'b0000111000110000000: color_data = Z;
		19'b0000111000110000001: color_data = Z;
		19'b0000111000110000010: color_data = Z;
		19'b0000111000110000011: color_data = Z;
		19'b0000111000110000100: color_data = Z;
		19'b0000111000110000101: color_data = Z;
		19'b0000111000110000110: color_data = Z;
		19'b0000111000110000111: color_data = Z;
		19'b0000111000110001000: color_data = Z;
		19'b0000111000110001001: color_data = Z;
		19'b0000111000110001010: color_data = Z;
		19'b0000111000110001011: color_data = Z;
		19'b0000111000110001100: color_data = Z;
		19'b0000111000110001101: color_data = Z;
		19'b0000111000110001110: color_data = Z;
		19'b0000111000110001111: color_data = Z;
		19'b0000111000110010000: color_data = Z;
		19'b0000111000110010001: color_data = Z;
		19'b0000111010011110100: color_data = Z;
		19'b0000111010011110101: color_data = Z;
		19'b0000111010011110110: color_data = Z;
		19'b0000111010011110111: color_data = Z;
		19'b0000111010011111100: color_data = Z;
		19'b0000111010011111101: color_data = Z;
		19'b0000111010011111110: color_data = Z;
		19'b0000111010011111111: color_data = Z;
		19'b0000111010100000000: color_data = Z;
		19'b0000111010100000001: color_data = Z;
		19'b0000111010100000010: color_data = Z;
		19'b0000111010100000011: color_data = Z;
		19'b0000111010100000100: color_data = Z;
		19'b0000111010100000101: color_data = Z;
		19'b0000111010100000110: color_data = Z;
		19'b0000111010100000111: color_data = Z;
		19'b0000111010100001000: color_data = Z;
		19'b0000111010100001001: color_data = Z;
		19'b0000111010100001010: color_data = Z;
		19'b0000111010100001011: color_data = Z;
		19'b0000111010100001100: color_data = Z;
		19'b0000111010100001101: color_data = Z;
		19'b0000111010100001110: color_data = Z;
		19'b0000111010100001111: color_data = Z;
		19'b0000111010100010000: color_data = Z;
		19'b0000111010100010001: color_data = Z;
		19'b0000111010100010010: color_data = Z;
		19'b0000111010100010011: color_data = Z;
		19'b0000111010100010100: color_data = Z;
		19'b0000111010100010101: color_data = Z;
		19'b0000111010100010110: color_data = Z;
		19'b0000111010100010111: color_data = Z;
		19'b0000111010100011000: color_data = Z;
		19'b0000111010100011001: color_data = Z;
		19'b0000111010100011010: color_data = Z;
		19'b0000111010100011011: color_data = Z;
		19'b0000111010100011100: color_data = Z;
		19'b0000111010100011101: color_data = Z;
		19'b0000111010100011110: color_data = Z;
		19'b0000111010100011111: color_data = Z;
		19'b0000111010100100000: color_data = Z;
		19'b0000111010100100001: color_data = Z;
		19'b0000111010100100010: color_data = Z;
		19'b0000111010100100011: color_data = Z;
		19'b0000111010100100100: color_data = Z;
		19'b0000111010100100101: color_data = Z;
		19'b0000111010100100110: color_data = Z;
		19'b0000111010100100111: color_data = Z;
		19'b0000111010100101000: color_data = Z;
		19'b0000111010100101001: color_data = Z;
		19'b0000111010100101010: color_data = Z;
		19'b0000111010100101011: color_data = Z;
		19'b0000111010100101100: color_data = Z;
		19'b0000111010100101101: color_data = Z;
		19'b0000111010100101110: color_data = Z;
		19'b0000111010100101111: color_data = Z;
		19'b0000111010100110000: color_data = Z;
		19'b0000111010100110001: color_data = Z;
		19'b0000111010100110010: color_data = Z;
		19'b0000111010100110011: color_data = Z;
		19'b0000111010100110100: color_data = Z;
		19'b0000111010100110101: color_data = Z;
		19'b0000111010100110110: color_data = Z;
		19'b0000111010100110111: color_data = Z;
		19'b0000111010100111000: color_data = Z;
		19'b0000111010100111001: color_data = Z;
		19'b0000111010100111010: color_data = Z;
		19'b0000111010100111011: color_data = Z;
		19'b0000111010100111100: color_data = Z;
		19'b0000111010100111101: color_data = Z;
		19'b0000111010100111110: color_data = Z;
		19'b0000111010100111111: color_data = Z;
		19'b0000111010101000000: color_data = Z;
		19'b0000111010101000001: color_data = Z;
		19'b0000111010101000010: color_data = Z;
		19'b0000111010101000011: color_data = Z;
		19'b0000111010101000100: color_data = Z;
		19'b0000111010101000101: color_data = Z;
		19'b0000111010101000110: color_data = Z;
		19'b0000111010101000111: color_data = Z;
		19'b0000111010101001000: color_data = Z;
		19'b0000111010101001001: color_data = Z;
		19'b0000111010101001010: color_data = Z;
		19'b0000111010101001011: color_data = Z;
		19'b0000111010101001100: color_data = Z;
		19'b0000111010101001101: color_data = Z;
		19'b0000111010101001110: color_data = Z;
		19'b0000111010101001111: color_data = Z;
		19'b0000111010101010000: color_data = Z;
		19'b0000111010101010001: color_data = Z;
		19'b0000111010101010010: color_data = Z;
		19'b0000111010101010011: color_data = Z;
		19'b0000111010101010100: color_data = Z;
		19'b0000111010101010101: color_data = Z;
		19'b0000111010101010110: color_data = Z;
		19'b0000111010101010111: color_data = Z;
		19'b0000111010101011000: color_data = Z;
		19'b0000111010101011001: color_data = Z;
		19'b0000111010101011010: color_data = Z;
		19'b0000111010101011011: color_data = Z;
		19'b0000111010101011100: color_data = Z;
		19'b0000111010101011101: color_data = Z;
		19'b0000111010101011110: color_data = Z;
		19'b0000111010101011111: color_data = Z;
		19'b0000111010101100000: color_data = Z;
		19'b0000111010101100001: color_data = Z;
		19'b0000111010101100010: color_data = Z;
		19'b0000111010101100011: color_data = Z;
		19'b0000111010101100100: color_data = Z;
		19'b0000111010101100101: color_data = Z;
		19'b0000111010101100110: color_data = Z;
		19'b0000111010101100111: color_data = Z;
		19'b0000111010101101000: color_data = Z;
		19'b0000111010101101001: color_data = Z;
		19'b0000111010101101010: color_data = Z;
		19'b0000111010101101011: color_data = Z;
		19'b0000111010101101100: color_data = Z;
		19'b0000111010101101101: color_data = Z;
		19'b0000111010101101110: color_data = Z;
		19'b0000111010101101111: color_data = Z;
		19'b0000111010101110000: color_data = Z;
		19'b0000111010101110001: color_data = Z;
		19'b0000111010101110010: color_data = Z;
		19'b0000111010101110011: color_data = Z;
		19'b0000111010101110100: color_data = Z;
		19'b0000111010101110101: color_data = Z;
		19'b0000111010101110110: color_data = Z;
		19'b0000111010101110111: color_data = Z;
		19'b0000111010101111000: color_data = Z;
		19'b0000111010101111001: color_data = Z;
		19'b0000111010101111010: color_data = Z;
		19'b0000111010101111011: color_data = Z;
		19'b0000111010101111100: color_data = Z;
		19'b0000111010101111101: color_data = Z;
		19'b0000111010101111110: color_data = Z;
		19'b0000111010101111111: color_data = Z;
		19'b0000111010110000000: color_data = Z;
		19'b0000111010110000001: color_data = Z;
		19'b0000111010110000010: color_data = Z;
		19'b0000111010110000011: color_data = Z;
		19'b0000111010110000100: color_data = Z;
		19'b0000111010110000101: color_data = Z;
		19'b0000111010110000110: color_data = Z;
		19'b0000111010110000111: color_data = Z;
		19'b0000111010110001000: color_data = Z;
		19'b0000111010110001001: color_data = Z;
		19'b0000111010110001010: color_data = Z;
		19'b0000111010110001011: color_data = Z;
		19'b0000111010110001100: color_data = Z;
		19'b0000111010110001101: color_data = Z;
		19'b0000111010110001110: color_data = Z;
		19'b0000111010110001111: color_data = Z;
		19'b0000111010110010000: color_data = Z;
		19'b0000111010110010001: color_data = Z;
		19'b0000111010110010010: color_data = Z;
		19'b0000111010110010011: color_data = Z;
		19'b0000111100011110010: color_data = Z;
		19'b0000111100011110011: color_data = Z;
		19'b0000111100011110100: color_data = Z;
		19'b0000111100011110101: color_data = Z;
		19'b0000111100011110110: color_data = Z;
		19'b0000111100011111010: color_data = Z;
		19'b0000111100011111011: color_data = Z;
		19'b0000111100011111100: color_data = Z;
		19'b0000111100011111101: color_data = Z;
		19'b0000111100011111110: color_data = Z;
		19'b0000111100011111111: color_data = Z;
		19'b0000111100100000000: color_data = Z;
		19'b0000111100100000001: color_data = Z;
		19'b0000111100100000010: color_data = Z;
		19'b0000111100100000011: color_data = Z;
		19'b0000111100100000100: color_data = Z;
		19'b0000111100100000101: color_data = Z;
		19'b0000111100100000110: color_data = Z;
		19'b0000111100100000111: color_data = Z;
		19'b0000111100100001000: color_data = Z;
		19'b0000111100100001001: color_data = Z;
		19'b0000111100100001010: color_data = Z;
		19'b0000111100100001011: color_data = Z;
		19'b0000111100100001100: color_data = Z;
		19'b0000111100100001101: color_data = Z;
		19'b0000111100100001110: color_data = Z;
		19'b0000111100100001111: color_data = Z;
		19'b0000111100100010000: color_data = Z;
		19'b0000111100100010001: color_data = Z;
		19'b0000111100100010010: color_data = Z;
		19'b0000111100100010011: color_data = Z;
		19'b0000111100100010100: color_data = Z;
		19'b0000111100100010101: color_data = Z;
		19'b0000111100100010110: color_data = Z;
		19'b0000111100100010111: color_data = Z;
		19'b0000111100100011000: color_data = Z;
		19'b0000111100100011001: color_data = Z;
		19'b0000111100100011010: color_data = Z;
		19'b0000111100100011011: color_data = Z;
		19'b0000111100100011100: color_data = Z;
		19'b0000111100100011101: color_data = Z;
		19'b0000111100100011110: color_data = Z;
		19'b0000111100100011111: color_data = Z;
		19'b0000111100100100000: color_data = Z;
		19'b0000111100100100001: color_data = Z;
		19'b0000111100100100010: color_data = Z;
		19'b0000111100100100011: color_data = Z;
		19'b0000111100100100100: color_data = Z;
		19'b0000111100100100101: color_data = Z;
		19'b0000111100100100110: color_data = Z;
		19'b0000111100100100111: color_data = Z;
		19'b0000111100100101000: color_data = Z;
		19'b0000111100100101001: color_data = Z;
		19'b0000111100100101010: color_data = Z;
		19'b0000111100100101011: color_data = Z;
		19'b0000111100100101100: color_data = Z;
		19'b0000111100100101101: color_data = Z;
		19'b0000111100100101110: color_data = Z;
		19'b0000111100100101111: color_data = Z;
		19'b0000111100100110000: color_data = Z;
		19'b0000111100100110001: color_data = Z;
		19'b0000111100100110010: color_data = Z;
		19'b0000111100100110011: color_data = Z;
		19'b0000111100100110100: color_data = Z;
		19'b0000111100100110101: color_data = Z;
		19'b0000111100100110110: color_data = Z;
		19'b0000111100100110111: color_data = Z;
		19'b0000111100100111000: color_data = Z;
		19'b0000111100100111001: color_data = Z;
		19'b0000111100100111010: color_data = Z;
		19'b0000111100100111011: color_data = Z;
		19'b0000111100100111100: color_data = Z;
		19'b0000111100100111101: color_data = Z;
		19'b0000111100100111110: color_data = Z;
		19'b0000111100100111111: color_data = Z;
		19'b0000111100101000000: color_data = Z;
		19'b0000111100101000001: color_data = Z;
		19'b0000111100101000010: color_data = Z;
		19'b0000111100101000011: color_data = Z;
		19'b0000111100101000100: color_data = Z;
		19'b0000111100101000101: color_data = Z;
		19'b0000111100101000110: color_data = Z;
		19'b0000111100101000111: color_data = Z;
		19'b0000111100101001000: color_data = Z;
		19'b0000111100101001001: color_data = Z;
		19'b0000111100101001010: color_data = Z;
		19'b0000111100101001011: color_data = Z;
		19'b0000111100101001100: color_data = Z;
		19'b0000111100101001101: color_data = Z;
		19'b0000111100101001110: color_data = Z;
		19'b0000111100101001111: color_data = Z;
		19'b0000111100101010000: color_data = Z;
		19'b0000111100101010001: color_data = Z;
		19'b0000111100101010010: color_data = Z;
		19'b0000111100101010011: color_data = Z;
		19'b0000111100101010100: color_data = Z;
		19'b0000111100101010101: color_data = Z;
		19'b0000111100101010110: color_data = Z;
		19'b0000111100101010111: color_data = Z;
		19'b0000111100101011000: color_data = Z;
		19'b0000111100101011001: color_data = Z;
		19'b0000111100101011010: color_data = Z;
		19'b0000111100101011011: color_data = Z;
		19'b0000111100101011100: color_data = Z;
		19'b0000111100101011101: color_data = Z;
		19'b0000111100101011110: color_data = Z;
		19'b0000111100101011111: color_data = Z;
		19'b0000111100101100000: color_data = Z;
		19'b0000111100101100001: color_data = Z;
		19'b0000111100101100010: color_data = Z;
		19'b0000111100101100011: color_data = Z;
		19'b0000111100101100100: color_data = Z;
		19'b0000111100101100101: color_data = Z;
		19'b0000111100101100110: color_data = Z;
		19'b0000111100101100111: color_data = Z;
		19'b0000111100101101000: color_data = Z;
		19'b0000111100101101001: color_data = Z;
		19'b0000111100101101010: color_data = Z;
		19'b0000111100101101011: color_data = Z;
		19'b0000111100101101100: color_data = Z;
		19'b0000111100101101101: color_data = Z;
		19'b0000111100101101110: color_data = Z;
		19'b0000111100101101111: color_data = Z;
		19'b0000111100101110000: color_data = Z;
		19'b0000111100101110001: color_data = Z;
		19'b0000111100101110010: color_data = Z;
		19'b0000111100101110011: color_data = Z;
		19'b0000111100101110100: color_data = Z;
		19'b0000111100101110101: color_data = Z;
		19'b0000111100101110110: color_data = Z;
		19'b0000111100101110111: color_data = Z;
		19'b0000111100101111000: color_data = Z;
		19'b0000111100101111001: color_data = Z;
		19'b0000111100101111010: color_data = Z;
		19'b0000111100101111011: color_data = Z;
		19'b0000111100101111100: color_data = Z;
		19'b0000111100101111101: color_data = Z;
		19'b0000111100101111110: color_data = Z;
		19'b0000111100101111111: color_data = Z;
		19'b0000111100110000000: color_data = Z;
		19'b0000111100110000001: color_data = Z;
		19'b0000111100110000010: color_data = Z;
		19'b0000111100110000011: color_data = Z;
		19'b0000111100110000100: color_data = Z;
		19'b0000111100110000101: color_data = Z;
		19'b0000111100110000110: color_data = Z;
		19'b0000111100110000111: color_data = Z;
		19'b0000111100110001000: color_data = Z;
		19'b0000111100110001001: color_data = Z;
		19'b0000111100110001010: color_data = Z;
		19'b0000111100110001011: color_data = Z;
		19'b0000111100110001100: color_data = Z;
		19'b0000111100110001101: color_data = Z;
		19'b0000111100110001110: color_data = Z;
		19'b0000111100110001111: color_data = Z;
		19'b0000111100110010000: color_data = Z;
		19'b0000111100110010001: color_data = Z;
		19'b0000111100110010010: color_data = Z;
		19'b0000111100110010011: color_data = Z;
		19'b0000111100110010100: color_data = Z;
		19'b0000111100110010101: color_data = Z;
		19'b0000111100110010110: color_data = Z;
		19'b0000111110011110001: color_data = Z;
		19'b0000111110011110010: color_data = Z;
		19'b0000111110011110011: color_data = Z;
		19'b0000111110011110100: color_data = Z;
		19'b0000111110011110101: color_data = Z;
		19'b0000111110011110110: color_data = Z;
		19'b0000111110011110111: color_data = Z;
		19'b0000111110011111000: color_data = Z;
		19'b0000111110011111001: color_data = Z;
		19'b0000111110011111010: color_data = Z;
		19'b0000111110011111011: color_data = Z;
		19'b0000111110011111100: color_data = Z;
		19'b0000111110011111101: color_data = Z;
		19'b0000111110011111110: color_data = Z;
		19'b0000111110011111111: color_data = Z;
		19'b0000111110100000000: color_data = Z;
		19'b0000111110100000001: color_data = Z;
		19'b0000111110100000010: color_data = Z;
		19'b0000111110100000011: color_data = Z;
		19'b0000111110100000100: color_data = Z;
		19'b0000111110100000101: color_data = Z;
		19'b0000111110100000110: color_data = Z;
		19'b0000111110100000111: color_data = Z;
		19'b0000111110100001000: color_data = Z;
		19'b0000111110100001001: color_data = Z;
		19'b0000111110100001010: color_data = Z;
		19'b0000111110100001011: color_data = Z;
		19'b0000111110100001100: color_data = Z;
		19'b0000111110100001101: color_data = Z;
		19'b0000111110100001110: color_data = Z;
		19'b0000111110100001111: color_data = Z;
		19'b0000111110100010000: color_data = Z;
		19'b0000111110100010001: color_data = Z;
		19'b0000111110100010010: color_data = Z;
		19'b0000111110100010011: color_data = Z;
		19'b0000111110100010100: color_data = Z;
		19'b0000111110100010101: color_data = Z;
		19'b0000111110100010110: color_data = Z;
		19'b0000111110100010111: color_data = Z;
		19'b0000111110100011000: color_data = Z;
		19'b0000111110100011001: color_data = Z;
		19'b0000111110100011010: color_data = Z;
		19'b0000111110100011011: color_data = Z;
		19'b0000111110100011100: color_data = Z;
		19'b0000111110100011101: color_data = Z;
		19'b0000111110100011110: color_data = Z;
		19'b0000111110100011111: color_data = Z;
		19'b0000111110100100000: color_data = Z;
		19'b0000111110100100001: color_data = Z;
		19'b0000111110100100010: color_data = Z;
		19'b0000111110100100011: color_data = Z;
		19'b0000111110100100100: color_data = Z;
		19'b0000111110100100101: color_data = Z;
		19'b0000111110100100110: color_data = Z;
		19'b0000111110100100111: color_data = Z;
		19'b0000111110100101000: color_data = Z;
		19'b0000111110100101001: color_data = Z;
		19'b0000111110100101010: color_data = Z;
		19'b0000111110100101011: color_data = Z;
		19'b0000111110100101100: color_data = Z;
		19'b0000111110100101101: color_data = Z;
		19'b0000111110100101110: color_data = Z;
		19'b0000111110100101111: color_data = Z;
		19'b0000111110100110000: color_data = Z;
		19'b0000111110100110001: color_data = Z;
		19'b0000111110100110010: color_data = Z;
		19'b0000111110100110011: color_data = Z;
		19'b0000111110100110100: color_data = Z;
		19'b0000111110100110101: color_data = Z;
		19'b0000111110100110110: color_data = Z;
		19'b0000111110100110111: color_data = Z;
		19'b0000111110100111000: color_data = Z;
		19'b0000111110100111001: color_data = Z;
		19'b0000111110100111010: color_data = Z;
		19'b0000111110100111011: color_data = Z;
		19'b0000111110100111100: color_data = Z;
		19'b0000111110100111101: color_data = Z;
		19'b0000111110100111110: color_data = Z;
		19'b0000111110100111111: color_data = Z;
		19'b0000111110101000000: color_data = Z;
		19'b0000111110101000001: color_data = Z;
		19'b0000111110101000010: color_data = Z;
		19'b0000111110101000011: color_data = Z;
		19'b0000111110101000100: color_data = Z;
		19'b0000111110101000101: color_data = Z;
		19'b0000111110101000110: color_data = Z;
		19'b0000111110101000111: color_data = Z;
		19'b0000111110101001000: color_data = Z;
		19'b0000111110101001001: color_data = Z;
		19'b0000111110101001010: color_data = Z;
		19'b0000111110101001011: color_data = Z;
		19'b0000111110101001100: color_data = Z;
		19'b0000111110101001101: color_data = Z;
		19'b0000111110101001110: color_data = Z;
		19'b0000111110101001111: color_data = Z;
		19'b0000111110101010000: color_data = Z;
		19'b0000111110101010001: color_data = Z;
		19'b0000111110101010010: color_data = Z;
		19'b0000111110101010011: color_data = Z;
		19'b0000111110101010100: color_data = Z;
		19'b0000111110101010101: color_data = Z;
		19'b0000111110101010110: color_data = Z;
		19'b0000111110101010111: color_data = Z;
		19'b0000111110101011000: color_data = Z;
		19'b0000111110101011001: color_data = Z;
		19'b0000111110101011010: color_data = Z;
		19'b0000111110101011011: color_data = Z;
		19'b0000111110101011100: color_data = Z;
		19'b0000111110101011101: color_data = Z;
		19'b0000111110101011110: color_data = Z;
		19'b0000111110101011111: color_data = Z;
		19'b0000111110101100000: color_data = Z;
		19'b0000111110101100001: color_data = Z;
		19'b0000111110101100010: color_data = Z;
		19'b0000111110101100011: color_data = Z;
		19'b0000111110101100100: color_data = Z;
		19'b0000111110101100101: color_data = Z;
		19'b0000111110101100110: color_data = Z;
		19'b0000111110101100111: color_data = Z;
		19'b0000111110101101000: color_data = Z;
		19'b0000111110101101001: color_data = Z;
		19'b0000111110101101010: color_data = Z;
		19'b0000111110101101011: color_data = Z;
		19'b0000111110101101100: color_data = Z;
		19'b0000111110101101101: color_data = Z;
		19'b0000111110101101110: color_data = Z;
		19'b0000111110101101111: color_data = Z;
		19'b0000111110101110000: color_data = Z;
		19'b0000111110101110001: color_data = Z;
		19'b0000111110101110010: color_data = Z;
		19'b0000111110101110011: color_data = Z;
		19'b0000111110101110100: color_data = Z;
		19'b0000111110101110101: color_data = Z;
		19'b0000111110101110110: color_data = Z;
		19'b0000111110101110111: color_data = Z;
		19'b0000111110101111000: color_data = Z;
		19'b0000111110101111001: color_data = Z;
		19'b0000111110101111010: color_data = Z;
		19'b0000111110101111011: color_data = Z;
		19'b0000111110101111100: color_data = Z;
		19'b0000111110101111101: color_data = Z;
		19'b0000111110101111110: color_data = Z;
		19'b0000111110101111111: color_data = Z;
		19'b0000111110110000000: color_data = Z;
		19'b0000111110110000001: color_data = Z;
		19'b0000111110110000010: color_data = Z;
		19'b0000111110110000011: color_data = Z;
		19'b0000111110110000100: color_data = Z;
		19'b0000111110110000101: color_data = Z;
		19'b0000111110110000110: color_data = Z;
		19'b0000111110110000111: color_data = Z;
		19'b0000111110110001000: color_data = Z;
		19'b0000111110110001001: color_data = Z;
		19'b0000111110110001010: color_data = Z;
		19'b0000111110110001011: color_data = Z;
		19'b0000111110110001100: color_data = Z;
		19'b0000111110110001101: color_data = Z;
		19'b0000111110110001110: color_data = Z;
		19'b0000111110110001111: color_data = Z;
		19'b0000111110110010000: color_data = Z;
		19'b0000111110110010001: color_data = Z;
		19'b0000111110110010010: color_data = Z;
		19'b0000111110110010011: color_data = Z;
		19'b0000111110110010100: color_data = Z;
		19'b0000111110110010101: color_data = Z;
		19'b0000111110110010110: color_data = Z;
		19'b0000111110110010111: color_data = Z;
		19'b0000111110110011000: color_data = Z;
		19'b0001000000011101111: color_data = Z;
		19'b0001000000011110000: color_data = Z;
		19'b0001000000011110001: color_data = Z;
		19'b0001000000011110010: color_data = Z;
		19'b0001000000011110011: color_data = Z;
		19'b0001000000011110100: color_data = Z;
		19'b0001000000011110101: color_data = Z;
		19'b0001000000011110110: color_data = Z;
		19'b0001000000011110111: color_data = Z;
		19'b0001000000011111000: color_data = Z;
		19'b0001000000011111001: color_data = Z;
		19'b0001000000011111010: color_data = Z;
		19'b0001000000011111011: color_data = Z;
		19'b0001000000011111100: color_data = Z;
		19'b0001000000011111101: color_data = Z;
		19'b0001000000011111110: color_data = Z;
		19'b0001000000011111111: color_data = Z;
		19'b0001000000100000000: color_data = Z;
		19'b0001000000100000001: color_data = Z;
		19'b0001000000100000010: color_data = Z;
		19'b0001000000100000011: color_data = Z;
		19'b0001000000100000100: color_data = Z;
		19'b0001000000100000101: color_data = Z;
		19'b0001000000100000110: color_data = Z;
		19'b0001000000100000111: color_data = Z;
		19'b0001000000100001000: color_data = Z;
		19'b0001000000100001001: color_data = Z;
		19'b0001000000100001010: color_data = Z;
		19'b0001000000100001011: color_data = Z;
		19'b0001000000100001100: color_data = Z;
		19'b0001000000100001101: color_data = Z;
		19'b0001000000100001110: color_data = Z;
		19'b0001000000100001111: color_data = Z;
		19'b0001000000100010000: color_data = Z;
		19'b0001000000100010001: color_data = Z;
		19'b0001000000100010010: color_data = Z;
		19'b0001000000100010011: color_data = Z;
		19'b0001000000100010100: color_data = Z;
		19'b0001000000100010101: color_data = Z;
		19'b0001000000100010110: color_data = Z;
		19'b0001000000100010111: color_data = Z;
		19'b0001000000100011000: color_data = Z;
		19'b0001000000100011001: color_data = Z;
		19'b0001000000100011010: color_data = Z;
		19'b0001000000100011011: color_data = Z;
		19'b0001000000100011100: color_data = Z;
		19'b0001000000100011101: color_data = Z;
		19'b0001000000100011110: color_data = Z;
		19'b0001000000100011111: color_data = Z;
		19'b0001000000100100000: color_data = Z;
		19'b0001000000100100001: color_data = Z;
		19'b0001000000100100010: color_data = Z;
		19'b0001000000100100011: color_data = Z;
		19'b0001000000100100100: color_data = Z;
		19'b0001000000100100101: color_data = Z;
		19'b0001000000100100110: color_data = Z;
		19'b0001000000100100111: color_data = Z;
		19'b0001000000100101000: color_data = Z;
		19'b0001000000100101001: color_data = Z;
		19'b0001000000100101010: color_data = Z;
		19'b0001000000100101011: color_data = Z;
		19'b0001000000100101100: color_data = Z;
		19'b0001000000100101101: color_data = Z;
		19'b0001000000100101110: color_data = Z;
		19'b0001000000100101111: color_data = Z;
		19'b0001000000100110000: color_data = Z;
		19'b0001000000100110001: color_data = Z;
		19'b0001000000100110010: color_data = Z;
		19'b0001000000100110011: color_data = Z;
		19'b0001000000100110100: color_data = Z;
		19'b0001000000100110101: color_data = Z;
		19'b0001000000100110110: color_data = Z;
		19'b0001000000100110111: color_data = Z;
		19'b0001000000100111000: color_data = Z;
		19'b0001000000100111001: color_data = Z;
		19'b0001000000100111010: color_data = Z;
		19'b0001000000100111011: color_data = Z;
		19'b0001000000100111100: color_data = Z;
		19'b0001000000100111101: color_data = Z;
		19'b0001000000100111110: color_data = Z;
		19'b0001000000100111111: color_data = Z;
		19'b0001000000101000000: color_data = Z;
		19'b0001000000101000001: color_data = Z;
		19'b0001000000101000010: color_data = Z;
		19'b0001000000101000011: color_data = Z;
		19'b0001000000101000100: color_data = Z;
		19'b0001000000101000101: color_data = Z;
		19'b0001000000101000110: color_data = Z;
		19'b0001000000101000111: color_data = Z;
		19'b0001000000101001000: color_data = Z;
		19'b0001000000101001001: color_data = Z;
		19'b0001000000101001010: color_data = Z;
		19'b0001000000101001011: color_data = Z;
		19'b0001000000101001100: color_data = Z;
		19'b0001000000101001101: color_data = Z;
		19'b0001000000101001110: color_data = Z;
		19'b0001000000101001111: color_data = Z;
		19'b0001000000101010000: color_data = Z;
		19'b0001000000101010001: color_data = Z;
		19'b0001000000101010010: color_data = Z;
		19'b0001000000101010011: color_data = Z;
		19'b0001000000101010100: color_data = Z;
		19'b0001000000101010101: color_data = Z;
		19'b0001000000101010110: color_data = Z;
		19'b0001000000101010111: color_data = Z;
		19'b0001000000101011000: color_data = Z;
		19'b0001000000101011001: color_data = Z;
		19'b0001000000101011010: color_data = Z;
		19'b0001000000101011011: color_data = Z;
		19'b0001000000101011100: color_data = Z;
		19'b0001000000101011101: color_data = Z;
		19'b0001000000101011110: color_data = Z;
		19'b0001000000101011111: color_data = Z;
		19'b0001000000101100000: color_data = Z;
		19'b0001000000101100001: color_data = Z;
		19'b0001000000101100010: color_data = Z;
		19'b0001000000101100011: color_data = Z;
		19'b0001000000101100100: color_data = Z;
		19'b0001000000101100101: color_data = Z;
		19'b0001000000101100110: color_data = Z;
		19'b0001000000101100111: color_data = Z;
		19'b0001000000101101000: color_data = Z;
		19'b0001000000101101001: color_data = Z;
		19'b0001000000101101010: color_data = Z;
		19'b0001000000101101011: color_data = Z;
		19'b0001000000101101100: color_data = Z;
		19'b0001000000101101101: color_data = Z;
		19'b0001000000101101110: color_data = Z;
		19'b0001000000101101111: color_data = Z;
		19'b0001000000101110000: color_data = Z;
		19'b0001000000101110001: color_data = Z;
		19'b0001000000101110010: color_data = Z;
		19'b0001000000101110011: color_data = Z;
		19'b0001000000101110100: color_data = Z;
		19'b0001000000101110101: color_data = Z;
		19'b0001000000101110110: color_data = Z;
		19'b0001000000101110111: color_data = Z;
		19'b0001000000101111000: color_data = Z;
		19'b0001000000101111001: color_data = Z;
		19'b0001000000101111010: color_data = Z;
		19'b0001000000101111011: color_data = Z;
		19'b0001000000101111100: color_data = Z;
		19'b0001000000101111101: color_data = Z;
		19'b0001000000101111110: color_data = Z;
		19'b0001000000101111111: color_data = Z;
		19'b0001000000110000000: color_data = Z;
		19'b0001000000110000001: color_data = Z;
		19'b0001000000110000010: color_data = Z;
		19'b0001000000110000011: color_data = Z;
		19'b0001000000110000100: color_data = Z;
		19'b0001000000110000101: color_data = Z;
		19'b0001000000110000110: color_data = Z;
		19'b0001000000110000111: color_data = Z;
		19'b0001000000110001000: color_data = Z;
		19'b0001000000110001001: color_data = Z;
		19'b0001000000110001010: color_data = Z;
		19'b0001000000110001011: color_data = Z;
		19'b0001000000110001100: color_data = Z;
		19'b0001000000110001101: color_data = Z;
		19'b0001000000110001110: color_data = Z;
		19'b0001000000110001111: color_data = Z;
		19'b0001000000110010000: color_data = Z;
		19'b0001000000110010001: color_data = Z;
		19'b0001000000110010010: color_data = Z;
		19'b0001000000110010011: color_data = Z;
		19'b0001000000110010100: color_data = Z;
		19'b0001000000110010101: color_data = Z;
		19'b0001000000110010110: color_data = Z;
		19'b0001000000110010111: color_data = Z;
		19'b0001000000110011000: color_data = Z;
		19'b0001000000110011001: color_data = Z;
		19'b0001000010011101110: color_data = Z;
		19'b0001000010011101111: color_data = Z;
		19'b0001000010011110000: color_data = Z;
		19'b0001000010011110001: color_data = Z;
		19'b0001000010011110010: color_data = Z;
		19'b0001000010011110011: color_data = Z;
		19'b0001000010011110100: color_data = Z;
		19'b0001000010011110101: color_data = Z;
		19'b0001000010011110110: color_data = Z;
		19'b0001000010011110111: color_data = Z;
		19'b0001000010011111000: color_data = Z;
		19'b0001000010011111001: color_data = Z;
		19'b0001000010011111010: color_data = Z;
		19'b0001000010011111011: color_data = Z;
		19'b0001000010011111100: color_data = Z;
		19'b0001000010011111101: color_data = Z;
		19'b0001000010011111110: color_data = Z;
		19'b0001000010011111111: color_data = Z;
		19'b0001000010100000000: color_data = Z;
		19'b0001000010100000001: color_data = Z;
		19'b0001000010100000010: color_data = Z;
		19'b0001000010100000011: color_data = Z;
		19'b0001000010100000100: color_data = Z;
		19'b0001000010100000101: color_data = Z;
		19'b0001000010100000110: color_data = Z;
		19'b0001000010100000111: color_data = Z;
		19'b0001000010100001000: color_data = Z;
		19'b0001000010100001001: color_data = Z;
		19'b0001000010100001010: color_data = Z;
		19'b0001000010100001011: color_data = Z;
		19'b0001000010100001100: color_data = Z;
		19'b0001000010100001101: color_data = Z;
		19'b0001000010100001110: color_data = Z;
		19'b0001000010100001111: color_data = Z;
		19'b0001000010100010000: color_data = Z;
		19'b0001000010100010001: color_data = Z;
		19'b0001000010100010010: color_data = Z;
		19'b0001000010100010011: color_data = Z;
		19'b0001000010100010100: color_data = Z;
		19'b0001000010100010101: color_data = Z;
		19'b0001000010100010110: color_data = Z;
		19'b0001000010100010111: color_data = Z;
		19'b0001000010100011000: color_data = Z;
		19'b0001000010100011001: color_data = Z;
		19'b0001000010100011010: color_data = Z;
		19'b0001000010100011011: color_data = Z;
		19'b0001000010100011100: color_data = Z;
		19'b0001000010100011101: color_data = Z;
		19'b0001000010100011110: color_data = Z;
		19'b0001000010100011111: color_data = Z;
		19'b0001000010100100000: color_data = Z;
		19'b0001000010100100001: color_data = Z;
		19'b0001000010100100010: color_data = Z;
		19'b0001000010100100011: color_data = Z;
		19'b0001000010100100100: color_data = Z;
		19'b0001000010100100101: color_data = Z;
		19'b0001000010100100110: color_data = Z;
		19'b0001000010100100111: color_data = Z;
		19'b0001000010100101000: color_data = Z;
		19'b0001000010100101001: color_data = Z;
		19'b0001000010100101010: color_data = Z;
		19'b0001000010100101011: color_data = Z;
		19'b0001000010100101100: color_data = Z;
		19'b0001000010100101101: color_data = Z;
		19'b0001000010100101110: color_data = Z;
		19'b0001000010100101111: color_data = Z;
		19'b0001000010100110000: color_data = Z;
		19'b0001000010100110001: color_data = Z;
		19'b0001000010100110010: color_data = Z;
		19'b0001000010100110011: color_data = Z;
		19'b0001000010100110100: color_data = Z;
		19'b0001000010100110101: color_data = Z;
		19'b0001000010100110110: color_data = Z;
		19'b0001000010100110111: color_data = Z;
		19'b0001000010100111000: color_data = Z;
		19'b0001000010100111001: color_data = Z;
		19'b0001000010100111010: color_data = Z;
		19'b0001000010100111011: color_data = Z;
		19'b0001000010100111100: color_data = Z;
		19'b0001000010100111101: color_data = Z;
		19'b0001000010100111110: color_data = Z;
		19'b0001000010100111111: color_data = Z;
		19'b0001000010101000000: color_data = Z;
		19'b0001000010101000001: color_data = Z;
		19'b0001000010101000010: color_data = Z;
		19'b0001000010101000011: color_data = Z;
		19'b0001000010101000100: color_data = Z;
		19'b0001000010101000101: color_data = Z;
		19'b0001000010101000110: color_data = Z;
		19'b0001000010101000111: color_data = Z;
		19'b0001000010101001000: color_data = Z;
		19'b0001000010101001001: color_data = Z;
		19'b0001000010101001010: color_data = Z;
		19'b0001000010101001011: color_data = Z;
		19'b0001000010101001100: color_data = Z;
		19'b0001000010101001101: color_data = Z;
		19'b0001000010101001110: color_data = Z;
		19'b0001000010101001111: color_data = Z;
		19'b0001000010101010000: color_data = Z;
		19'b0001000010101010001: color_data = Z;
		19'b0001000010101010010: color_data = Z;
		19'b0001000010101010011: color_data = Z;
		19'b0001000010101010100: color_data = Z;
		19'b0001000010101010101: color_data = Z;
		19'b0001000010101010110: color_data = Z;
		19'b0001000010101010111: color_data = Z;
		19'b0001000010101011000: color_data = Z;
		19'b0001000010101011001: color_data = Z;
		19'b0001000010101011010: color_data = Z;
		19'b0001000010101011011: color_data = Z;
		19'b0001000010101011100: color_data = Z;
		19'b0001000010101011101: color_data = Z;
		19'b0001000010101011110: color_data = Z;
		19'b0001000010101011111: color_data = Z;
		19'b0001000010101100000: color_data = Z;
		19'b0001000010101100001: color_data = Z;
		19'b0001000010101100010: color_data = Z;
		19'b0001000010101100011: color_data = Z;
		19'b0001000010101100100: color_data = Z;
		19'b0001000010101100101: color_data = Z;
		19'b0001000010101100110: color_data = Z;
		19'b0001000010101100111: color_data = Z;
		19'b0001000010101101000: color_data = Z;
		19'b0001000010101101001: color_data = Z;
		19'b0001000010101101010: color_data = Z;
		19'b0001000010101101011: color_data = Z;
		19'b0001000010101101100: color_data = Z;
		19'b0001000010101101101: color_data = Z;
		19'b0001000010101101110: color_data = Z;
		19'b0001000010101101111: color_data = Z;
		19'b0001000010101110000: color_data = Z;
		19'b0001000010101110001: color_data = Z;
		19'b0001000010101110010: color_data = Z;
		19'b0001000010101110011: color_data = Z;
		19'b0001000010101110100: color_data = Z;
		19'b0001000010101110101: color_data = Z;
		19'b0001000010101110110: color_data = Z;
		19'b0001000010101110111: color_data = Z;
		19'b0001000010101111000: color_data = Z;
		19'b0001000010101111001: color_data = Z;
		19'b0001000010101111010: color_data = Z;
		19'b0001000010101111011: color_data = Z;
		19'b0001000010101111100: color_data = Z;
		19'b0001000010101111101: color_data = Z;
		19'b0001000010101111110: color_data = Z;
		19'b0001000010101111111: color_data = Z;
		19'b0001000010110000000: color_data = Z;
		19'b0001000010110000001: color_data = Z;
		19'b0001000010110000010: color_data = Z;
		19'b0001000010110000011: color_data = Z;
		19'b0001000010110000100: color_data = Z;
		19'b0001000010110000101: color_data = Z;
		19'b0001000010110000110: color_data = Z;
		19'b0001000010110000111: color_data = Z;
		19'b0001000010110001000: color_data = Z;
		19'b0001000010110001001: color_data = Z;
		19'b0001000010110001010: color_data = Z;
		19'b0001000010110001011: color_data = Z;
		19'b0001000010110001100: color_data = Z;
		19'b0001000010110001101: color_data = Z;
		19'b0001000010110001110: color_data = Z;
		19'b0001000010110001111: color_data = Z;
		19'b0001000010110010000: color_data = Z;
		19'b0001000010110010001: color_data = Z;
		19'b0001000010110010010: color_data = Z;
		19'b0001000010110010011: color_data = Z;
		19'b0001000010110010100: color_data = Z;
		19'b0001000010110010101: color_data = Z;
		19'b0001000010110010110: color_data = Z;
		19'b0001000010110010111: color_data = Z;
		19'b0001000010110011000: color_data = Z;
		19'b0001000010110011001: color_data = Z;
		19'b0001000010110011010: color_data = Z;
		19'b0001000100011101100: color_data = Z;
		19'b0001000100011101101: color_data = Z;
		19'b0001000100011101110: color_data = Z;
		19'b0001000100011101111: color_data = Z;
		19'b0001000100011110000: color_data = Z;
		19'b0001000100011110001: color_data = Z;
		19'b0001000100011110010: color_data = Z;
		19'b0001000100011110011: color_data = Z;
		19'b0001000100011110100: color_data = Z;
		19'b0001000100011110101: color_data = Z;
		19'b0001000100011110110: color_data = Z;
		19'b0001000100011110111: color_data = Z;
		19'b0001000100011111000: color_data = Z;
		19'b0001000100011111001: color_data = Z;
		19'b0001000100011111010: color_data = Z;
		19'b0001000100011111011: color_data = Z;
		19'b0001000100011111100: color_data = Z;
		19'b0001000100011111101: color_data = Z;
		19'b0001000100011111110: color_data = Z;
		19'b0001000100011111111: color_data = Z;
		19'b0001000100100000000: color_data = Z;
		19'b0001000100100000001: color_data = Z;
		19'b0001000100100000010: color_data = Z;
		19'b0001000100100000011: color_data = Z;
		19'b0001000100100000100: color_data = Z;
		19'b0001000100100000101: color_data = Z;
		19'b0001000100100000110: color_data = Z;
		19'b0001000100100000111: color_data = Z;
		19'b0001000100100001000: color_data = Z;
		19'b0001000100100001001: color_data = Z;
		19'b0001000100100001010: color_data = Z;
		19'b0001000100100001011: color_data = Z;
		19'b0001000100100001100: color_data = Z;
		19'b0001000100100001101: color_data = Z;
		19'b0001000100100001110: color_data = Z;
		19'b0001000100100001111: color_data = Z;
		19'b0001000100100010000: color_data = Z;
		19'b0001000100100010001: color_data = Z;
		19'b0001000100100010010: color_data = Z;
		19'b0001000100100010011: color_data = Z;
		19'b0001000100100010100: color_data = Z;
		19'b0001000100100010101: color_data = Z;
		19'b0001000100100010110: color_data = Z;
		19'b0001000100100010111: color_data = Z;
		19'b0001000100100011000: color_data = Z;
		19'b0001000100100011001: color_data = Z;
		19'b0001000100100011010: color_data = Z;
		19'b0001000100100011011: color_data = Z;
		19'b0001000100100011100: color_data = Z;
		19'b0001000100100011101: color_data = Z;
		19'b0001000100100011110: color_data = Z;
		19'b0001000100100011111: color_data = Z;
		19'b0001000100100100000: color_data = Z;
		19'b0001000100100100001: color_data = Z;
		19'b0001000100100100010: color_data = Z;
		19'b0001000100100100011: color_data = Z;
		19'b0001000100100100100: color_data = Z;
		19'b0001000100100100101: color_data = Z;
		19'b0001000100100100110: color_data = Z;
		19'b0001000100100100111: color_data = Z;
		19'b0001000100100101000: color_data = Z;
		19'b0001000100100101001: color_data = Z;
		19'b0001000100100101010: color_data = Z;
		19'b0001000100100101011: color_data = Z;
		19'b0001000100100101100: color_data = Z;
		19'b0001000100100101101: color_data = Z;
		19'b0001000100100101110: color_data = Z;
		19'b0001000100100101111: color_data = Z;
		19'b0001000100100110000: color_data = Z;
		19'b0001000100100110001: color_data = Z;
		19'b0001000100100110010: color_data = Z;
		19'b0001000100100110011: color_data = Z;
		19'b0001000100100110100: color_data = Z;
		19'b0001000100100110101: color_data = Z;
		19'b0001000100100110110: color_data = Z;
		19'b0001000100100110111: color_data = Z;
		19'b0001000100100111000: color_data = Z;
		19'b0001000100100111001: color_data = Z;
		19'b0001000100100111010: color_data = Z;
		19'b0001000100100111011: color_data = Z;
		19'b0001000100100111100: color_data = Z;
		19'b0001000100100111101: color_data = Z;
		19'b0001000100100111110: color_data = Z;
		19'b0001000100100111111: color_data = Z;
		19'b0001000100101000000: color_data = Z;
		19'b0001000100101000001: color_data = Z;
		19'b0001000100101000010: color_data = Z;
		19'b0001000100101000011: color_data = Z;
		19'b0001000100101000100: color_data = Z;
		19'b0001000100101000101: color_data = Z;
		19'b0001000100101000110: color_data = Z;
		19'b0001000100101000111: color_data = Z;
		19'b0001000100101001000: color_data = Z;
		19'b0001000100101001001: color_data = Z;
		19'b0001000100101001010: color_data = Z;
		19'b0001000100101001011: color_data = Z;
		19'b0001000100101001100: color_data = Z;
		19'b0001000100101001101: color_data = Z;
		19'b0001000100101001110: color_data = Z;
		19'b0001000100101001111: color_data = Z;
		19'b0001000100101010000: color_data = Z;
		19'b0001000100101010001: color_data = Z;
		19'b0001000100101010010: color_data = Z;
		19'b0001000100101010011: color_data = Z;
		19'b0001000100101010100: color_data = Z;
		19'b0001000100101010101: color_data = Z;
		19'b0001000100101010110: color_data = Z;
		19'b0001000100101010111: color_data = Z;
		19'b0001000100101011000: color_data = Z;
		19'b0001000100101011001: color_data = Z;
		19'b0001000100101011010: color_data = Z;
		19'b0001000100101011011: color_data = Z;
		19'b0001000100101011100: color_data = Z;
		19'b0001000100101011101: color_data = Z;
		19'b0001000100101011110: color_data = Z;
		19'b0001000100101011111: color_data = Z;
		19'b0001000100101100000: color_data = Z;
		19'b0001000100101100001: color_data = Z;
		19'b0001000100101100010: color_data = Z;
		19'b0001000100101100011: color_data = Z;
		19'b0001000100101100100: color_data = Z;
		19'b0001000100101100101: color_data = Z;
		19'b0001000100101100110: color_data = Z;
		19'b0001000100101100111: color_data = Z;
		19'b0001000100101101000: color_data = Z;
		19'b0001000100101101001: color_data = Z;
		19'b0001000100101101010: color_data = Z;
		19'b0001000100101101011: color_data = Z;
		19'b0001000100101101100: color_data = Z;
		19'b0001000100101101101: color_data = Z;
		19'b0001000100101101110: color_data = Z;
		19'b0001000100101101111: color_data = Z;
		19'b0001000100101110000: color_data = Z;
		19'b0001000100101110001: color_data = Z;
		19'b0001000100101110010: color_data = Z;
		19'b0001000100101110011: color_data = Z;
		19'b0001000100101110100: color_data = Z;
		19'b0001000100101110101: color_data = Z;
		19'b0001000100101110110: color_data = Z;
		19'b0001000100101110111: color_data = Z;
		19'b0001000100101111000: color_data = Z;
		19'b0001000100101111001: color_data = Z;
		19'b0001000100101111010: color_data = Z;
		19'b0001000100101111011: color_data = Z;
		19'b0001000100101111100: color_data = Z;
		19'b0001000100101111101: color_data = Z;
		19'b0001000100101111110: color_data = Z;
		19'b0001000100101111111: color_data = Z;
		19'b0001000100110000000: color_data = Z;
		19'b0001000100110000001: color_data = Z;
		19'b0001000100110000010: color_data = Z;
		19'b0001000100110000011: color_data = Z;
		19'b0001000100110000100: color_data = Z;
		19'b0001000100110000101: color_data = Z;
		19'b0001000100110000110: color_data = Z;
		19'b0001000100110000111: color_data = Z;
		19'b0001000100110001000: color_data = Z;
		19'b0001000100110001001: color_data = Z;
		19'b0001000100110001010: color_data = Z;
		19'b0001000100110001011: color_data = Z;
		19'b0001000100110001100: color_data = Z;
		19'b0001000100110001101: color_data = Z;
		19'b0001000100110001110: color_data = Z;
		19'b0001000100110001111: color_data = Z;
		19'b0001000100110010000: color_data = Z;
		19'b0001000100110010001: color_data = Z;
		19'b0001000100110010010: color_data = Z;
		19'b0001000100110010011: color_data = Z;
		19'b0001000100110010100: color_data = Z;
		19'b0001000100110010101: color_data = Z;
		19'b0001000100110010110: color_data = Z;
		19'b0001000100110010111: color_data = Z;
		19'b0001000100110011000: color_data = Z;
		19'b0001000100110011001: color_data = Z;
		19'b0001000100110011010: color_data = Z;
		19'b0001000110011101100: color_data = Z;
		19'b0001000110011101101: color_data = Z;
		19'b0001000110011101110: color_data = Z;
		19'b0001000110011101111: color_data = Z;
		19'b0001000110011110000: color_data = Z;
		19'b0001000110011110001: color_data = Z;
		19'b0001000110011110010: color_data = Z;
		19'b0001000110011110011: color_data = Z;
		19'b0001000110011110100: color_data = Z;
		19'b0001000110011110101: color_data = Z;
		19'b0001000110011110110: color_data = Z;
		19'b0001000110011110111: color_data = Z;
		19'b0001000110011111000: color_data = Z;
		19'b0001000110011111001: color_data = Z;
		19'b0001000110011111010: color_data = Z;
		19'b0001000110011111011: color_data = Z;
		19'b0001000110011111100: color_data = Z;
		19'b0001000110011111101: color_data = Z;
		19'b0001000110011111110: color_data = Z;
		19'b0001000110011111111: color_data = Z;
		19'b0001000110100000000: color_data = Z;
		19'b0001000110100000001: color_data = Z;
		19'b0001000110100000010: color_data = Z;
		19'b0001000110100000011: color_data = Z;
		19'b0001000110100000100: color_data = Z;
		19'b0001000110100000101: color_data = Z;
		19'b0001000110100000110: color_data = Z;
		19'b0001000110100000111: color_data = Z;
		19'b0001000110100001000: color_data = Z;
		19'b0001000110100001001: color_data = Z;
		19'b0001000110100001010: color_data = Z;
		19'b0001000110100001011: color_data = Z;
		19'b0001000110100001100: color_data = Z;
		19'b0001000110100001101: color_data = Z;
		19'b0001000110100001110: color_data = Z;
		19'b0001000110100001111: color_data = Z;
		19'b0001000110100010000: color_data = Z;
		19'b0001000110100010001: color_data = Z;
		19'b0001000110100010010: color_data = Z;
		19'b0001000110100010011: color_data = Z;
		19'b0001000110100010100: color_data = Z;
		19'b0001000110100010101: color_data = Z;
		19'b0001000110100010110: color_data = Z;
		19'b0001000110100010111: color_data = Z;
		19'b0001000110100011000: color_data = Z;
		19'b0001000110100011001: color_data = Z;
		19'b0001000110100011010: color_data = Z;
		19'b0001000110100011011: color_data = Z;
		19'b0001000110100011100: color_data = Z;
		19'b0001000110100011101: color_data = Z;
		19'b0001000110100011110: color_data = Z;
		19'b0001000110100011111: color_data = Z;
		19'b0001000110100100000: color_data = Z;
		19'b0001000110100100001: color_data = Z;
		19'b0001000110100100010: color_data = Z;
		19'b0001000110100100011: color_data = Z;
		19'b0001000110100100100: color_data = Z;
		19'b0001000110100100101: color_data = Z;
		19'b0001000110100100110: color_data = Z;
		19'b0001000110100100111: color_data = Z;
		19'b0001000110100101000: color_data = Z;
		19'b0001000110100101001: color_data = Z;
		19'b0001000110100101010: color_data = Z;
		19'b0001000110100101011: color_data = Z;
		19'b0001000110100101100: color_data = Z;
		19'b0001000110100101101: color_data = Z;
		19'b0001000110100101110: color_data = Z;
		19'b0001000110100101111: color_data = Z;
		19'b0001000110100110000: color_data = Z;
		19'b0001000110100110001: color_data = Z;
		19'b0001000110100110010: color_data = Z;
		19'b0001000110100110011: color_data = Z;
		19'b0001000110100110100: color_data = Z;
		19'b0001000110100110101: color_data = Z;
		19'b0001000110100110110: color_data = Z;
		19'b0001000110100110111: color_data = Z;
		19'b0001000110100111000: color_data = Z;
		19'b0001000110100111001: color_data = Z;
		19'b0001000110100111010: color_data = Z;
		19'b0001000110100111011: color_data = Z;
		19'b0001000110100111100: color_data = Z;
		19'b0001000110100111101: color_data = Z;
		19'b0001000110100111110: color_data = Z;
		19'b0001000110100111111: color_data = Z;
		19'b0001000110101000000: color_data = Z;
		19'b0001000110101000001: color_data = Z;
		19'b0001000110101000010: color_data = Z;
		19'b0001000110101000011: color_data = Z;
		19'b0001000110101000100: color_data = Z;
		19'b0001000110101000101: color_data = Z;
		19'b0001000110101000110: color_data = Z;
		19'b0001000110101000111: color_data = Z;
		19'b0001000110101001000: color_data = Z;
		19'b0001000110101001001: color_data = Z;
		19'b0001000110101001010: color_data = Z;
		19'b0001000110101001011: color_data = Z;
		19'b0001000110101001100: color_data = Z;
		19'b0001000110101001101: color_data = Z;
		19'b0001000110101001110: color_data = Z;
		19'b0001000110101001111: color_data = Z;
		19'b0001000110101010000: color_data = Z;
		19'b0001000110101010001: color_data = Z;
		19'b0001000110101010010: color_data = Z;
		19'b0001000110101010011: color_data = Z;
		19'b0001000110101010100: color_data = Z;
		19'b0001000110101010101: color_data = Z;
		19'b0001000110101010110: color_data = Z;
		19'b0001000110101010111: color_data = Z;
		19'b0001000110101011000: color_data = Z;
		19'b0001000110101011001: color_data = Z;
		19'b0001000110101011010: color_data = Z;
		19'b0001000110101011011: color_data = Z;
		19'b0001000110101011100: color_data = Z;
		19'b0001000110101011101: color_data = Z;
		19'b0001000110101011110: color_data = Z;
		19'b0001000110101011111: color_data = Z;
		19'b0001000110101100000: color_data = Z;
		19'b0001000110101100001: color_data = Z;
		19'b0001000110101100010: color_data = Z;
		19'b0001000110101100011: color_data = Z;
		19'b0001000110101100100: color_data = Z;
		19'b0001000110101100101: color_data = Z;
		19'b0001000110101100110: color_data = Z;
		19'b0001000110101100111: color_data = Z;
		19'b0001000110101101000: color_data = Z;
		19'b0001000110101101001: color_data = Z;
		19'b0001000110101101010: color_data = Z;
		19'b0001000110101101011: color_data = Z;
		19'b0001000110101101100: color_data = Z;
		19'b0001000110101101101: color_data = Z;
		19'b0001000110101101110: color_data = Z;
		19'b0001000110101101111: color_data = Z;
		19'b0001000110101110000: color_data = Z;
		19'b0001000110101110001: color_data = Z;
		19'b0001000110101110010: color_data = Z;
		19'b0001000110101110011: color_data = Z;
		19'b0001000110101110100: color_data = Z;
		19'b0001000110101110101: color_data = Z;
		19'b0001000110101110110: color_data = Z;
		19'b0001000110101110111: color_data = Z;
		19'b0001000110101111000: color_data = Z;
		19'b0001000110101111001: color_data = Z;
		19'b0001000110101111010: color_data = Z;
		19'b0001000110101111011: color_data = Z;
		19'b0001000110101111100: color_data = Z;
		19'b0001000110101111101: color_data = Z;
		19'b0001000110101111110: color_data = Z;
		19'b0001000110101111111: color_data = Z;
		19'b0001000110110000000: color_data = Z;
		19'b0001000110110000001: color_data = Z;
		19'b0001000110110000010: color_data = Z;
		19'b0001000110110000011: color_data = Z;
		19'b0001000110110000100: color_data = Z;
		19'b0001000110110000101: color_data = Z;
		19'b0001000110110000110: color_data = Z;
		19'b0001000110110000111: color_data = Z;
		19'b0001000110110001000: color_data = Z;
		19'b0001000110110001001: color_data = Z;
		19'b0001000110110001010: color_data = Z;
		19'b0001000110110001011: color_data = Z;
		19'b0001000110110001100: color_data = Z;
		19'b0001000110110001101: color_data = Z;
		19'b0001000110110001110: color_data = Z;
		19'b0001000110110001111: color_data = Z;
		19'b0001000110110010000: color_data = Z;
		19'b0001000110110010001: color_data = Z;
		19'b0001000110110010010: color_data = Z;
		19'b0001000110110010011: color_data = Z;
		19'b0001000110110010100: color_data = Z;
		19'b0001000110110010101: color_data = Z;
		19'b0001000110110010110: color_data = Z;
		19'b0001000110110010111: color_data = Z;
		19'b0001000110110011000: color_data = Z;
		19'b0001000110110011001: color_data = Z;
		19'b0001000110110011010: color_data = Z;
		19'b0001000110110011011: color_data = Z;
		19'b0001001000011101011: color_data = Z;
		19'b0001001000011101100: color_data = Z;
		19'b0001001000011101101: color_data = Z;
		19'b0001001000011101110: color_data = Z;
		19'b0001001000011101111: color_data = Z;
		19'b0001001000011110000: color_data = Z;
		19'b0001001000011110001: color_data = Z;
		19'b0001001000011110010: color_data = Z;
		19'b0001001000011110011: color_data = Z;
		19'b0001001000011110100: color_data = Z;
		19'b0001001000011110101: color_data = Z;
		19'b0001001000011110110: color_data = Z;
		19'b0001001000011110111: color_data = Z;
		19'b0001001000011111000: color_data = Z;
		19'b0001001000011111001: color_data = Z;
		19'b0001001000011111010: color_data = Z;
		19'b0001001000011111011: color_data = Z;
		19'b0001001000011111100: color_data = Z;
		19'b0001001000011111101: color_data = Z;
		19'b0001001000011111110: color_data = Z;
		19'b0001001000011111111: color_data = Z;
		19'b0001001000100000000: color_data = Z;
		19'b0001001000100000001: color_data = Z;
		19'b0001001000100000010: color_data = Z;
		19'b0001001000100000011: color_data = Z;
		19'b0001001000100000100: color_data = Z;
		19'b0001001000100000101: color_data = Z;
		19'b0001001000100000110: color_data = Z;
		19'b0001001000100000111: color_data = Z;
		19'b0001001000100001000: color_data = Z;
		19'b0001001000100001001: color_data = Z;
		19'b0001001000100001010: color_data = Z;
		19'b0001001000100001011: color_data = Z;
		19'b0001001000100001100: color_data = Z;
		19'b0001001000100001101: color_data = Z;
		19'b0001001000100001110: color_data = Z;
		19'b0001001000100001111: color_data = Z;
		19'b0001001000100010000: color_data = Z;
		19'b0001001000100010001: color_data = Z;
		19'b0001001000100010010: color_data = Z;
		19'b0001001000100010011: color_data = Z;
		19'b0001001000100010100: color_data = Z;
		19'b0001001000100010101: color_data = Z;
		19'b0001001000100010110: color_data = Z;
		19'b0001001000100010111: color_data = Z;
		19'b0001001000100011000: color_data = Z;
		19'b0001001000100011001: color_data = Z;
		19'b0001001000100011010: color_data = Z;
		19'b0001001000100011011: color_data = Z;
		19'b0001001000100011100: color_data = Z;
		19'b0001001000100011101: color_data = Z;
		19'b0001001000100011110: color_data = Z;
		19'b0001001000100011111: color_data = Z;
		19'b0001001000100100000: color_data = Z;
		19'b0001001000100100001: color_data = Z;
		19'b0001001000100100010: color_data = Z;
		19'b0001001000100100011: color_data = Z;
		19'b0001001000100100100: color_data = Z;
		19'b0001001000100100101: color_data = Z;
		19'b0001001000100100110: color_data = Z;
		19'b0001001000100100111: color_data = Z;
		19'b0001001000100101000: color_data = Z;
		19'b0001001000100101001: color_data = Z;
		19'b0001001000100101010: color_data = Z;
		19'b0001001000100101011: color_data = Z;
		19'b0001001000100101100: color_data = Z;
		19'b0001001000100101101: color_data = Z;
		19'b0001001000100101110: color_data = Z;
		19'b0001001000100101111: color_data = Z;
		19'b0001001000100110000: color_data = Z;
		19'b0001001000100110001: color_data = Z;
		19'b0001001000100110010: color_data = Z;
		19'b0001001000100110011: color_data = Z;
		19'b0001001000100110100: color_data = Z;
		19'b0001001000100110101: color_data = Z;
		19'b0001001000100110110: color_data = Z;
		19'b0001001000100110111: color_data = Z;
		19'b0001001000100111000: color_data = Z;
		19'b0001001000100111001: color_data = Z;
		19'b0001001000100111010: color_data = Z;
		19'b0001001000100111011: color_data = Z;
		19'b0001001000100111100: color_data = Z;
		19'b0001001000100111101: color_data = Z;
		19'b0001001000100111110: color_data = Z;
		19'b0001001000100111111: color_data = Z;
		19'b0001001000101000000: color_data = Z;
		19'b0001001000101000001: color_data = Z;
		19'b0001001000101000010: color_data = Z;
		19'b0001001000101000011: color_data = Z;
		19'b0001001000101000100: color_data = Z;
		19'b0001001000101000101: color_data = Z;
		19'b0001001000101000110: color_data = Z;
		19'b0001001000101000111: color_data = Z;
		19'b0001001000101001000: color_data = Z;
		19'b0001001000101001001: color_data = Z;
		19'b0001001000101001010: color_data = Z;
		19'b0001001000101001011: color_data = Z;
		19'b0001001000101001100: color_data = Z;
		19'b0001001000101001101: color_data = Z;
		19'b0001001000101001110: color_data = Z;
		19'b0001001000101001111: color_data = Z;
		19'b0001001000101010000: color_data = Z;
		19'b0001001000101010001: color_data = Z;
		19'b0001001000101010010: color_data = Z;
		19'b0001001000101010011: color_data = Z;
		19'b0001001000101010100: color_data = Z;
		19'b0001001000101010101: color_data = Z;
		19'b0001001000101010110: color_data = Z;
		19'b0001001000101010111: color_data = Z;
		19'b0001001000101011000: color_data = Z;
		19'b0001001000101011001: color_data = Z;
		19'b0001001000101011010: color_data = Z;
		19'b0001001000101011011: color_data = Z;
		19'b0001001000101011100: color_data = Z;
		19'b0001001000101011101: color_data = Z;
		19'b0001001000101011110: color_data = Z;
		19'b0001001000101011111: color_data = Z;
		19'b0001001000101100000: color_data = Z;
		19'b0001001000101100001: color_data = Z;
		19'b0001001000101100010: color_data = Z;
		19'b0001001000101100011: color_data = Z;
		19'b0001001000101100100: color_data = Z;
		19'b0001001000101100101: color_data = Z;
		19'b0001001000101100110: color_data = Z;
		19'b0001001000101100111: color_data = Z;
		19'b0001001000101101000: color_data = Z;
		19'b0001001000101101001: color_data = Z;
		19'b0001001000101101010: color_data = Z;
		19'b0001001000101101011: color_data = Z;
		19'b0001001000101101100: color_data = Z;
		19'b0001001000101101101: color_data = Z;
		19'b0001001000101101110: color_data = Z;
		19'b0001001000101101111: color_data = Z;
		19'b0001001000101110000: color_data = Z;
		19'b0001001000101110001: color_data = Z;
		19'b0001001000101110010: color_data = Z;
		19'b0001001000101110011: color_data = Z;
		19'b0001001000101110100: color_data = Z;
		19'b0001001000101110101: color_data = Z;
		19'b0001001000101110110: color_data = Z;
		19'b0001001000101110111: color_data = Z;
		19'b0001001000101111000: color_data = Z;
		19'b0001001000101111001: color_data = Z;
		19'b0001001000101111010: color_data = Z;
		19'b0001001000101111011: color_data = Z;
		19'b0001001000101111100: color_data = Z;
		19'b0001001000101111101: color_data = Z;
		19'b0001001000101111110: color_data = Z;
		19'b0001001000101111111: color_data = Z;
		19'b0001001000110000000: color_data = Z;
		19'b0001001000110000001: color_data = Z;
		19'b0001001000110000010: color_data = Z;
		19'b0001001000110000011: color_data = Z;
		19'b0001001000110000100: color_data = Z;
		19'b0001001000110000101: color_data = Z;
		19'b0001001000110000110: color_data = Z;
		19'b0001001000110000111: color_data = Z;
		19'b0001001000110001000: color_data = Z;
		19'b0001001000110001001: color_data = Z;
		19'b0001001000110001010: color_data = Z;
		19'b0001001000110001011: color_data = Z;
		19'b0001001000110001100: color_data = Z;
		19'b0001001000110001101: color_data = Z;
		19'b0001001000110001110: color_data = Z;
		19'b0001001000110001111: color_data = Z;
		19'b0001001000110010000: color_data = Z;
		19'b0001001000110010001: color_data = Z;
		19'b0001001000110010010: color_data = Z;
		19'b0001001000110010011: color_data = Z;
		19'b0001001000110010100: color_data = Z;
		19'b0001001000110010101: color_data = Z;
		19'b0001001000110010110: color_data = Z;
		19'b0001001000110010111: color_data = Z;
		19'b0001001000110011000: color_data = Z;
		19'b0001001000110011001: color_data = Z;
		19'b0001001000110011010: color_data = Z;
		19'b0001001000110011011: color_data = Z;
		19'b0001001010011101011: color_data = Z;
		19'b0001001010011101100: color_data = Z;
		19'b0001001010011101101: color_data = Z;
		19'b0001001010011101110: color_data = Z;
		19'b0001001010011101111: color_data = Z;
		19'b0001001010011110000: color_data = Z;
		19'b0001001010011110001: color_data = Z;
		19'b0001001010011110010: color_data = Z;
		19'b0001001010011110011: color_data = Z;
		19'b0001001010011110100: color_data = Z;
		19'b0001001010011110101: color_data = Z;
		19'b0001001010011110110: color_data = Z;
		19'b0001001010011110111: color_data = Z;
		19'b0001001010011111000: color_data = Z;
		19'b0001001010011111001: color_data = Z;
		19'b0001001010011111010: color_data = Z;
		19'b0001001010011111011: color_data = Z;
		19'b0001001010011111100: color_data = Z;
		19'b0001001010011111101: color_data = Z;
		19'b0001001010011111110: color_data = Z;
		19'b0001001010011111111: color_data = Z;
		19'b0001001010100000000: color_data = Z;
		19'b0001001010100000001: color_data = Z;
		19'b0001001010100000010: color_data = Z;
		19'b0001001010100000011: color_data = Z;
		19'b0001001010100000100: color_data = Z;
		19'b0001001010100000101: color_data = Z;
		19'b0001001010100000110: color_data = Z;
		19'b0001001010100000111: color_data = Z;
		19'b0001001010100001000: color_data = Z;
		19'b0001001010100001001: color_data = Z;
		19'b0001001010100001010: color_data = Z;
		19'b0001001010100001011: color_data = Z;
		19'b0001001010100001100: color_data = Z;
		19'b0001001010100001101: color_data = Z;
		19'b0001001010100001110: color_data = Z;
		19'b0001001010100001111: color_data = Z;
		19'b0001001010100010000: color_data = Z;
		19'b0001001010100010001: color_data = Z;
		19'b0001001010100010010: color_data = Z;
		19'b0001001010100010011: color_data = Z;
		19'b0001001010100010100: color_data = Z;
		19'b0001001010100010101: color_data = Z;
		19'b0001001010100010110: color_data = Z;
		19'b0001001010100010111: color_data = Z;
		19'b0001001010100011000: color_data = Z;
		19'b0001001010100011001: color_data = Z;
		19'b0001001010100011010: color_data = Z;
		19'b0001001010100011011: color_data = Z;
		19'b0001001010100011100: color_data = Z;
		19'b0001001010100011101: color_data = Z;
		19'b0001001010100011110: color_data = Z;
		19'b0001001010100011111: color_data = Z;
		19'b0001001010100100000: color_data = Z;
		19'b0001001010100100001: color_data = Z;
		19'b0001001010100100010: color_data = Z;
		19'b0001001010100100011: color_data = Z;
		19'b0001001010100100100: color_data = Z;
		19'b0001001010100100101: color_data = Z;
		19'b0001001010100100110: color_data = Z;
		19'b0001001010100100111: color_data = Z;
		19'b0001001010100101000: color_data = Z;
		19'b0001001010100101001: color_data = Z;
		19'b0001001010100101010: color_data = Z;
		19'b0001001010100101011: color_data = Z;
		19'b0001001010100101100: color_data = Z;
		19'b0001001010100101101: color_data = Z;
		19'b0001001010100101110: color_data = Z;
		19'b0001001010100101111: color_data = Z;
		19'b0001001010100110000: color_data = Z;
		19'b0001001010100110001: color_data = Z;
		19'b0001001010100110010: color_data = Z;
		19'b0001001010100110011: color_data = Z;
		19'b0001001010100110100: color_data = Z;
		19'b0001001010100110101: color_data = Z;
		19'b0001001010100110110: color_data = Z;
		19'b0001001010100110111: color_data = Z;
		19'b0001001010100111000: color_data = Z;
		19'b0001001010100111001: color_data = Z;
		19'b0001001010100111010: color_data = Z;
		19'b0001001010100111011: color_data = Z;
		19'b0001001010100111100: color_data = Z;
		19'b0001001010100111101: color_data = Z;
		19'b0001001010100111110: color_data = Z;
		19'b0001001010100111111: color_data = Z;
		19'b0001001010101000000: color_data = Z;
		19'b0001001010101000001: color_data = Z;
		19'b0001001010101000010: color_data = Z;
		19'b0001001010101000011: color_data = Z;
		19'b0001001010101000100: color_data = Z;
		19'b0001001010101000101: color_data = Z;
		19'b0001001010101000110: color_data = Z;
		19'b0001001010101000111: color_data = Z;
		19'b0001001010101001000: color_data = Z;
		19'b0001001010101001001: color_data = Z;
		19'b0001001010101001010: color_data = Z;
		19'b0001001010101001011: color_data = Z;
		19'b0001001010101001100: color_data = Z;
		19'b0001001010101001101: color_data = Z;
		19'b0001001010101001110: color_data = Z;
		19'b0001001010101001111: color_data = Z;
		19'b0001001010101010000: color_data = Z;
		19'b0001001010101010001: color_data = Z;
		19'b0001001010101010010: color_data = Z;
		19'b0001001010101010011: color_data = Z;
		19'b0001001010101010100: color_data = Z;
		19'b0001001010101010101: color_data = Z;
		19'b0001001010101010110: color_data = Z;
		19'b0001001010101010111: color_data = Z;
		19'b0001001010101011000: color_data = Z;
		19'b0001001010101011001: color_data = Z;
		19'b0001001010101011010: color_data = Z;
		19'b0001001010101011011: color_data = Z;
		19'b0001001010101011100: color_data = Z;
		19'b0001001010101011101: color_data = Z;
		19'b0001001010101011110: color_data = Z;
		19'b0001001010101011111: color_data = Z;
		19'b0001001010101100000: color_data = Z;
		19'b0001001010101100001: color_data = Z;
		19'b0001001010101100010: color_data = Z;
		19'b0001001010101100011: color_data = Z;
		19'b0001001010101100100: color_data = Z;
		19'b0001001010101100101: color_data = Z;
		19'b0001001010101100110: color_data = Z;
		19'b0001001010101100111: color_data = Z;
		19'b0001001010101101000: color_data = Z;
		19'b0001001010101101001: color_data = Z;
		19'b0001001010101101010: color_data = Z;
		19'b0001001010101101011: color_data = Z;
		19'b0001001010101101100: color_data = Z;
		19'b0001001010101101101: color_data = Z;
		19'b0001001010101101110: color_data = Z;
		19'b0001001010101101111: color_data = Z;
		19'b0001001010101110000: color_data = Z;
		19'b0001001010101110001: color_data = Z;
		19'b0001001010101110010: color_data = Z;
		19'b0001001010101110011: color_data = Z;
		19'b0001001010101110100: color_data = Z;
		19'b0001001010101110101: color_data = Z;
		19'b0001001010101110110: color_data = Z;
		19'b0001001010101110111: color_data = Z;
		19'b0001001010101111000: color_data = Z;
		19'b0001001010101111001: color_data = Z;
		19'b0001001010101111010: color_data = Z;
		19'b0001001010101111011: color_data = Z;
		19'b0001001010101111100: color_data = Z;
		19'b0001001010101111101: color_data = Z;
		19'b0001001010101111110: color_data = Z;
		19'b0001001010101111111: color_data = Z;
		19'b0001001010110000000: color_data = Z;
		19'b0001001010110000001: color_data = Z;
		19'b0001001010110000010: color_data = Z;
		19'b0001001010110000011: color_data = Z;
		19'b0001001010110000100: color_data = Z;
		19'b0001001010110000101: color_data = Z;
		19'b0001001010110000110: color_data = Z;
		19'b0001001010110000111: color_data = Z;
		19'b0001001010110001000: color_data = Z;
		19'b0001001010110001001: color_data = Z;
		19'b0001001010110001010: color_data = Z;
		19'b0001001010110001011: color_data = Z;
		19'b0001001010110001100: color_data = Z;
		19'b0001001010110001101: color_data = Z;
		19'b0001001010110001110: color_data = Z;
		19'b0001001010110001111: color_data = Z;
		19'b0001001010110010000: color_data = Z;
		19'b0001001010110010001: color_data = Z;
		19'b0001001010110010010: color_data = Z;
		19'b0001001010110010011: color_data = Z;
		19'b0001001010110010100: color_data = Z;
		19'b0001001010110010101: color_data = Z;
		19'b0001001010110010110: color_data = Z;
		19'b0001001010110010111: color_data = Z;
		19'b0001001010110011000: color_data = Z;
		19'b0001001010110011001: color_data = Z;
		19'b0001001010110011010: color_data = Z;
		19'b0001001010110011011: color_data = Z;
		19'b0001001010110100000: color_data = Z;
		19'b0001001010110100001: color_data = Z;
		19'b0001001010110100010: color_data = Z;
		19'b0001001100011101010: color_data = Z;
		19'b0001001100011101011: color_data = Z;
		19'b0001001100011101100: color_data = Z;
		19'b0001001100011101101: color_data = Z;
		19'b0001001100011101110: color_data = Z;
		19'b0001001100011101111: color_data = Z;
		19'b0001001100011110000: color_data = Z;
		19'b0001001100011110001: color_data = Z;
		19'b0001001100011110010: color_data = Z;
		19'b0001001100011110011: color_data = Z;
		19'b0001001100011110100: color_data = Z;
		19'b0001001100011110101: color_data = Z;
		19'b0001001100011110110: color_data = Z;
		19'b0001001100011110111: color_data = Z;
		19'b0001001100011111000: color_data = Z;
		19'b0001001100011111001: color_data = Z;
		19'b0001001100011111010: color_data = Z;
		19'b0001001100011111011: color_data = Z;
		19'b0001001100011111100: color_data = Z;
		19'b0001001100011111101: color_data = Z;
		19'b0001001100011111110: color_data = Z;
		19'b0001001100011111111: color_data = Z;
		19'b0001001100100000000: color_data = Z;
		19'b0001001100100000001: color_data = Z;
		19'b0001001100100000010: color_data = Z;
		19'b0001001100100000011: color_data = Z;
		19'b0001001100100000100: color_data = Z;
		19'b0001001100100000101: color_data = Z;
		19'b0001001100100000110: color_data = Z;
		19'b0001001100100000111: color_data = Z;
		19'b0001001100100001000: color_data = Z;
		19'b0001001100100001001: color_data = Z;
		19'b0001001100100001010: color_data = Z;
		19'b0001001100100001011: color_data = Z;
		19'b0001001100100001100: color_data = Z;
		19'b0001001100100001101: color_data = Z;
		19'b0001001100100001110: color_data = Z;
		19'b0001001100100001111: color_data = Z;
		19'b0001001100100010000: color_data = Z;
		19'b0001001100100010001: color_data = Z;
		19'b0001001100100010010: color_data = Z;
		19'b0001001100100010011: color_data = Z;
		19'b0001001100100010100: color_data = Z;
		19'b0001001100100010101: color_data = Z;
		19'b0001001100100010110: color_data = Z;
		19'b0001001100100010111: color_data = Z;
		19'b0001001100100011000: color_data = Z;
		19'b0001001100100011001: color_data = Z;
		19'b0001001100100011010: color_data = Z;
		19'b0001001100100011011: color_data = Z;
		19'b0001001100100011100: color_data = Z;
		19'b0001001100100011101: color_data = Z;
		19'b0001001100100011110: color_data = Z;
		19'b0001001100100011111: color_data = Z;
		19'b0001001100100100000: color_data = Z;
		19'b0001001100100100001: color_data = Z;
		19'b0001001100100100010: color_data = Z;
		19'b0001001100100100011: color_data = Z;
		19'b0001001100100100100: color_data = Z;
		19'b0001001100100100101: color_data = Z;
		19'b0001001100100100110: color_data = Z;
		19'b0001001100100100111: color_data = Z;
		19'b0001001100100101000: color_data = Z;
		19'b0001001100100101001: color_data = Z;
		19'b0001001100100101010: color_data = Z;
		19'b0001001100100101011: color_data = Z;
		19'b0001001100100101100: color_data = Z;
		19'b0001001100100101101: color_data = Z;
		19'b0001001100100101110: color_data = Z;
		19'b0001001100100101111: color_data = Z;
		19'b0001001100100110000: color_data = Z;
		19'b0001001100100110001: color_data = Z;
		19'b0001001100100110010: color_data = Z;
		19'b0001001100100110011: color_data = Z;
		19'b0001001100100110100: color_data = Z;
		19'b0001001100100110101: color_data = Z;
		19'b0001001100100110110: color_data = Z;
		19'b0001001100100110111: color_data = Z;
		19'b0001001100100111000: color_data = Z;
		19'b0001001100100111001: color_data = Z;
		19'b0001001100100111010: color_data = Z;
		19'b0001001100100111011: color_data = Z;
		19'b0001001100100111100: color_data = Z;
		19'b0001001100100111101: color_data = Z;
		19'b0001001100100111110: color_data = Z;
		19'b0001001100100111111: color_data = Z;
		19'b0001001100101000000: color_data = Z;
		19'b0001001100101000001: color_data = Z;
		19'b0001001100101000010: color_data = Z;
		19'b0001001100101000011: color_data = Z;
		19'b0001001100101000100: color_data = Z;
		19'b0001001100101000101: color_data = Z;
		19'b0001001100101000110: color_data = Z;
		19'b0001001100101000111: color_data = Z;
		19'b0001001100101001000: color_data = Z;
		19'b0001001100101001001: color_data = Z;
		19'b0001001100101001010: color_data = Z;
		19'b0001001100101001011: color_data = Z;
		19'b0001001100101001100: color_data = Z;
		19'b0001001100101001101: color_data = Z;
		19'b0001001100101001110: color_data = Z;
		19'b0001001100101001111: color_data = Z;
		19'b0001001100101010000: color_data = Z;
		19'b0001001100101010001: color_data = Z;
		19'b0001001100101010010: color_data = Z;
		19'b0001001100101010011: color_data = Z;
		19'b0001001100101010100: color_data = Z;
		19'b0001001100101010101: color_data = Z;
		19'b0001001100101010110: color_data = Z;
		19'b0001001100101010111: color_data = Z;
		19'b0001001100101011000: color_data = Z;
		19'b0001001100101011001: color_data = Z;
		19'b0001001100101011010: color_data = Z;
		19'b0001001100101011011: color_data = Z;
		19'b0001001100101011100: color_data = Z;
		19'b0001001100101011101: color_data = Z;
		19'b0001001100101011110: color_data = Z;
		19'b0001001100101011111: color_data = Z;
		19'b0001001100101100000: color_data = Z;
		19'b0001001100101100001: color_data = Z;
		19'b0001001100101100010: color_data = Z;
		19'b0001001100101100011: color_data = Z;
		19'b0001001100101100100: color_data = Z;
		19'b0001001100101100101: color_data = Z;
		19'b0001001100101100110: color_data = Z;
		19'b0001001100101100111: color_data = Z;
		19'b0001001100101101000: color_data = Z;
		19'b0001001100101101001: color_data = Z;
		19'b0001001100101101010: color_data = Z;
		19'b0001001100101101011: color_data = Z;
		19'b0001001100101101100: color_data = Z;
		19'b0001001100101101101: color_data = Z;
		19'b0001001100101101110: color_data = Z;
		19'b0001001100101101111: color_data = Z;
		19'b0001001100101110000: color_data = Z;
		19'b0001001100101110001: color_data = Z;
		19'b0001001100101110010: color_data = Z;
		19'b0001001100101110011: color_data = Z;
		19'b0001001100101110100: color_data = Z;
		19'b0001001100101110101: color_data = Z;
		19'b0001001100101110110: color_data = Z;
		19'b0001001100101110111: color_data = Z;
		19'b0001001100101111000: color_data = Z;
		19'b0001001100101111001: color_data = Z;
		19'b0001001100101111010: color_data = Z;
		19'b0001001100101111011: color_data = Z;
		19'b0001001100101111100: color_data = Z;
		19'b0001001100101111101: color_data = Z;
		19'b0001001100101111110: color_data = Z;
		19'b0001001100101111111: color_data = Z;
		19'b0001001100110000000: color_data = Z;
		19'b0001001100110000001: color_data = Z;
		19'b0001001100110000010: color_data = Z;
		19'b0001001100110000011: color_data = Z;
		19'b0001001100110000100: color_data = Z;
		19'b0001001100110000101: color_data = Z;
		19'b0001001100110000110: color_data = Z;
		19'b0001001100110000111: color_data = Z;
		19'b0001001100110001000: color_data = Z;
		19'b0001001100110001001: color_data = Z;
		19'b0001001100110001010: color_data = Z;
		19'b0001001100110001011: color_data = Z;
		19'b0001001100110001100: color_data = Z;
		19'b0001001100110001101: color_data = Z;
		19'b0001001100110001110: color_data = Z;
		19'b0001001100110001111: color_data = Z;
		19'b0001001100110010000: color_data = Z;
		19'b0001001100110010001: color_data = Z;
		19'b0001001100110010010: color_data = Z;
		19'b0001001100110010011: color_data = Z;
		19'b0001001100110010100: color_data = Z;
		19'b0001001100110010101: color_data = Z;
		19'b0001001100110010110: color_data = Z;
		19'b0001001100110010111: color_data = Z;
		19'b0001001100110011000: color_data = Z;
		19'b0001001100110011001: color_data = Z;
		19'b0001001100110011010: color_data = Z;
		19'b0001001100110011011: color_data = Z;
		19'b0001001100110100000: color_data = Z;
		19'b0001001100110100001: color_data = Z;
		19'b0001001100110100010: color_data = Z;
		19'b0001001100110100011: color_data = Z;
		19'b0001001100110100100: color_data = Z;
		19'b0001001100110100101: color_data = Z;
		19'b0001001110011101001: color_data = Z;
		19'b0001001110011101010: color_data = Z;
		19'b0001001110011101011: color_data = Z;
		19'b0001001110011101100: color_data = Z;
		19'b0001001110011101101: color_data = Z;
		19'b0001001110011101110: color_data = Z;
		19'b0001001110011101111: color_data = Z;
		19'b0001001110011110000: color_data = Z;
		19'b0001001110011110001: color_data = Z;
		19'b0001001110011110010: color_data = Z;
		19'b0001001110011110011: color_data = Z;
		19'b0001001110011110100: color_data = Z;
		19'b0001001110011110101: color_data = Z;
		19'b0001001110011110110: color_data = Z;
		19'b0001001110011110111: color_data = Z;
		19'b0001001110011111000: color_data = Z;
		19'b0001001110011111001: color_data = Z;
		19'b0001001110011111010: color_data = Z;
		19'b0001001110011111011: color_data = Z;
		19'b0001001110011111100: color_data = Z;
		19'b0001001110011111101: color_data = Z;
		19'b0001001110011111110: color_data = Z;
		19'b0001001110011111111: color_data = Z;
		19'b0001001110100000000: color_data = Z;
		19'b0001001110100000001: color_data = Z;
		19'b0001001110100000010: color_data = Z;
		19'b0001001110100000011: color_data = Z;
		19'b0001001110100000100: color_data = Z;
		19'b0001001110100000101: color_data = Z;
		19'b0001001110100000110: color_data = Z;
		19'b0001001110100000111: color_data = Z;
		19'b0001001110100001000: color_data = Z;
		19'b0001001110100001001: color_data = Z;
		19'b0001001110100001010: color_data = Z;
		19'b0001001110100001011: color_data = Z;
		19'b0001001110100001100: color_data = Z;
		19'b0001001110100001101: color_data = Z;
		19'b0001001110100001110: color_data = Z;
		19'b0001001110100001111: color_data = Z;
		19'b0001001110100010000: color_data = Z;
		19'b0001001110100010001: color_data = Z;
		19'b0001001110100010010: color_data = Z;
		19'b0001001110100010011: color_data = Z;
		19'b0001001110100010100: color_data = Z;
		19'b0001001110100010101: color_data = Z;
		19'b0001001110100010110: color_data = Z;
		19'b0001001110100010111: color_data = Z;
		19'b0001001110100011000: color_data = Z;
		19'b0001001110100011001: color_data = Z;
		19'b0001001110100011010: color_data = Z;
		19'b0001001110100011011: color_data = Z;
		19'b0001001110100011100: color_data = Z;
		19'b0001001110100011101: color_data = Z;
		19'b0001001110100011110: color_data = Z;
		19'b0001001110100011111: color_data = Z;
		19'b0001001110100100000: color_data = Z;
		19'b0001001110100100001: color_data = Z;
		19'b0001001110100100010: color_data = Z;
		19'b0001001110100100011: color_data = Z;
		19'b0001001110100100100: color_data = Z;
		19'b0001001110100100101: color_data = Z;
		19'b0001001110100100110: color_data = Z;
		19'b0001001110100100111: color_data = Z;
		19'b0001001110100101000: color_data = Z;
		19'b0001001110100101001: color_data = Z;
		19'b0001001110100101010: color_data = Z;
		19'b0001001110100101011: color_data = Z;
		19'b0001001110100101100: color_data = Z;
		19'b0001001110100101101: color_data = Z;
		19'b0001001110100101110: color_data = Z;
		19'b0001001110100101111: color_data = Z;
		19'b0001001110100110000: color_data = Z;
		19'b0001001110100110001: color_data = Z;
		19'b0001001110100110010: color_data = Z;
		19'b0001001110100110011: color_data = Z;
		19'b0001001110100110100: color_data = Z;
		19'b0001001110100110101: color_data = Z;
		19'b0001001110100110110: color_data = Z;
		19'b0001001110100110111: color_data = Z;
		19'b0001001110100111000: color_data = Z;
		19'b0001001110100111001: color_data = Z;
		19'b0001001110100111010: color_data = Z;
		19'b0001001110100111011: color_data = Z;
		19'b0001001110100111100: color_data = Z;
		19'b0001001110100111101: color_data = Z;
		19'b0001001110100111110: color_data = Z;
		19'b0001001110100111111: color_data = Z;
		19'b0001001110101000000: color_data = Z;
		19'b0001001110101000001: color_data = Z;
		19'b0001001110101000010: color_data = Z;
		19'b0001001110101000011: color_data = Z;
		19'b0001001110101000100: color_data = Z;
		19'b0001001110101000101: color_data = Z;
		19'b0001001110101000110: color_data = Z;
		19'b0001001110101000111: color_data = Z;
		19'b0001001110101001000: color_data = Z;
		19'b0001001110101001001: color_data = Z;
		19'b0001001110101001010: color_data = Z;
		19'b0001001110101001011: color_data = Z;
		19'b0001001110101001100: color_data = Z;
		19'b0001001110101001101: color_data = Z;
		19'b0001001110101001110: color_data = Z;
		19'b0001001110101001111: color_data = Z;
		19'b0001001110101010000: color_data = Z;
		19'b0001001110101010001: color_data = Z;
		19'b0001001110101010010: color_data = Z;
		19'b0001001110101010011: color_data = Z;
		19'b0001001110101010100: color_data = Z;
		19'b0001001110101010101: color_data = Z;
		19'b0001001110101010110: color_data = Z;
		19'b0001001110101010111: color_data = Z;
		19'b0001001110101011000: color_data = Z;
		19'b0001001110101011001: color_data = Z;
		19'b0001001110101011010: color_data = Z;
		19'b0001001110101011011: color_data = Z;
		19'b0001001110101011100: color_data = Z;
		19'b0001001110101011101: color_data = Z;
		19'b0001001110101011110: color_data = Z;
		19'b0001001110101011111: color_data = Z;
		19'b0001001110101100000: color_data = Z;
		19'b0001001110101100001: color_data = Z;
		19'b0001001110101100010: color_data = Z;
		19'b0001001110101100011: color_data = Z;
		19'b0001001110101100100: color_data = Z;
		19'b0001001110101100101: color_data = Z;
		19'b0001001110101100110: color_data = Z;
		19'b0001001110101100111: color_data = Z;
		19'b0001001110101101000: color_data = Z;
		19'b0001001110101101001: color_data = Z;
		19'b0001001110101101010: color_data = Z;
		19'b0001001110101101011: color_data = Z;
		19'b0001001110101101100: color_data = Z;
		19'b0001001110101101101: color_data = Z;
		19'b0001001110101101110: color_data = Z;
		19'b0001001110101101111: color_data = Z;
		19'b0001001110101110000: color_data = Z;
		19'b0001001110101110001: color_data = Z;
		19'b0001001110101110010: color_data = Z;
		19'b0001001110101110011: color_data = Z;
		19'b0001001110101110100: color_data = Z;
		19'b0001001110101110101: color_data = Z;
		19'b0001001110101110110: color_data = Z;
		19'b0001001110101110111: color_data = Z;
		19'b0001001110101111000: color_data = Z;
		19'b0001001110101111001: color_data = Z;
		19'b0001001110101111010: color_data = Z;
		19'b0001001110101111011: color_data = Z;
		19'b0001001110101111100: color_data = Z;
		19'b0001001110101111101: color_data = Z;
		19'b0001001110101111110: color_data = Z;
		19'b0001001110101111111: color_data = Z;
		19'b0001001110110000000: color_data = Z;
		19'b0001001110110000001: color_data = Z;
		19'b0001001110110000010: color_data = Z;
		19'b0001001110110000011: color_data = Z;
		19'b0001001110110000100: color_data = Z;
		19'b0001001110110000101: color_data = Z;
		19'b0001001110110000110: color_data = Z;
		19'b0001001110110000111: color_data = Z;
		19'b0001001110110001000: color_data = Z;
		19'b0001001110110001001: color_data = Z;
		19'b0001001110110001010: color_data = Z;
		19'b0001001110110001011: color_data = Z;
		19'b0001001110110001100: color_data = Z;
		19'b0001001110110001101: color_data = Z;
		19'b0001001110110001110: color_data = Z;
		19'b0001001110110001111: color_data = Z;
		19'b0001001110110010000: color_data = Z;
		19'b0001001110110010001: color_data = Z;
		19'b0001001110110010010: color_data = Z;
		19'b0001001110110010011: color_data = Z;
		19'b0001001110110010100: color_data = Z;
		19'b0001001110110010101: color_data = Z;
		19'b0001001110110010110: color_data = Z;
		19'b0001001110110010111: color_data = Z;
		19'b0001001110110011000: color_data = Z;
		19'b0001001110110011001: color_data = Z;
		19'b0001001110110011010: color_data = Z;
		19'b0001001110110011011: color_data = Z;
		19'b0001001110110100000: color_data = Z;
		19'b0001001110110100001: color_data = Z;
		19'b0001001110110100010: color_data = Z;
		19'b0001001110110100011: color_data = Z;
		19'b0001001110110100100: color_data = Z;
		19'b0001001110110100101: color_data = Z;
		19'b0001001110110100110: color_data = Z;
		19'b0001001110110100111: color_data = Z;
		19'b0001010000011100111: color_data = Z;
		19'b0001010000011101000: color_data = Z;
		19'b0001010000011101001: color_data = Z;
		19'b0001010000011101010: color_data = Z;
		19'b0001010000011101011: color_data = Z;
		19'b0001010000011101100: color_data = Z;
		19'b0001010000011101101: color_data = Z;
		19'b0001010000011101110: color_data = Z;
		19'b0001010000011101111: color_data = Z;
		19'b0001010000011110000: color_data = Z;
		19'b0001010000011110001: color_data = Z;
		19'b0001010000011110010: color_data = Z;
		19'b0001010000011110011: color_data = Z;
		19'b0001010000011110100: color_data = Z;
		19'b0001010000011110101: color_data = Z;
		19'b0001010000011110110: color_data = Z;
		19'b0001010000011110111: color_data = Z;
		19'b0001010000011111000: color_data = Z;
		19'b0001010000011111001: color_data = Z;
		19'b0001010000011111010: color_data = Z;
		19'b0001010000011111011: color_data = Z;
		19'b0001010000011111100: color_data = Z;
		19'b0001010000011111101: color_data = Z;
		19'b0001010000011111110: color_data = Z;
		19'b0001010000011111111: color_data = Z;
		19'b0001010000100000000: color_data = Z;
		19'b0001010000100000001: color_data = Z;
		19'b0001010000100000010: color_data = Z;
		19'b0001010000100000011: color_data = Z;
		19'b0001010000100000100: color_data = Z;
		19'b0001010000100000101: color_data = Z;
		19'b0001010000100000110: color_data = Z;
		19'b0001010000100000111: color_data = Z;
		19'b0001010000100001000: color_data = Z;
		19'b0001010000100001001: color_data = Z;
		19'b0001010000100001010: color_data = Z;
		19'b0001010000100001011: color_data = Z;
		19'b0001010000100001100: color_data = Z;
		19'b0001010000100001101: color_data = Z;
		19'b0001010000100001110: color_data = Z;
		19'b0001010000100001111: color_data = Z;
		19'b0001010000100010000: color_data = Z;
		19'b0001010000100010001: color_data = Z;
		19'b0001010000100010010: color_data = Z;
		19'b0001010000100010011: color_data = Z;
		19'b0001010000100010100: color_data = Z;
		19'b0001010000100010101: color_data = Z;
		19'b0001010000100010110: color_data = Z;
		19'b0001010000100010111: color_data = Z;
		19'b0001010000100011000: color_data = Z;
		19'b0001010000100011001: color_data = Z;
		19'b0001010000100011010: color_data = Z;
		19'b0001010000100011011: color_data = Z;
		19'b0001010000100011100: color_data = Z;
		19'b0001010000100011101: color_data = Z;
		19'b0001010000100011110: color_data = Z;
		19'b0001010000100011111: color_data = Z;
		19'b0001010000100100000: color_data = Z;
		19'b0001010000100100001: color_data = Z;
		19'b0001010000100100010: color_data = Z;
		19'b0001010000100100011: color_data = Z;
		19'b0001010000100100100: color_data = Z;
		19'b0001010000100100101: color_data = Z;
		19'b0001010000100100110: color_data = Z;
		19'b0001010000100100111: color_data = Z;
		19'b0001010000100101000: color_data = Z;
		19'b0001010000100101001: color_data = Z;
		19'b0001010000100101010: color_data = Z;
		19'b0001010000100101011: color_data = Z;
		19'b0001010000100101100: color_data = Z;
		19'b0001010000100101101: color_data = Z;
		19'b0001010000100101110: color_data = Z;
		19'b0001010000100101111: color_data = Z;
		19'b0001010000100110000: color_data = Z;
		19'b0001010000100110001: color_data = Z;
		19'b0001010000100110010: color_data = Z;
		19'b0001010000100110011: color_data = Z;
		19'b0001010000100110100: color_data = Z;
		19'b0001010000100110101: color_data = Z;
		19'b0001010000100110110: color_data = Z;
		19'b0001010000100110111: color_data = Z;
		19'b0001010000100111000: color_data = Z;
		19'b0001010000100111001: color_data = Z;
		19'b0001010000100111010: color_data = Z;
		19'b0001010000100111011: color_data = Z;
		19'b0001010000100111100: color_data = Z;
		19'b0001010000100111101: color_data = Z;
		19'b0001010000100111110: color_data = Z;
		19'b0001010000100111111: color_data = Z;
		19'b0001010000101000000: color_data = Z;
		19'b0001010000101000001: color_data = Z;
		19'b0001010000101000010: color_data = Z;
		19'b0001010000101000011: color_data = Z;
		19'b0001010000101000100: color_data = Z;
		19'b0001010000101000101: color_data = Z;
		19'b0001010000101000110: color_data = Z;
		19'b0001010000101000111: color_data = Z;
		19'b0001010000101001000: color_data = Z;
		19'b0001010000101001001: color_data = Z;
		19'b0001010000101001010: color_data = Z;
		19'b0001010000101001011: color_data = Z;
		19'b0001010000101001100: color_data = Z;
		19'b0001010000101001101: color_data = Z;
		19'b0001010000101001110: color_data = Z;
		19'b0001010000101001111: color_data = Z;
		19'b0001010000101010000: color_data = Z;
		19'b0001010000101010001: color_data = Z;
		19'b0001010000101010010: color_data = Z;
		19'b0001010000101010011: color_data = Z;
		19'b0001010000101010100: color_data = Z;
		19'b0001010000101010101: color_data = Z;
		19'b0001010000101010110: color_data = Z;
		19'b0001010000101010111: color_data = Z;
		19'b0001010000101011000: color_data = Z;
		19'b0001010000101011001: color_data = Z;
		19'b0001010000101011010: color_data = Z;
		19'b0001010000101011011: color_data = Z;
		19'b0001010000101011100: color_data = Z;
		19'b0001010000101011101: color_data = Z;
		19'b0001010000101011110: color_data = Z;
		19'b0001010000101011111: color_data = Z;
		19'b0001010000101100000: color_data = Z;
		19'b0001010000101100001: color_data = Z;
		19'b0001010000101100010: color_data = Z;
		19'b0001010000101100011: color_data = Z;
		19'b0001010000101100100: color_data = Z;
		19'b0001010000101100101: color_data = Z;
		19'b0001010000101100110: color_data = Z;
		19'b0001010000101100111: color_data = Z;
		19'b0001010000101101000: color_data = Z;
		19'b0001010000101101001: color_data = Z;
		19'b0001010000101101010: color_data = Z;
		19'b0001010000101101011: color_data = Z;
		19'b0001010000101101100: color_data = Z;
		19'b0001010000101101101: color_data = Z;
		19'b0001010000101101110: color_data = Z;
		19'b0001010000101101111: color_data = Z;
		19'b0001010000101110000: color_data = Z;
		19'b0001010000101110001: color_data = Z;
		19'b0001010000101110010: color_data = Z;
		19'b0001010000101110011: color_data = Z;
		19'b0001010000101110100: color_data = Z;
		19'b0001010000101110101: color_data = Z;
		19'b0001010000101110110: color_data = Z;
		19'b0001010000101110111: color_data = Z;
		19'b0001010000101111000: color_data = Z;
		19'b0001010000101111001: color_data = Z;
		19'b0001010000101111010: color_data = Z;
		19'b0001010000101111011: color_data = Z;
		19'b0001010000101111100: color_data = Z;
		19'b0001010000101111101: color_data = Z;
		19'b0001010000101111110: color_data = Z;
		19'b0001010000101111111: color_data = Z;
		19'b0001010000110000000: color_data = Z;
		19'b0001010000110000001: color_data = Z;
		19'b0001010000110000010: color_data = Z;
		19'b0001010000110000011: color_data = Z;
		19'b0001010000110000100: color_data = Z;
		19'b0001010000110000101: color_data = Z;
		19'b0001010000110000110: color_data = Z;
		19'b0001010000110000111: color_data = Z;
		19'b0001010000110001000: color_data = Z;
		19'b0001010000110001001: color_data = Z;
		19'b0001010000110001010: color_data = Z;
		19'b0001010000110001011: color_data = Z;
		19'b0001010000110001100: color_data = Z;
		19'b0001010000110001101: color_data = Z;
		19'b0001010000110001110: color_data = Z;
		19'b0001010000110001111: color_data = Z;
		19'b0001010000110010000: color_data = Z;
		19'b0001010000110010001: color_data = Z;
		19'b0001010000110010010: color_data = Z;
		19'b0001010000110010011: color_data = Z;
		19'b0001010000110010100: color_data = Z;
		19'b0001010000110010101: color_data = Z;
		19'b0001010000110010110: color_data = Z;
		19'b0001010000110010111: color_data = Z;
		19'b0001010000110011000: color_data = Z;
		19'b0001010000110011001: color_data = Z;
		19'b0001010000110011010: color_data = Z;
		19'b0001010000110011011: color_data = Z;
		19'b0001010000110100001: color_data = Z;
		19'b0001010000110100010: color_data = Z;
		19'b0001010000110100011: color_data = Z;
		19'b0001010000110100100: color_data = Z;
		19'b0001010000110100101: color_data = Z;
		19'b0001010000110100110: color_data = Z;
		19'b0001010000110100111: color_data = Z;
		19'b0001010000110101000: color_data = Z;
		19'b0001010010011100101: color_data = Z;
		19'b0001010010011100110: color_data = Z;
		19'b0001010010011100111: color_data = Z;
		19'b0001010010011101000: color_data = Z;
		19'b0001010010011101001: color_data = Z;
		19'b0001010010011101010: color_data = Z;
		19'b0001010010011101011: color_data = Z;
		19'b0001010010011101100: color_data = Z;
		19'b0001010010011101101: color_data = Z;
		19'b0001010010011101110: color_data = Z;
		19'b0001010010011101111: color_data = Z;
		19'b0001010010011110000: color_data = Z;
		19'b0001010010011110001: color_data = Z;
		19'b0001010010011110010: color_data = Z;
		19'b0001010010011110011: color_data = Z;
		19'b0001010010011110100: color_data = Z;
		19'b0001010010011110101: color_data = Z;
		19'b0001010010011110110: color_data = Z;
		19'b0001010010011110111: color_data = Z;
		19'b0001010010011111000: color_data = Z;
		19'b0001010010011111001: color_data = Z;
		19'b0001010010011111010: color_data = Z;
		19'b0001010010011111011: color_data = Z;
		19'b0001010010011111100: color_data = Z;
		19'b0001010010011111101: color_data = Z;
		19'b0001010010011111110: color_data = Z;
		19'b0001010010011111111: color_data = Z;
		19'b0001010010100000000: color_data = Z;
		19'b0001010010100000001: color_data = Z;
		19'b0001010010100000010: color_data = Z;
		19'b0001010010100000011: color_data = Z;
		19'b0001010010100000100: color_data = Z;
		19'b0001010010100000101: color_data = Z;
		19'b0001010010100000110: color_data = Z;
		19'b0001010010100000111: color_data = Z;
		19'b0001010010100001000: color_data = Z;
		19'b0001010010100001001: color_data = Z;
		19'b0001010010100001010: color_data = Z;
		19'b0001010010100001011: color_data = Z;
		19'b0001010010100001100: color_data = Z;
		19'b0001010010100001101: color_data = Z;
		19'b0001010010100001110: color_data = Z;
		19'b0001010010100001111: color_data = Z;
		19'b0001010010100010000: color_data = Z;
		19'b0001010010100010001: color_data = Z;
		19'b0001010010100010010: color_data = Z;
		19'b0001010010100010011: color_data = Z;
		19'b0001010010100010100: color_data = Z;
		19'b0001010010100010101: color_data = Z;
		19'b0001010010100010110: color_data = Z;
		19'b0001010010100010111: color_data = Z;
		19'b0001010010100011000: color_data = Z;
		19'b0001010010100011001: color_data = Z;
		19'b0001010010100011010: color_data = Z;
		19'b0001010010100011011: color_data = Z;
		19'b0001010010100011100: color_data = Z;
		19'b0001010010100011101: color_data = Z;
		19'b0001010010100011110: color_data = Z;
		19'b0001010010100011111: color_data = Z;
		19'b0001010010100100000: color_data = Z;
		19'b0001010010100100001: color_data = Z;
		19'b0001010010100100010: color_data = Z;
		19'b0001010010100100011: color_data = Z;
		19'b0001010010100100100: color_data = Z;
		19'b0001010010100100101: color_data = Z;
		19'b0001010010100100110: color_data = Z;
		19'b0001010010100100111: color_data = Z;
		19'b0001010010100101000: color_data = Z;
		19'b0001010010100101001: color_data = Z;
		19'b0001010010100101010: color_data = Z;
		19'b0001010010100101011: color_data = Z;
		19'b0001010010100101100: color_data = Z;
		19'b0001010010100101101: color_data = Z;
		19'b0001010010100101110: color_data = Z;
		19'b0001010010100101111: color_data = Z;
		19'b0001010010100110000: color_data = Z;
		19'b0001010010100110001: color_data = Z;
		19'b0001010010100110010: color_data = Z;
		19'b0001010010100110011: color_data = Z;
		19'b0001010010100110100: color_data = Z;
		19'b0001010010100110101: color_data = Z;
		19'b0001010010100110110: color_data = Z;
		19'b0001010010100110111: color_data = Z;
		19'b0001010010100111000: color_data = Z;
		19'b0001010010100111001: color_data = Z;
		19'b0001010010100111010: color_data = Z;
		19'b0001010010100111011: color_data = Z;
		19'b0001010010100111100: color_data = Z;
		19'b0001010010100111101: color_data = Z;
		19'b0001010010100111110: color_data = Z;
		19'b0001010010100111111: color_data = Z;
		19'b0001010010101000000: color_data = Z;
		19'b0001010010101000001: color_data = Z;
		19'b0001010010101000010: color_data = Z;
		19'b0001010010101000011: color_data = Z;
		19'b0001010010101000100: color_data = Z;
		19'b0001010010101000101: color_data = Z;
		19'b0001010010101000110: color_data = Z;
		19'b0001010010101000111: color_data = Z;
		19'b0001010010101001000: color_data = Z;
		19'b0001010010101001001: color_data = Z;
		19'b0001010010101001010: color_data = Z;
		19'b0001010010101001011: color_data = Z;
		19'b0001010010101001100: color_data = Z;
		19'b0001010010101001101: color_data = Z;
		19'b0001010010101001110: color_data = Z;
		19'b0001010010101001111: color_data = Z;
		19'b0001010010101010000: color_data = Z;
		19'b0001010010101010001: color_data = Z;
		19'b0001010010101010010: color_data = Z;
		19'b0001010010101010011: color_data = Z;
		19'b0001010010101010100: color_data = Z;
		19'b0001010010101010101: color_data = Z;
		19'b0001010010101010110: color_data = Z;
		19'b0001010010101010111: color_data = Z;
		19'b0001010010101011000: color_data = Z;
		19'b0001010010101011001: color_data = Z;
		19'b0001010010101011010: color_data = Z;
		19'b0001010010101011011: color_data = Z;
		19'b0001010010101011100: color_data = Z;
		19'b0001010010101011101: color_data = Z;
		19'b0001010010101011110: color_data = Z;
		19'b0001010010101011111: color_data = Z;
		19'b0001010010101100000: color_data = Z;
		19'b0001010010101100001: color_data = Z;
		19'b0001010010101100010: color_data = Z;
		19'b0001010010101100011: color_data = Z;
		19'b0001010010101100100: color_data = Z;
		19'b0001010010101100101: color_data = Z;
		19'b0001010010101100110: color_data = Z;
		19'b0001010010101100111: color_data = Z;
		19'b0001010010101101000: color_data = Z;
		19'b0001010010101101001: color_data = Z;
		19'b0001010010101101010: color_data = Z;
		19'b0001010010101101011: color_data = Z;
		19'b0001010010101101100: color_data = Z;
		19'b0001010010101101101: color_data = Z;
		19'b0001010010101101110: color_data = Z;
		19'b0001010010101101111: color_data = Z;
		19'b0001010010101110000: color_data = Z;
		19'b0001010010101110001: color_data = Z;
		19'b0001010010101110010: color_data = Z;
		19'b0001010010101110011: color_data = Z;
		19'b0001010010101110100: color_data = Z;
		19'b0001010010101110101: color_data = Z;
		19'b0001010010101110110: color_data = Z;
		19'b0001010010101110111: color_data = Z;
		19'b0001010010101111000: color_data = Z;
		19'b0001010010101111001: color_data = Z;
		19'b0001010010101111010: color_data = Z;
		19'b0001010010101111011: color_data = Z;
		19'b0001010010101111100: color_data = Z;
		19'b0001010010101111101: color_data = Z;
		19'b0001010010101111110: color_data = Z;
		19'b0001010010101111111: color_data = Z;
		19'b0001010010110000000: color_data = Z;
		19'b0001010010110000001: color_data = Z;
		19'b0001010010110000010: color_data = Z;
		19'b0001010010110000011: color_data = Z;
		19'b0001010010110000100: color_data = Z;
		19'b0001010010110000101: color_data = Z;
		19'b0001010010110000110: color_data = Z;
		19'b0001010010110000111: color_data = Z;
		19'b0001010010110001000: color_data = Z;
		19'b0001010010110001001: color_data = Z;
		19'b0001010010110001010: color_data = Z;
		19'b0001010010110001011: color_data = Z;
		19'b0001010010110001100: color_data = Z;
		19'b0001010010110001101: color_data = Z;
		19'b0001010010110001110: color_data = Z;
		19'b0001010010110001111: color_data = Z;
		19'b0001010010110010000: color_data = Z;
		19'b0001010010110010001: color_data = Z;
		19'b0001010010110010010: color_data = Z;
		19'b0001010010110010011: color_data = Z;
		19'b0001010010110010100: color_data = Z;
		19'b0001010010110010101: color_data = Z;
		19'b0001010010110010110: color_data = Z;
		19'b0001010010110010111: color_data = Z;
		19'b0001010010110011000: color_data = Z;
		19'b0001010010110011001: color_data = Z;
		19'b0001010010110011010: color_data = Z;
		19'b0001010010110011011: color_data = Z;
		19'b0001010010110100001: color_data = Z;
		19'b0001010010110100010: color_data = Z;
		19'b0001010010110100011: color_data = Z;
		19'b0001010010110100100: color_data = Z;
		19'b0001010010110100101: color_data = Z;
		19'b0001010010110100110: color_data = Z;
		19'b0001010010110100111: color_data = Z;
		19'b0001010010110101000: color_data = Z;
		19'b0001010010110101001: color_data = Z;
		19'b0001010100011100101: color_data = Z;
		19'b0001010100011100110: color_data = Z;
		19'b0001010100011100111: color_data = Z;
		19'b0001010100011101000: color_data = Z;
		19'b0001010100011101001: color_data = Z;
		19'b0001010100011101010: color_data = Z;
		19'b0001010100011101011: color_data = Z;
		19'b0001010100011101100: color_data = Z;
		19'b0001010100011101101: color_data = Z;
		19'b0001010100011101110: color_data = Z;
		19'b0001010100011101111: color_data = Z;
		19'b0001010100011110000: color_data = Z;
		19'b0001010100011110001: color_data = Z;
		19'b0001010100011110010: color_data = Z;
		19'b0001010100011110011: color_data = Z;
		19'b0001010100011110100: color_data = Z;
		19'b0001010100011110101: color_data = Z;
		19'b0001010100011110110: color_data = Z;
		19'b0001010100011110111: color_data = Z;
		19'b0001010100011111000: color_data = Z;
		19'b0001010100011111001: color_data = Z;
		19'b0001010100011111010: color_data = Z;
		19'b0001010100011111011: color_data = Z;
		19'b0001010100011111100: color_data = Z;
		19'b0001010100011111101: color_data = Z;
		19'b0001010100011111110: color_data = Z;
		19'b0001010100011111111: color_data = Z;
		19'b0001010100100000000: color_data = Z;
		19'b0001010100100000001: color_data = Z;
		19'b0001010100100000010: color_data = Z;
		19'b0001010100100000011: color_data = Z;
		19'b0001010100100000100: color_data = Z;
		19'b0001010100100000101: color_data = Z;
		19'b0001010100100000110: color_data = Z;
		19'b0001010100100000111: color_data = Z;
		19'b0001010100100001000: color_data = Z;
		19'b0001010100100001001: color_data = Z;
		19'b0001010100100001010: color_data = Z;
		19'b0001010100100001011: color_data = Z;
		19'b0001010100100001100: color_data = Z;
		19'b0001010100100001101: color_data = Z;
		19'b0001010100100001110: color_data = Z;
		19'b0001010100100001111: color_data = Z;
		19'b0001010100100010000: color_data = Z;
		19'b0001010100100010001: color_data = Z;
		19'b0001010100100010010: color_data = Z;
		19'b0001010100100010011: color_data = Z;
		19'b0001010100100010100: color_data = Z;
		19'b0001010100100010101: color_data = Z;
		19'b0001010100100010110: color_data = Z;
		19'b0001010100100010111: color_data = Z;
		19'b0001010100100011000: color_data = Z;
		19'b0001010100100011001: color_data = Z;
		19'b0001010100100011010: color_data = Z;
		19'b0001010100100011011: color_data = Z;
		19'b0001010100100011100: color_data = Z;
		19'b0001010100100011101: color_data = Z;
		19'b0001010100100011110: color_data = Z;
		19'b0001010100100011111: color_data = Z;
		19'b0001010100100100000: color_data = Z;
		19'b0001010100100100001: color_data = Z;
		19'b0001010100100100010: color_data = Z;
		19'b0001010100100100011: color_data = Z;
		19'b0001010100100100100: color_data = Z;
		19'b0001010100100100101: color_data = Z;
		19'b0001010100100100110: color_data = Z;
		19'b0001010100100100111: color_data = Z;
		19'b0001010100100101000: color_data = Z;
		19'b0001010100100101001: color_data = Z;
		19'b0001010100100101010: color_data = Z;
		19'b0001010100100101011: color_data = Z;
		19'b0001010100100101100: color_data = Z;
		19'b0001010100100101101: color_data = Z;
		19'b0001010100100101110: color_data = Z;
		19'b0001010100100101111: color_data = Z;
		19'b0001010100100110000: color_data = Z;
		19'b0001010100100110001: color_data = Z;
		19'b0001010100100110010: color_data = Z;
		19'b0001010100100110011: color_data = Z;
		19'b0001010100100110100: color_data = Z;
		19'b0001010100100110101: color_data = Z;
		19'b0001010100100110110: color_data = Z;
		19'b0001010100100110111: color_data = Z;
		19'b0001010100100111000: color_data = Z;
		19'b0001010100100111001: color_data = Z;
		19'b0001010100100111010: color_data = Z;
		19'b0001010100100111011: color_data = Z;
		19'b0001010100100111100: color_data = Z;
		19'b0001010100100111101: color_data = Z;
		19'b0001010100100111110: color_data = Z;
		19'b0001010100100111111: color_data = Z;
		19'b0001010100101000000: color_data = Z;
		19'b0001010100101000001: color_data = Z;
		19'b0001010100101000010: color_data = Z;
		19'b0001010100101000011: color_data = Z;
		19'b0001010100101000100: color_data = Z;
		19'b0001010100101000101: color_data = Z;
		19'b0001010100101000110: color_data = Z;
		19'b0001010100101000111: color_data = Z;
		19'b0001010100101001000: color_data = Z;
		19'b0001010100101001001: color_data = Z;
		19'b0001010100101001010: color_data = Z;
		19'b0001010100101001011: color_data = Z;
		19'b0001010100101001100: color_data = Z;
		19'b0001010100101001101: color_data = Z;
		19'b0001010100101001110: color_data = Z;
		19'b0001010100101001111: color_data = Z;
		19'b0001010100101010000: color_data = Z;
		19'b0001010100101010001: color_data = Z;
		19'b0001010100101010010: color_data = Z;
		19'b0001010100101010011: color_data = Z;
		19'b0001010100101010100: color_data = Z;
		19'b0001010100101010101: color_data = Z;
		19'b0001010100101010110: color_data = Z;
		19'b0001010100101010111: color_data = Z;
		19'b0001010100101011000: color_data = Z;
		19'b0001010100101011001: color_data = Z;
		19'b0001010100101011010: color_data = Z;
		19'b0001010100101011011: color_data = Z;
		19'b0001010100101011100: color_data = Z;
		19'b0001010100101011101: color_data = Z;
		19'b0001010100101011110: color_data = Z;
		19'b0001010100101011111: color_data = Z;
		19'b0001010100101100000: color_data = Z;
		19'b0001010100101100001: color_data = Z;
		19'b0001010100101100010: color_data = Z;
		19'b0001010100101100011: color_data = Z;
		19'b0001010100101100100: color_data = Z;
		19'b0001010100101100101: color_data = Z;
		19'b0001010100101100110: color_data = Z;
		19'b0001010100101100111: color_data = Z;
		19'b0001010100101101000: color_data = Z;
		19'b0001010100101101001: color_data = Z;
		19'b0001010100101101010: color_data = Z;
		19'b0001010100101101011: color_data = Z;
		19'b0001010100101101100: color_data = Z;
		19'b0001010100101101101: color_data = Z;
		19'b0001010100101101110: color_data = Z;
		19'b0001010100101101111: color_data = Z;
		19'b0001010100101110000: color_data = Z;
		19'b0001010100101110001: color_data = Z;
		19'b0001010100101110010: color_data = Z;
		19'b0001010100101110011: color_data = Z;
		19'b0001010100101110100: color_data = Z;
		19'b0001010100101110101: color_data = Z;
		19'b0001010100101110110: color_data = Z;
		19'b0001010100101110111: color_data = Z;
		19'b0001010100101111000: color_data = Z;
		19'b0001010100101111001: color_data = Z;
		19'b0001010100101111010: color_data = Z;
		19'b0001010100101111011: color_data = Z;
		19'b0001010100101111100: color_data = Z;
		19'b0001010100101111101: color_data = Z;
		19'b0001010100101111110: color_data = Z;
		19'b0001010100101111111: color_data = Z;
		19'b0001010100110000000: color_data = Z;
		19'b0001010100110000001: color_data = Z;
		19'b0001010100110000010: color_data = Z;
		19'b0001010100110000011: color_data = Z;
		19'b0001010100110000100: color_data = Z;
		19'b0001010100110000101: color_data = Z;
		19'b0001010100110000110: color_data = Z;
		19'b0001010100110000111: color_data = Z;
		19'b0001010100110001000: color_data = Z;
		19'b0001010100110001001: color_data = Z;
		19'b0001010100110001010: color_data = Z;
		19'b0001010100110001011: color_data = Z;
		19'b0001010100110001100: color_data = Z;
		19'b0001010100110001101: color_data = Z;
		19'b0001010100110001110: color_data = Z;
		19'b0001010100110001111: color_data = Z;
		19'b0001010100110010000: color_data = Z;
		19'b0001010100110010001: color_data = Z;
		19'b0001010100110010010: color_data = Z;
		19'b0001010100110010011: color_data = Z;
		19'b0001010100110010100: color_data = Z;
		19'b0001010100110010101: color_data = Z;
		19'b0001010100110010110: color_data = Z;
		19'b0001010100110010111: color_data = Z;
		19'b0001010100110011000: color_data = Z;
		19'b0001010100110011001: color_data = Z;
		19'b0001010100110011010: color_data = Z;
		19'b0001010100110011011: color_data = Z;
		19'b0001010100110100001: color_data = Z;
		19'b0001010100110100010: color_data = Z;
		19'b0001010100110100011: color_data = Z;
		19'b0001010100110100100: color_data = Z;
		19'b0001010100110100101: color_data = Z;
		19'b0001010100110100110: color_data = Z;
		19'b0001010100110101000: color_data = Z;
		19'b0001010100110101001: color_data = Z;
		19'b0001010100110101010: color_data = Z;
		19'b0001010100110101011: color_data = Z;
		19'b0001010110011100010: color_data = Z;
		19'b0001010110011100011: color_data = Z;
		19'b0001010110011100100: color_data = Z;
		19'b0001010110011100101: color_data = Z;
		19'b0001010110011100110: color_data = Z;
		19'b0001010110011100111: color_data = Z;
		19'b0001010110011101000: color_data = Z;
		19'b0001010110011101001: color_data = Z;
		19'b0001010110011101010: color_data = Z;
		19'b0001010110011101011: color_data = Z;
		19'b0001010110011101100: color_data = Z;
		19'b0001010110011101101: color_data = Z;
		19'b0001010110011101110: color_data = Z;
		19'b0001010110011101111: color_data = Z;
		19'b0001010110011110000: color_data = Z;
		19'b0001010110011110001: color_data = Z;
		19'b0001010110011110010: color_data = Z;
		19'b0001010110011110011: color_data = Z;
		19'b0001010110011110100: color_data = Z;
		19'b0001010110011110101: color_data = Z;
		19'b0001010110011110110: color_data = Z;
		19'b0001010110011110111: color_data = Z;
		19'b0001010110011111000: color_data = Z;
		19'b0001010110011111001: color_data = Z;
		19'b0001010110011111010: color_data = Z;
		19'b0001010110011111011: color_data = Z;
		19'b0001010110011111100: color_data = Z;
		19'b0001010110011111101: color_data = Z;
		19'b0001010110011111110: color_data = Z;
		19'b0001010110011111111: color_data = Z;
		19'b0001010110100000000: color_data = Z;
		19'b0001010110100000001: color_data = Z;
		19'b0001010110100000010: color_data = Z;
		19'b0001010110100000011: color_data = Z;
		19'b0001010110100000100: color_data = Z;
		19'b0001010110100000101: color_data = Z;
		19'b0001010110100000110: color_data = Z;
		19'b0001010110100000111: color_data = Z;
		19'b0001010110100001000: color_data = Z;
		19'b0001010110100001001: color_data = Z;
		19'b0001010110100001010: color_data = Z;
		19'b0001010110100001011: color_data = Z;
		19'b0001010110100001100: color_data = Z;
		19'b0001010110100001101: color_data = Z;
		19'b0001010110100001110: color_data = Z;
		19'b0001010110100001111: color_data = Z;
		19'b0001010110100010000: color_data = Z;
		19'b0001010110100010001: color_data = Z;
		19'b0001010110100010010: color_data = Z;
		19'b0001010110100010011: color_data = Z;
		19'b0001010110100010100: color_data = Z;
		19'b0001010110100010101: color_data = Z;
		19'b0001010110100010110: color_data = Z;
		19'b0001010110100010111: color_data = Z;
		19'b0001010110100011000: color_data = Z;
		19'b0001010110100011001: color_data = Z;
		19'b0001010110100011010: color_data = Z;
		19'b0001010110100011011: color_data = Z;
		19'b0001010110100011100: color_data = Z;
		19'b0001010110100011101: color_data = Z;
		19'b0001010110100011110: color_data = Z;
		19'b0001010110100011111: color_data = Z;
		19'b0001010110100100000: color_data = Z;
		19'b0001010110100100001: color_data = Z;
		19'b0001010110100100010: color_data = Z;
		19'b0001010110100100011: color_data = Z;
		19'b0001010110100100100: color_data = Z;
		19'b0001010110100100101: color_data = Z;
		19'b0001010110100100110: color_data = Z;
		19'b0001010110100100111: color_data = Z;
		19'b0001010110100101000: color_data = Z;
		19'b0001010110100101001: color_data = Z;
		19'b0001010110100101010: color_data = Z;
		19'b0001010110100101011: color_data = Z;
		19'b0001010110100101100: color_data = Z;
		19'b0001010110100101101: color_data = Z;
		19'b0001010110100101110: color_data = Z;
		19'b0001010110100101111: color_data = Z;
		19'b0001010110100110000: color_data = Z;
		19'b0001010110100110001: color_data = Z;
		19'b0001010110100110010: color_data = Z;
		19'b0001010110100110011: color_data = Z;
		19'b0001010110100110100: color_data = Z;
		19'b0001010110100110101: color_data = Z;
		19'b0001010110100110110: color_data = Z;
		19'b0001010110100110111: color_data = Z;
		19'b0001010110100111000: color_data = Z;
		19'b0001010110100111001: color_data = Z;
		19'b0001010110100111010: color_data = Z;
		19'b0001010110100111011: color_data = Z;
		19'b0001010110100111100: color_data = Z;
		19'b0001010110100111101: color_data = Z;
		19'b0001010110100111110: color_data = Z;
		19'b0001010110100111111: color_data = Z;
		19'b0001010110101000000: color_data = Z;
		19'b0001010110101000001: color_data = Z;
		19'b0001010110101000010: color_data = Z;
		19'b0001010110101000011: color_data = Z;
		19'b0001010110101000100: color_data = Z;
		19'b0001010110101000101: color_data = Z;
		19'b0001010110101000110: color_data = Z;
		19'b0001010110101000111: color_data = Z;
		19'b0001010110101001000: color_data = Z;
		19'b0001010110101001001: color_data = Z;
		19'b0001010110101001010: color_data = Z;
		19'b0001010110101001011: color_data = Z;
		19'b0001010110101001100: color_data = Z;
		19'b0001010110101001101: color_data = Z;
		19'b0001010110101001110: color_data = Z;
		19'b0001010110101001111: color_data = Z;
		19'b0001010110101010000: color_data = Z;
		19'b0001010110101010001: color_data = Z;
		19'b0001010110101010010: color_data = Z;
		19'b0001010110101010011: color_data = Z;
		19'b0001010110101010100: color_data = Z;
		19'b0001010110101010101: color_data = Z;
		19'b0001010110101010110: color_data = Z;
		19'b0001010110101010111: color_data = Z;
		19'b0001010110101011000: color_data = Z;
		19'b0001010110101011001: color_data = Z;
		19'b0001010110101011010: color_data = Z;
		19'b0001010110101011011: color_data = Z;
		19'b0001010110101011100: color_data = Z;
		19'b0001010110101011101: color_data = Z;
		19'b0001010110101011110: color_data = Z;
		19'b0001010110101011111: color_data = Z;
		19'b0001010110101100000: color_data = Z;
		19'b0001010110101100001: color_data = Z;
		19'b0001010110101100010: color_data = Z;
		19'b0001010110101100011: color_data = Z;
		19'b0001010110101100100: color_data = Z;
		19'b0001010110101100101: color_data = Z;
		19'b0001010110101100110: color_data = Z;
		19'b0001010110101100111: color_data = Z;
		19'b0001010110101101000: color_data = Z;
		19'b0001010110101101001: color_data = Z;
		19'b0001010110101101010: color_data = Z;
		19'b0001010110101101011: color_data = Z;
		19'b0001010110101101100: color_data = Z;
		19'b0001010110101101101: color_data = Z;
		19'b0001010110101101110: color_data = Z;
		19'b0001010110101101111: color_data = Z;
		19'b0001010110101110000: color_data = Z;
		19'b0001010110101110001: color_data = Z;
		19'b0001010110101110010: color_data = Z;
		19'b0001010110101110011: color_data = Z;
		19'b0001010110101110100: color_data = Z;
		19'b0001010110101110101: color_data = Z;
		19'b0001010110101110110: color_data = Z;
		19'b0001010110101110111: color_data = Z;
		19'b0001010110101111000: color_data = Z;
		19'b0001010110101111001: color_data = Z;
		19'b0001010110101111010: color_data = Z;
		19'b0001010110101111011: color_data = Z;
		19'b0001010110101111100: color_data = Z;
		19'b0001010110101111101: color_data = Z;
		19'b0001010110101111110: color_data = Z;
		19'b0001010110101111111: color_data = Z;
		19'b0001010110110000000: color_data = Z;
		19'b0001010110110000001: color_data = Z;
		19'b0001010110110000010: color_data = Z;
		19'b0001010110110000011: color_data = Z;
		19'b0001010110110000100: color_data = Z;
		19'b0001010110110000101: color_data = Z;
		19'b0001010110110000110: color_data = Z;
		19'b0001010110110000111: color_data = Z;
		19'b0001010110110001000: color_data = Z;
		19'b0001010110110001001: color_data = Z;
		19'b0001010110110001010: color_data = Z;
		19'b0001010110110001011: color_data = Z;
		19'b0001010110110001100: color_data = Z;
		19'b0001010110110001101: color_data = Z;
		19'b0001010110110001110: color_data = Z;
		19'b0001010110110001111: color_data = Z;
		19'b0001010110110010000: color_data = Z;
		19'b0001010110110010001: color_data = Z;
		19'b0001010110110010010: color_data = Z;
		19'b0001010110110010011: color_data = Z;
		19'b0001010110110010100: color_data = Z;
		19'b0001010110110010101: color_data = Z;
		19'b0001010110110010110: color_data = Z;
		19'b0001010110110010111: color_data = Z;
		19'b0001010110110011000: color_data = Z;
		19'b0001010110110011001: color_data = Z;
		19'b0001010110110011010: color_data = Z;
		19'b0001010110110011011: color_data = Z;
		19'b0001010110110011100: color_data = Z;
		19'b0001010110110100001: color_data = Z;
		19'b0001010110110100010: color_data = Z;
		19'b0001010110110100011: color_data = Z;
		19'b0001010110110100100: color_data = Z;
		19'b0001010110110100101: color_data = Z;
		19'b0001010110110100110: color_data = Z;
		19'b0001010110110101000: color_data = Z;
		19'b0001010110110101001: color_data = Z;
		19'b0001010110110101010: color_data = Z;
		19'b0001010110110101011: color_data = Z;
		19'b0001010110110101100: color_data = Z;
		19'b0001011000011100001: color_data = Z;
		19'b0001011000011100010: color_data = Z;
		19'b0001011000011100011: color_data = Z;
		19'b0001011000011100100: color_data = Z;
		19'b0001011000011100101: color_data = Z;
		19'b0001011000011100110: color_data = Z;
		19'b0001011000011100111: color_data = Z;
		19'b0001011000011101000: color_data = Z;
		19'b0001011000011101001: color_data = Z;
		19'b0001011000011101010: color_data = Z;
		19'b0001011000011101011: color_data = Z;
		19'b0001011000011101100: color_data = Z;
		19'b0001011000011101101: color_data = Z;
		19'b0001011000011101110: color_data = Z;
		19'b0001011000011101111: color_data = Z;
		19'b0001011000011110000: color_data = Z;
		19'b0001011000011110001: color_data = Z;
		19'b0001011000011110010: color_data = Z;
		19'b0001011000011110011: color_data = Z;
		19'b0001011000011110100: color_data = Z;
		19'b0001011000011110101: color_data = Z;
		19'b0001011000011110110: color_data = Z;
		19'b0001011000011110111: color_data = Z;
		19'b0001011000011111000: color_data = Z;
		19'b0001011000011111001: color_data = Z;
		19'b0001011000011111010: color_data = Z;
		19'b0001011000011111011: color_data = Z;
		19'b0001011000011111100: color_data = Z;
		19'b0001011000011111101: color_data = Z;
		19'b0001011000011111110: color_data = Z;
		19'b0001011000011111111: color_data = Z;
		19'b0001011000100000000: color_data = Z;
		19'b0001011000100000001: color_data = Z;
		19'b0001011000100000010: color_data = Z;
		19'b0001011000100000011: color_data = Z;
		19'b0001011000100000100: color_data = Z;
		19'b0001011000100000101: color_data = Z;
		19'b0001011000100000110: color_data = Z;
		19'b0001011000100000111: color_data = Z;
		19'b0001011000100001000: color_data = Z;
		19'b0001011000100001001: color_data = Z;
		19'b0001011000100001010: color_data = Z;
		19'b0001011000100001011: color_data = Z;
		19'b0001011000100001100: color_data = Z;
		19'b0001011000100001101: color_data = Z;
		19'b0001011000100001110: color_data = Z;
		19'b0001011000100001111: color_data = Z;
		19'b0001011000100010000: color_data = Z;
		19'b0001011000100010001: color_data = Z;
		19'b0001011000100010010: color_data = Z;
		19'b0001011000100010011: color_data = Z;
		19'b0001011000100010100: color_data = Z;
		19'b0001011000100010101: color_data = Z;
		19'b0001011000100010110: color_data = Z;
		19'b0001011000100010111: color_data = Z;
		19'b0001011000100011000: color_data = Z;
		19'b0001011000100011001: color_data = Z;
		19'b0001011000100011010: color_data = Z;
		19'b0001011000100011011: color_data = Z;
		19'b0001011000100011100: color_data = Z;
		19'b0001011000100011101: color_data = Z;
		19'b0001011000100011110: color_data = Z;
		19'b0001011000100011111: color_data = Z;
		19'b0001011000100100000: color_data = Z;
		19'b0001011000100100001: color_data = Z;
		19'b0001011000100100010: color_data = Z;
		19'b0001011000100100011: color_data = Z;
		19'b0001011000100100100: color_data = Z;
		19'b0001011000100100101: color_data = Z;
		19'b0001011000100100110: color_data = Z;
		19'b0001011000100100111: color_data = Z;
		19'b0001011000100101000: color_data = Z;
		19'b0001011000100101001: color_data = Z;
		19'b0001011000100101010: color_data = Z;
		19'b0001011000100101011: color_data = Z;
		19'b0001011000100101100: color_data = Z;
		19'b0001011000100101101: color_data = Z;
		19'b0001011000100101110: color_data = Z;
		19'b0001011000100101111: color_data = Z;
		19'b0001011000100110000: color_data = Z;
		19'b0001011000100110001: color_data = Z;
		19'b0001011000100110010: color_data = Z;
		19'b0001011000100110011: color_data = Z;
		19'b0001011000100110100: color_data = Z;
		19'b0001011000100110101: color_data = Z;
		19'b0001011000100110110: color_data = Z;
		19'b0001011000100110111: color_data = Z;
		19'b0001011000100111000: color_data = Z;
		19'b0001011000100111001: color_data = Z;
		19'b0001011000100111010: color_data = Z;
		19'b0001011000100111011: color_data = Z;
		19'b0001011000100111100: color_data = Z;
		19'b0001011000100111101: color_data = Z;
		19'b0001011000100111110: color_data = Z;
		19'b0001011000100111111: color_data = Z;
		19'b0001011000101000000: color_data = Z;
		19'b0001011000101000001: color_data = Z;
		19'b0001011000101000010: color_data = Z;
		19'b0001011000101000011: color_data = Z;
		19'b0001011000101000100: color_data = Z;
		19'b0001011000101000101: color_data = Z;
		19'b0001011000101000110: color_data = Z;
		19'b0001011000101000111: color_data = Z;
		19'b0001011000101001000: color_data = Z;
		19'b0001011000101001001: color_data = Z;
		19'b0001011000101001010: color_data = Z;
		19'b0001011000101001011: color_data = Z;
		19'b0001011000101001100: color_data = Z;
		19'b0001011000101001101: color_data = Z;
		19'b0001011000101001110: color_data = Z;
		19'b0001011000101001111: color_data = Z;
		19'b0001011000101010000: color_data = Z;
		19'b0001011000101010001: color_data = Z;
		19'b0001011000101010010: color_data = Z;
		19'b0001011000101010011: color_data = Z;
		19'b0001011000101010100: color_data = Z;
		19'b0001011000101010101: color_data = Z;
		19'b0001011000101010110: color_data = Z;
		19'b0001011000101010111: color_data = Z;
		19'b0001011000101011000: color_data = Z;
		19'b0001011000101011001: color_data = Z;
		19'b0001011000101011010: color_data = Z;
		19'b0001011000101011011: color_data = Z;
		19'b0001011000101011100: color_data = Z;
		19'b0001011000101011101: color_data = Z;
		19'b0001011000101011110: color_data = Z;
		19'b0001011000101011111: color_data = Z;
		19'b0001011000101100000: color_data = Z;
		19'b0001011000101100001: color_data = Z;
		19'b0001011000101100010: color_data = Z;
		19'b0001011000101100011: color_data = Z;
		19'b0001011000101100100: color_data = Z;
		19'b0001011000101100101: color_data = Z;
		19'b0001011000101100110: color_data = Z;
		19'b0001011000101100111: color_data = Z;
		19'b0001011000101101000: color_data = Z;
		19'b0001011000101101001: color_data = Z;
		19'b0001011000101101010: color_data = Z;
		19'b0001011000101101011: color_data = Z;
		19'b0001011000101101100: color_data = Z;
		19'b0001011000101101101: color_data = Z;
		19'b0001011000101101110: color_data = Z;
		19'b0001011000101101111: color_data = Z;
		19'b0001011000101110000: color_data = Z;
		19'b0001011000101110001: color_data = Z;
		19'b0001011000101110010: color_data = Z;
		19'b0001011000101110011: color_data = Z;
		19'b0001011000101110100: color_data = Z;
		19'b0001011000101110101: color_data = Z;
		19'b0001011000101110110: color_data = Z;
		19'b0001011000101110111: color_data = Z;
		19'b0001011000101111000: color_data = Z;
		19'b0001011000101111001: color_data = Z;
		19'b0001011000101111010: color_data = Z;
		19'b0001011000101111011: color_data = Z;
		19'b0001011000101111100: color_data = Z;
		19'b0001011000101111101: color_data = Z;
		19'b0001011000101111110: color_data = Z;
		19'b0001011000101111111: color_data = Z;
		19'b0001011000110000000: color_data = Z;
		19'b0001011000110000001: color_data = Z;
		19'b0001011000110000010: color_data = Z;
		19'b0001011000110000011: color_data = Z;
		19'b0001011000110000100: color_data = Z;
		19'b0001011000110000101: color_data = Z;
		19'b0001011000110000110: color_data = Z;
		19'b0001011000110000111: color_data = Z;
		19'b0001011000110001000: color_data = Z;
		19'b0001011000110001001: color_data = Z;
		19'b0001011000110001010: color_data = Z;
		19'b0001011000110001011: color_data = Z;
		19'b0001011000110001100: color_data = Z;
		19'b0001011000110001101: color_data = Z;
		19'b0001011000110001110: color_data = Z;
		19'b0001011000110001111: color_data = Z;
		19'b0001011000110010000: color_data = Z;
		19'b0001011000110010001: color_data = Z;
		19'b0001011000110010010: color_data = Z;
		19'b0001011000110010011: color_data = Z;
		19'b0001011000110010100: color_data = Z;
		19'b0001011000110010101: color_data = Z;
		19'b0001011000110010110: color_data = Z;
		19'b0001011000110010111: color_data = Z;
		19'b0001011000110011000: color_data = Z;
		19'b0001011000110011001: color_data = Z;
		19'b0001011000110011010: color_data = Z;
		19'b0001011000110011011: color_data = Z;
		19'b0001011000110011100: color_data = Z;
		19'b0001011000110100001: color_data = Z;
		19'b0001011000110100010: color_data = Z;
		19'b0001011000110100011: color_data = Z;
		19'b0001011000110100100: color_data = Z;
		19'b0001011000110100101: color_data = Z;
		19'b0001011000110101001: color_data = Z;
		19'b0001011000110101010: color_data = Z;
		19'b0001011000110101011: color_data = Z;
		19'b0001011000110101100: color_data = Z;
		19'b0001011000110101101: color_data = Z;
		19'b0001011010011100000: color_data = Z;
		19'b0001011010011100001: color_data = Z;
		19'b0001011010011100010: color_data = Z;
		19'b0001011010011100011: color_data = Z;
		19'b0001011010011100100: color_data = Z;
		19'b0001011010011100101: color_data = Z;
		19'b0001011010011100110: color_data = Z;
		19'b0001011010011100111: color_data = Z;
		19'b0001011010011101000: color_data = Z;
		19'b0001011010011101001: color_data = Z;
		19'b0001011010011101010: color_data = Z;
		19'b0001011010011101011: color_data = Z;
		19'b0001011010011101100: color_data = Z;
		19'b0001011010011101101: color_data = Z;
		19'b0001011010011101110: color_data = Z;
		19'b0001011010011101111: color_data = Z;
		19'b0001011010011110000: color_data = Z;
		19'b0001011010011110001: color_data = Z;
		19'b0001011010011110010: color_data = Z;
		19'b0001011010011110011: color_data = Z;
		19'b0001011010011110100: color_data = Z;
		19'b0001011010011110101: color_data = Z;
		19'b0001011010011110110: color_data = Z;
		19'b0001011010011110111: color_data = Z;
		19'b0001011010011111000: color_data = Z;
		19'b0001011010011111001: color_data = Z;
		19'b0001011010011111010: color_data = Z;
		19'b0001011010011111011: color_data = Z;
		19'b0001011010011111100: color_data = Z;
		19'b0001011010011111101: color_data = Z;
		19'b0001011010011111110: color_data = Z;
		19'b0001011010011111111: color_data = Z;
		19'b0001011010100000000: color_data = Z;
		19'b0001011010100000001: color_data = Z;
		19'b0001011010100000010: color_data = Z;
		19'b0001011010100000011: color_data = Z;
		19'b0001011010100000100: color_data = Z;
		19'b0001011010100000101: color_data = Z;
		19'b0001011010100000110: color_data = Z;
		19'b0001011010100000111: color_data = Z;
		19'b0001011010100001000: color_data = Z;
		19'b0001011010100001001: color_data = Z;
		19'b0001011010100001010: color_data = Z;
		19'b0001011010100001011: color_data = Z;
		19'b0001011010100001100: color_data = Z;
		19'b0001011010100001101: color_data = Z;
		19'b0001011010100001110: color_data = Z;
		19'b0001011010100001111: color_data = Z;
		19'b0001011010100010000: color_data = Z;
		19'b0001011010100010001: color_data = Z;
		19'b0001011010100010010: color_data = Z;
		19'b0001011010100010011: color_data = Z;
		19'b0001011010100010100: color_data = Z;
		19'b0001011010100010101: color_data = Z;
		19'b0001011010100010110: color_data = Z;
		19'b0001011010100010111: color_data = Z;
		19'b0001011010100011000: color_data = Z;
		19'b0001011010100011001: color_data = Z;
		19'b0001011010100011010: color_data = Z;
		19'b0001011010100011011: color_data = Z;
		19'b0001011010100011100: color_data = Z;
		19'b0001011010100011101: color_data = Z;
		19'b0001011010100011110: color_data = Z;
		19'b0001011010100011111: color_data = Z;
		19'b0001011010100100000: color_data = Z;
		19'b0001011010100100001: color_data = Z;
		19'b0001011010100100010: color_data = Z;
		19'b0001011010100100011: color_data = Z;
		19'b0001011010100100100: color_data = Z;
		19'b0001011010100100101: color_data = Z;
		19'b0001011010100100110: color_data = Z;
		19'b0001011010100100111: color_data = Z;
		19'b0001011010100101000: color_data = Z;
		19'b0001011010100101001: color_data = Z;
		19'b0001011010100101010: color_data = Z;
		19'b0001011010100101011: color_data = Z;
		19'b0001011010100101100: color_data = Z;
		19'b0001011010100101101: color_data = Z;
		19'b0001011010100101110: color_data = Z;
		19'b0001011010100101111: color_data = Z;
		19'b0001011010100110000: color_data = Z;
		19'b0001011010100110001: color_data = Z;
		19'b0001011010100110010: color_data = Z;
		19'b0001011010100110011: color_data = Z;
		19'b0001011010100110100: color_data = Z;
		19'b0001011010100110101: color_data = Z;
		19'b0001011010100110110: color_data = Z;
		19'b0001011010100110111: color_data = Z;
		19'b0001011010100111000: color_data = Z;
		19'b0001011010100111001: color_data = Z;
		19'b0001011010100111010: color_data = Z;
		19'b0001011010100111011: color_data = Z;
		19'b0001011010100111100: color_data = Z;
		19'b0001011010100111101: color_data = Z;
		19'b0001011010100111110: color_data = Z;
		19'b0001011010100111111: color_data = Z;
		19'b0001011010101000000: color_data = Z;
		19'b0001011010101000001: color_data = Z;
		19'b0001011010101000010: color_data = Z;
		19'b0001011010101000011: color_data = Z;
		19'b0001011010101000100: color_data = Z;
		19'b0001011010101000101: color_data = Z;
		19'b0001011010101000110: color_data = Z;
		19'b0001011010101000111: color_data = Z;
		19'b0001011010101001000: color_data = Z;
		19'b0001011010101001001: color_data = Z;
		19'b0001011010101001010: color_data = Z;
		19'b0001011010101001011: color_data = Z;
		19'b0001011010101001100: color_data = Z;
		19'b0001011010101001101: color_data = Z;
		19'b0001011010101001110: color_data = Z;
		19'b0001011010101001111: color_data = Z;
		19'b0001011010101010000: color_data = Z;
		19'b0001011010101010001: color_data = Z;
		19'b0001011010101010010: color_data = Z;
		19'b0001011010101010011: color_data = Z;
		19'b0001011010101010100: color_data = Z;
		19'b0001011010101010101: color_data = Z;
		19'b0001011010101010110: color_data = Z;
		19'b0001011010101010111: color_data = Z;
		19'b0001011010101011000: color_data = Z;
		19'b0001011010101011001: color_data = Z;
		19'b0001011010101011010: color_data = Z;
		19'b0001011010101011011: color_data = Z;
		19'b0001011010101011100: color_data = Z;
		19'b0001011010101011101: color_data = Z;
		19'b0001011010101011110: color_data = Z;
		19'b0001011010101011111: color_data = Z;
		19'b0001011010101100000: color_data = Z;
		19'b0001011010101100001: color_data = Z;
		19'b0001011010101100010: color_data = Z;
		19'b0001011010101100011: color_data = Z;
		19'b0001011010101100100: color_data = Z;
		19'b0001011010101100101: color_data = Z;
		19'b0001011010101100110: color_data = Z;
		19'b0001011010101100111: color_data = Z;
		19'b0001011010101101000: color_data = Z;
		19'b0001011010101101001: color_data = Z;
		19'b0001011010101101010: color_data = Z;
		19'b0001011010101101011: color_data = Z;
		19'b0001011010101101100: color_data = Z;
		19'b0001011010101101101: color_data = Z;
		19'b0001011010101101110: color_data = Z;
		19'b0001011010101101111: color_data = Z;
		19'b0001011010101110000: color_data = Z;
		19'b0001011010101110001: color_data = Z;
		19'b0001011010101110010: color_data = Z;
		19'b0001011010101110011: color_data = Z;
		19'b0001011010101110100: color_data = Z;
		19'b0001011010101110101: color_data = Z;
		19'b0001011010101110110: color_data = Z;
		19'b0001011010101110111: color_data = Z;
		19'b0001011010101111000: color_data = Z;
		19'b0001011010101111001: color_data = Z;
		19'b0001011010101111010: color_data = Z;
		19'b0001011010101111011: color_data = Z;
		19'b0001011010101111100: color_data = Z;
		19'b0001011010101111101: color_data = Z;
		19'b0001011010101111110: color_data = Z;
		19'b0001011010101111111: color_data = Z;
		19'b0001011010110000000: color_data = Z;
		19'b0001011010110000001: color_data = Z;
		19'b0001011010110000010: color_data = Z;
		19'b0001011010110000011: color_data = Z;
		19'b0001011010110000100: color_data = Z;
		19'b0001011010110000101: color_data = Z;
		19'b0001011010110000110: color_data = Z;
		19'b0001011010110000111: color_data = Z;
		19'b0001011010110001000: color_data = Z;
		19'b0001011010110001001: color_data = Z;
		19'b0001011010110001010: color_data = Z;
		19'b0001011010110001011: color_data = Z;
		19'b0001011010110001100: color_data = Z;
		19'b0001011010110001101: color_data = Z;
		19'b0001011010110001110: color_data = Z;
		19'b0001011010110001111: color_data = Z;
		19'b0001011010110010000: color_data = Z;
		19'b0001011010110010001: color_data = Z;
		19'b0001011010110010010: color_data = Z;
		19'b0001011010110010011: color_data = Z;
		19'b0001011010110010100: color_data = Z;
		19'b0001011010110010101: color_data = Z;
		19'b0001011010110010110: color_data = Z;
		19'b0001011010110010111: color_data = Z;
		19'b0001011010110011000: color_data = Z;
		19'b0001011010110011001: color_data = Z;
		19'b0001011010110011010: color_data = Z;
		19'b0001011010110011011: color_data = Z;
		19'b0001011010110011100: color_data = Z;
		19'b0001011010110100001: color_data = Z;
		19'b0001011010110100010: color_data = Z;
		19'b0001011010110100011: color_data = Z;
		19'b0001011010110100100: color_data = Z;
		19'b0001011010110100101: color_data = Z;
		19'b0001011010110101001: color_data = Z;
		19'b0001011010110101010: color_data = Z;
		19'b0001011010110101011: color_data = Z;
		19'b0001011010110101100: color_data = Z;
		19'b0001011010110101101: color_data = Z;
		19'b0001011010110101110: color_data = Z;
		19'b0001011100011100000: color_data = Z;
		19'b0001011100011100001: color_data = Z;
		19'b0001011100011100010: color_data = Z;
		19'b0001011100011100011: color_data = Z;
		19'b0001011100011100100: color_data = Z;
		19'b0001011100011100101: color_data = Z;
		19'b0001011100011100110: color_data = Z;
		19'b0001011100011100111: color_data = Z;
		19'b0001011100011101000: color_data = Z;
		19'b0001011100011101001: color_data = Z;
		19'b0001011100011101010: color_data = Z;
		19'b0001011100011101011: color_data = Z;
		19'b0001011100011101100: color_data = Z;
		19'b0001011100011101101: color_data = Z;
		19'b0001011100011101110: color_data = Z;
		19'b0001011100011101111: color_data = Z;
		19'b0001011100011110000: color_data = Z;
		19'b0001011100011110001: color_data = Z;
		19'b0001011100011110010: color_data = Z;
		19'b0001011100011110011: color_data = Z;
		19'b0001011100011110100: color_data = Z;
		19'b0001011100011110101: color_data = Z;
		19'b0001011100011110110: color_data = Z;
		19'b0001011100011110111: color_data = Z;
		19'b0001011100011111000: color_data = Z;
		19'b0001011100011111001: color_data = Z;
		19'b0001011100011111010: color_data = Z;
		19'b0001011100011111011: color_data = Z;
		19'b0001011100011111100: color_data = Z;
		19'b0001011100011111101: color_data = Z;
		19'b0001011100011111110: color_data = Z;
		19'b0001011100011111111: color_data = Z;
		19'b0001011100100000000: color_data = Z;
		19'b0001011100100000001: color_data = Z;
		19'b0001011100100000010: color_data = Z;
		19'b0001011100100000011: color_data = Z;
		19'b0001011100100000100: color_data = Z;
		19'b0001011100100000101: color_data = Z;
		19'b0001011100100000110: color_data = Z;
		19'b0001011100100000111: color_data = Z;
		19'b0001011100100001000: color_data = Z;
		19'b0001011100100001001: color_data = Z;
		19'b0001011100100001010: color_data = Z;
		19'b0001011100100001011: color_data = Z;
		19'b0001011100100001100: color_data = Z;
		19'b0001011100100001101: color_data = Z;
		19'b0001011100100001110: color_data = Z;
		19'b0001011100100001111: color_data = Z;
		19'b0001011100100010000: color_data = Z;
		19'b0001011100100010001: color_data = Z;
		19'b0001011100100010010: color_data = Z;
		19'b0001011100100010011: color_data = Z;
		19'b0001011100100010100: color_data = Z;
		19'b0001011100100010101: color_data = Z;
		19'b0001011100100010110: color_data = Z;
		19'b0001011100100010111: color_data = Z;
		19'b0001011100100011000: color_data = Z;
		19'b0001011100100011001: color_data = Z;
		19'b0001011100100011010: color_data = Z;
		19'b0001011100100011011: color_data = Z;
		19'b0001011100100011100: color_data = Z;
		19'b0001011100100011101: color_data = Z;
		19'b0001011100100011110: color_data = Z;
		19'b0001011100100011111: color_data = Z;
		19'b0001011100100100000: color_data = Z;
		19'b0001011100100100001: color_data = Z;
		19'b0001011100100100010: color_data = Z;
		19'b0001011100100100011: color_data = Z;
		19'b0001011100100100100: color_data = Z;
		19'b0001011100100100101: color_data = Z;
		19'b0001011100100100110: color_data = Z;
		19'b0001011100100100111: color_data = Z;
		19'b0001011100100101000: color_data = Z;
		19'b0001011100100101001: color_data = Z;
		19'b0001011100100101010: color_data = Z;
		19'b0001011100100101011: color_data = Z;
		19'b0001011100100101100: color_data = Z;
		19'b0001011100100101101: color_data = Z;
		19'b0001011100100101110: color_data = Z;
		19'b0001011100100101111: color_data = Z;
		19'b0001011100100110000: color_data = Z;
		19'b0001011100100110001: color_data = Z;
		19'b0001011100100110010: color_data = Z;
		19'b0001011100100110011: color_data = Z;
		19'b0001011100100110100: color_data = Z;
		19'b0001011100100110101: color_data = Z;
		19'b0001011100100110110: color_data = Z;
		19'b0001011100100110111: color_data = Z;
		19'b0001011100100111000: color_data = Z;
		19'b0001011100100111001: color_data = Z;
		19'b0001011100100111010: color_data = Z;
		19'b0001011100100111011: color_data = Z;
		19'b0001011100100111100: color_data = Z;
		19'b0001011100100111101: color_data = Z;
		19'b0001011100100111110: color_data = Z;
		19'b0001011100100111111: color_data = Z;
		19'b0001011100101000000: color_data = Z;
		19'b0001011100101000001: color_data = Z;
		19'b0001011100101000010: color_data = Z;
		19'b0001011100101000011: color_data = Z;
		19'b0001011100101000100: color_data = Z;
		19'b0001011100101000101: color_data = Z;
		19'b0001011100101000110: color_data = Z;
		19'b0001011100101000111: color_data = Z;
		19'b0001011100101001000: color_data = Z;
		19'b0001011100101001001: color_data = Z;
		19'b0001011100101001010: color_data = Z;
		19'b0001011100101001011: color_data = Z;
		19'b0001011100101001100: color_data = Z;
		19'b0001011100101001101: color_data = Z;
		19'b0001011100101001110: color_data = Z;
		19'b0001011100101001111: color_data = Z;
		19'b0001011100101010000: color_data = Z;
		19'b0001011100101010001: color_data = Z;
		19'b0001011100101010010: color_data = Z;
		19'b0001011100101010011: color_data = Z;
		19'b0001011100101010100: color_data = Z;
		19'b0001011100101010101: color_data = Z;
		19'b0001011100101010110: color_data = Z;
		19'b0001011100101010111: color_data = Z;
		19'b0001011100101011000: color_data = Z;
		19'b0001011100101011001: color_data = Z;
		19'b0001011100101011010: color_data = Z;
		19'b0001011100101011011: color_data = Z;
		19'b0001011100101011100: color_data = Z;
		19'b0001011100101011101: color_data = Z;
		19'b0001011100101011110: color_data = Z;
		19'b0001011100101011111: color_data = Z;
		19'b0001011100101100000: color_data = Z;
		19'b0001011100101100001: color_data = Z;
		19'b0001011100101100010: color_data = Z;
		19'b0001011100101100011: color_data = Z;
		19'b0001011100101100100: color_data = Z;
		19'b0001011100101100101: color_data = Z;
		19'b0001011100101100110: color_data = Z;
		19'b0001011100101100111: color_data = Z;
		19'b0001011100101101000: color_data = Z;
		19'b0001011100101101001: color_data = Z;
		19'b0001011100101101010: color_data = Z;
		19'b0001011100101101011: color_data = Z;
		19'b0001011100101101100: color_data = Z;
		19'b0001011100101101101: color_data = Z;
		19'b0001011100101101110: color_data = Z;
		19'b0001011100101101111: color_data = Z;
		19'b0001011100101110000: color_data = Z;
		19'b0001011100101110001: color_data = Z;
		19'b0001011100101110010: color_data = Z;
		19'b0001011100101110011: color_data = Z;
		19'b0001011100101110100: color_data = Z;
		19'b0001011100101110101: color_data = Z;
		19'b0001011100101110110: color_data = Z;
		19'b0001011100101110111: color_data = Z;
		19'b0001011100101111000: color_data = Z;
		19'b0001011100101111001: color_data = Z;
		19'b0001011100101111010: color_data = Z;
		19'b0001011100101111011: color_data = Z;
		19'b0001011100101111100: color_data = Z;
		19'b0001011100101111101: color_data = Z;
		19'b0001011100101111110: color_data = Z;
		19'b0001011100101111111: color_data = Z;
		19'b0001011100110000000: color_data = Z;
		19'b0001011100110000001: color_data = Z;
		19'b0001011100110000010: color_data = Z;
		19'b0001011100110000011: color_data = Z;
		19'b0001011100110000100: color_data = Z;
		19'b0001011100110000101: color_data = Z;
		19'b0001011100110000110: color_data = Z;
		19'b0001011100110000111: color_data = Z;
		19'b0001011100110001000: color_data = Z;
		19'b0001011100110001001: color_data = Z;
		19'b0001011100110001010: color_data = Z;
		19'b0001011100110001011: color_data = Z;
		19'b0001011100110001100: color_data = Z;
		19'b0001011100110001101: color_data = Z;
		19'b0001011100110001110: color_data = Z;
		19'b0001011100110001111: color_data = Z;
		19'b0001011100110010000: color_data = Z;
		19'b0001011100110010001: color_data = Z;
		19'b0001011100110010010: color_data = Z;
		19'b0001011100110010011: color_data = Z;
		19'b0001011100110010100: color_data = Z;
		19'b0001011100110010101: color_data = Z;
		19'b0001011100110010110: color_data = Z;
		19'b0001011100110010111: color_data = Z;
		19'b0001011100110011000: color_data = Z;
		19'b0001011100110011001: color_data = Z;
		19'b0001011100110011010: color_data = Z;
		19'b0001011100110011011: color_data = Z;
		19'b0001011100110011100: color_data = Z;
		19'b0001011100110100011: color_data = Z;
		19'b0001011100110100100: color_data = Z;
		19'b0001011100110100101: color_data = Z;
		19'b0001011100110101010: color_data = Z;
		19'b0001011100110101011: color_data = Z;
		19'b0001011100110101100: color_data = Z;
		19'b0001011100110101101: color_data = Z;
		19'b0001011100110101110: color_data = Z;
		19'b0001011100110101111: color_data = Z;
		19'b0001011110011011111: color_data = Z;
		19'b0001011110011100000: color_data = Z;
		19'b0001011110011100001: color_data = Z;
		19'b0001011110011100010: color_data = Z;
		19'b0001011110011100011: color_data = Z;
		19'b0001011110011100100: color_data = Z;
		19'b0001011110011100101: color_data = Z;
		19'b0001011110011100110: color_data = Z;
		19'b0001011110011100111: color_data = Z;
		19'b0001011110011101000: color_data = Z;
		19'b0001011110011101001: color_data = Z;
		19'b0001011110011101010: color_data = Z;
		19'b0001011110011101011: color_data = Z;
		19'b0001011110011101100: color_data = Z;
		19'b0001011110011101101: color_data = Z;
		19'b0001011110011101110: color_data = Z;
		19'b0001011110011101111: color_data = Z;
		19'b0001011110011110000: color_data = Z;
		19'b0001011110011110001: color_data = Z;
		19'b0001011110011110010: color_data = Z;
		19'b0001011110011110011: color_data = Z;
		19'b0001011110011110100: color_data = Z;
		19'b0001011110011110101: color_data = Z;
		19'b0001011110011110110: color_data = Z;
		19'b0001011110011110111: color_data = Z;
		19'b0001011110011111000: color_data = Z;
		19'b0001011110011111001: color_data = Z;
		19'b0001011110011111010: color_data = Z;
		19'b0001011110011111011: color_data = Z;
		19'b0001011110011111100: color_data = Z;
		19'b0001011110011111101: color_data = Z;
		19'b0001011110011111110: color_data = Z;
		19'b0001011110011111111: color_data = Z;
		19'b0001011110100000000: color_data = Z;
		19'b0001011110100000001: color_data = Z;
		19'b0001011110100000010: color_data = Z;
		19'b0001011110100000011: color_data = Z;
		19'b0001011110100000100: color_data = Z;
		19'b0001011110100000101: color_data = Z;
		19'b0001011110100000110: color_data = Z;
		19'b0001011110100000111: color_data = Z;
		19'b0001011110100001000: color_data = Z;
		19'b0001011110100001001: color_data = Z;
		19'b0001011110100001010: color_data = Z;
		19'b0001011110100001011: color_data = Z;
		19'b0001011110100001100: color_data = Z;
		19'b0001011110100001101: color_data = Z;
		19'b0001011110100001110: color_data = Z;
		19'b0001011110100001111: color_data = Z;
		19'b0001011110100010000: color_data = Z;
		19'b0001011110100010001: color_data = Z;
		19'b0001011110100010010: color_data = Z;
		19'b0001011110100010011: color_data = Z;
		19'b0001011110100010100: color_data = Z;
		19'b0001011110100010101: color_data = Z;
		19'b0001011110100010110: color_data = Z;
		19'b0001011110100010111: color_data = Z;
		19'b0001011110100011000: color_data = Z;
		19'b0001011110100011001: color_data = Z;
		19'b0001011110100011010: color_data = Z;
		19'b0001011110100011011: color_data = Z;
		19'b0001011110100011100: color_data = Z;
		19'b0001011110100011101: color_data = Z;
		19'b0001011110100011110: color_data = Z;
		19'b0001011110100011111: color_data = Z;
		19'b0001011110100100000: color_data = Z;
		19'b0001011110100100001: color_data = Z;
		19'b0001011110100100010: color_data = Z;
		19'b0001011110100100011: color_data = Z;
		19'b0001011110100100100: color_data = Z;
		19'b0001011110100100101: color_data = Z;
		19'b0001011110100100110: color_data = Z;
		19'b0001011110100100111: color_data = Z;
		19'b0001011110100101000: color_data = Z;
		19'b0001011110100101001: color_data = Z;
		19'b0001011110100101010: color_data = Z;
		19'b0001011110100101011: color_data = Z;
		19'b0001011110100101100: color_data = Z;
		19'b0001011110100101101: color_data = Z;
		19'b0001011110100101110: color_data = Z;
		19'b0001011110100101111: color_data = Z;
		19'b0001011110100110000: color_data = Z;
		19'b0001011110100110001: color_data = Z;
		19'b0001011110100110010: color_data = Z;
		19'b0001011110100110011: color_data = Z;
		19'b0001011110100110100: color_data = Z;
		19'b0001011110100110101: color_data = Z;
		19'b0001011110100110110: color_data = Z;
		19'b0001011110100110111: color_data = Z;
		19'b0001011110100111000: color_data = Z;
		19'b0001011110100111001: color_data = Z;
		19'b0001011110100111010: color_data = Z;
		19'b0001011110100111011: color_data = Z;
		19'b0001011110100111100: color_data = Z;
		19'b0001011110100111101: color_data = Z;
		19'b0001011110100111110: color_data = Z;
		19'b0001011110100111111: color_data = Z;
		19'b0001011110101000000: color_data = Z;
		19'b0001011110101000001: color_data = Z;
		19'b0001011110101000010: color_data = Z;
		19'b0001011110101000011: color_data = Z;
		19'b0001011110101000100: color_data = Z;
		19'b0001011110101000101: color_data = Z;
		19'b0001011110101000110: color_data = Z;
		19'b0001011110101000111: color_data = Z;
		19'b0001011110101001000: color_data = Z;
		19'b0001011110101001001: color_data = Z;
		19'b0001011110101001010: color_data = Z;
		19'b0001011110101001011: color_data = Z;
		19'b0001011110101001100: color_data = Z;
		19'b0001011110101001101: color_data = Z;
		19'b0001011110101001110: color_data = Z;
		19'b0001011110101001111: color_data = Z;
		19'b0001011110101010000: color_data = Z;
		19'b0001011110101010001: color_data = Z;
		19'b0001011110101010010: color_data = Z;
		19'b0001011110101010011: color_data = Z;
		19'b0001011110101010100: color_data = Z;
		19'b0001011110101010101: color_data = Z;
		19'b0001011110101010110: color_data = Z;
		19'b0001011110101010111: color_data = Z;
		19'b0001011110101011000: color_data = Z;
		19'b0001011110101011001: color_data = Z;
		19'b0001011110101011010: color_data = Z;
		19'b0001011110101011011: color_data = Z;
		19'b0001011110101011100: color_data = Z;
		19'b0001011110101011101: color_data = Z;
		19'b0001011110101011110: color_data = Z;
		19'b0001011110101011111: color_data = Z;
		19'b0001011110101100000: color_data = Z;
		19'b0001011110101100001: color_data = Z;
		19'b0001011110101100010: color_data = Z;
		19'b0001011110101100011: color_data = Z;
		19'b0001011110101100100: color_data = Z;
		19'b0001011110101100101: color_data = Z;
		19'b0001011110101100110: color_data = Z;
		19'b0001011110101100111: color_data = Z;
		19'b0001011110101101000: color_data = Z;
		19'b0001011110101101001: color_data = Z;
		19'b0001011110101101010: color_data = Z;
		19'b0001011110101101011: color_data = Z;
		19'b0001011110101101100: color_data = Z;
		19'b0001011110101101101: color_data = Z;
		19'b0001011110101101110: color_data = Z;
		19'b0001011110101101111: color_data = Z;
		19'b0001011110101110000: color_data = Z;
		19'b0001011110101110001: color_data = Z;
		19'b0001011110101110010: color_data = Z;
		19'b0001011110101110011: color_data = Z;
		19'b0001011110101110100: color_data = Z;
		19'b0001011110101110101: color_data = Z;
		19'b0001011110101110110: color_data = Z;
		19'b0001011110101110111: color_data = Z;
		19'b0001011110101111000: color_data = Z;
		19'b0001011110101111001: color_data = Z;
		19'b0001011110101111010: color_data = Z;
		19'b0001011110101111011: color_data = Z;
		19'b0001011110101111100: color_data = Z;
		19'b0001011110101111101: color_data = Z;
		19'b0001011110101111110: color_data = Z;
		19'b0001011110101111111: color_data = Z;
		19'b0001011110110000000: color_data = Z;
		19'b0001011110110000001: color_data = Z;
		19'b0001011110110000010: color_data = Z;
		19'b0001011110110000011: color_data = Z;
		19'b0001011110110000100: color_data = Z;
		19'b0001011110110000101: color_data = Z;
		19'b0001011110110000110: color_data = Z;
		19'b0001011110110000111: color_data = Z;
		19'b0001011110110001000: color_data = Z;
		19'b0001011110110001001: color_data = Z;
		19'b0001011110110001010: color_data = Z;
		19'b0001011110110001011: color_data = Z;
		19'b0001011110110001100: color_data = Z;
		19'b0001011110110001101: color_data = Z;
		19'b0001011110110001110: color_data = Z;
		19'b0001011110110001111: color_data = Z;
		19'b0001011110110010000: color_data = Z;
		19'b0001011110110010001: color_data = Z;
		19'b0001011110110010010: color_data = Z;
		19'b0001011110110010011: color_data = Z;
		19'b0001011110110010100: color_data = Z;
		19'b0001011110110010101: color_data = Z;
		19'b0001011110110010110: color_data = Z;
		19'b0001011110110010111: color_data = Z;
		19'b0001011110110011000: color_data = Z;
		19'b0001011110110011001: color_data = Z;
		19'b0001011110110011010: color_data = Z;
		19'b0001011110110011011: color_data = Z;
		19'b0001011110110011100: color_data = Z;
		19'b0001011110110100011: color_data = Z;
		19'b0001011110110100100: color_data = Z;
		19'b0001011110110100101: color_data = Z;
		19'b0001011110110100110: color_data = Z;
		19'b0001011110110101010: color_data = Z;
		19'b0001011110110101011: color_data = Z;
		19'b0001011110110101100: color_data = Z;
		19'b0001011110110101101: color_data = Z;
		19'b0001011110110101110: color_data = Z;
		19'b0001011110110101111: color_data = Z;
		19'b0001011110110110000: color_data = Z;
		19'b0001100000011011110: color_data = Z;
		19'b0001100000011011111: color_data = Z;
		19'b0001100000011100000: color_data = Z;
		19'b0001100000011100001: color_data = Z;
		19'b0001100000011100010: color_data = Z;
		19'b0001100000011100011: color_data = Z;
		19'b0001100000011100100: color_data = Z;
		19'b0001100000011100101: color_data = Z;
		19'b0001100000011100110: color_data = Z;
		19'b0001100000011100111: color_data = Z;
		19'b0001100000011101000: color_data = Z;
		19'b0001100000011101001: color_data = Z;
		19'b0001100000011101010: color_data = Z;
		19'b0001100000011101011: color_data = Z;
		19'b0001100000011101100: color_data = Z;
		19'b0001100000011101101: color_data = Z;
		19'b0001100000011101110: color_data = Z;
		19'b0001100000011101111: color_data = Z;
		19'b0001100000011110000: color_data = Z;
		19'b0001100000011110001: color_data = Z;
		19'b0001100000011110010: color_data = Z;
		19'b0001100000011110011: color_data = Z;
		19'b0001100000011110100: color_data = Z;
		19'b0001100000011110101: color_data = Z;
		19'b0001100000011110110: color_data = Z;
		19'b0001100000011110111: color_data = Z;
		19'b0001100000011111000: color_data = Z;
		19'b0001100000011111001: color_data = Z;
		19'b0001100000011111010: color_data = Z;
		19'b0001100000011111011: color_data = Z;
		19'b0001100000011111100: color_data = Z;
		19'b0001100000011111101: color_data = Z;
		19'b0001100000011111110: color_data = Z;
		19'b0001100000011111111: color_data = Z;
		19'b0001100000100000000: color_data = Z;
		19'b0001100000100000001: color_data = Z;
		19'b0001100000100000010: color_data = Z;
		19'b0001100000100000011: color_data = Z;
		19'b0001100000100000100: color_data = Z;
		19'b0001100000100000101: color_data = Z;
		19'b0001100000100000110: color_data = Z;
		19'b0001100000100000111: color_data = Z;
		19'b0001100000100001000: color_data = Z;
		19'b0001100000100001001: color_data = Z;
		19'b0001100000100001010: color_data = Z;
		19'b0001100000100001011: color_data = Z;
		19'b0001100000100001100: color_data = Z;
		19'b0001100000100001101: color_data = Z;
		19'b0001100000100001110: color_data = Z;
		19'b0001100000100001111: color_data = Z;
		19'b0001100000100010000: color_data = Z;
		19'b0001100000100010001: color_data = Z;
		19'b0001100000100010010: color_data = Z;
		19'b0001100000100010011: color_data = Z;
		19'b0001100000100010100: color_data = Z;
		19'b0001100000100010101: color_data = Z;
		19'b0001100000100010110: color_data = Z;
		19'b0001100000100010111: color_data = Z;
		19'b0001100000100011000: color_data = Z;
		19'b0001100000100011001: color_data = Z;
		19'b0001100000100011010: color_data = Z;
		19'b0001100000100011011: color_data = Z;
		19'b0001100000100011100: color_data = Z;
		19'b0001100000100011101: color_data = Z;
		19'b0001100000100011110: color_data = Z;
		19'b0001100000100011111: color_data = Z;
		19'b0001100000100100000: color_data = Z;
		19'b0001100000100100001: color_data = Z;
		19'b0001100000100100010: color_data = Z;
		19'b0001100000100100011: color_data = Z;
		19'b0001100000100100100: color_data = Z;
		19'b0001100000100100101: color_data = Z;
		19'b0001100000100100110: color_data = Z;
		19'b0001100000100100111: color_data = Z;
		19'b0001100000100101000: color_data = Z;
		19'b0001100000100101001: color_data = Z;
		19'b0001100000100101010: color_data = Z;
		19'b0001100000100101011: color_data = Z;
		19'b0001100000100101100: color_data = Z;
		19'b0001100000100101101: color_data = Z;
		19'b0001100000100101110: color_data = Z;
		19'b0001100000100101111: color_data = Z;
		19'b0001100000100110000: color_data = Z;
		19'b0001100000100110001: color_data = Z;
		19'b0001100000100110010: color_data = Z;
		19'b0001100000100110011: color_data = Z;
		19'b0001100000100110100: color_data = Z;
		19'b0001100000100110101: color_data = Z;
		19'b0001100000100110110: color_data = Z;
		19'b0001100000100110111: color_data = Z;
		19'b0001100000100111000: color_data = Z;
		19'b0001100000100111001: color_data = Z;
		19'b0001100000100111010: color_data = Z;
		19'b0001100000100111011: color_data = Z;
		19'b0001100000100111100: color_data = Z;
		19'b0001100000100111101: color_data = Z;
		19'b0001100000100111110: color_data = Z;
		19'b0001100000100111111: color_data = Z;
		19'b0001100000101000000: color_data = Z;
		19'b0001100000101000001: color_data = Z;
		19'b0001100000101000010: color_data = Z;
		19'b0001100000101000011: color_data = Z;
		19'b0001100000101000100: color_data = Z;
		19'b0001100000101000101: color_data = Z;
		19'b0001100000101000110: color_data = Z;
		19'b0001100000101000111: color_data = Z;
		19'b0001100000101001000: color_data = Z;
		19'b0001100000101001001: color_data = Z;
		19'b0001100000101001010: color_data = Z;
		19'b0001100000101001011: color_data = Z;
		19'b0001100000101001100: color_data = Z;
		19'b0001100000101001101: color_data = Z;
		19'b0001100000101001110: color_data = Z;
		19'b0001100000101001111: color_data = Z;
		19'b0001100000101010000: color_data = Z;
		19'b0001100000101010001: color_data = Z;
		19'b0001100000101010010: color_data = Z;
		19'b0001100000101010011: color_data = Z;
		19'b0001100000101010100: color_data = Z;
		19'b0001100000101010101: color_data = Z;
		19'b0001100000101010110: color_data = Z;
		19'b0001100000101010111: color_data = Z;
		19'b0001100000101011000: color_data = Z;
		19'b0001100000101011001: color_data = Z;
		19'b0001100000101011010: color_data = Z;
		19'b0001100000101011011: color_data = Z;
		19'b0001100000101011100: color_data = Z;
		19'b0001100000101011101: color_data = Z;
		19'b0001100000101011110: color_data = Z;
		19'b0001100000101011111: color_data = Z;
		19'b0001100000101100000: color_data = Z;
		19'b0001100000101100001: color_data = Z;
		19'b0001100000101100010: color_data = Z;
		19'b0001100000101100011: color_data = Z;
		19'b0001100000101100100: color_data = Z;
		19'b0001100000101100101: color_data = Z;
		19'b0001100000101100110: color_data = Z;
		19'b0001100000101100111: color_data = Z;
		19'b0001100000101101000: color_data = Z;
		19'b0001100000101101001: color_data = Z;
		19'b0001100000101101010: color_data = Z;
		19'b0001100000101101011: color_data = Z;
		19'b0001100000101101100: color_data = Z;
		19'b0001100000101101101: color_data = Z;
		19'b0001100000101101110: color_data = Z;
		19'b0001100000101101111: color_data = Z;
		19'b0001100000101110000: color_data = Z;
		19'b0001100000101110001: color_data = Z;
		19'b0001100000101110010: color_data = Z;
		19'b0001100000101110011: color_data = Z;
		19'b0001100000101110100: color_data = Z;
		19'b0001100000101110101: color_data = Z;
		19'b0001100000101110110: color_data = Z;
		19'b0001100000101110111: color_data = Z;
		19'b0001100000101111000: color_data = Z;
		19'b0001100000101111001: color_data = Z;
		19'b0001100000101111010: color_data = Z;
		19'b0001100000101111011: color_data = Z;
		19'b0001100000101111100: color_data = Z;
		19'b0001100000101111101: color_data = Z;
		19'b0001100000101111110: color_data = Z;
		19'b0001100000101111111: color_data = Z;
		19'b0001100000110000000: color_data = Z;
		19'b0001100000110000001: color_data = Z;
		19'b0001100000110000010: color_data = Z;
		19'b0001100000110000011: color_data = Z;
		19'b0001100000110000100: color_data = Z;
		19'b0001100000110000101: color_data = Z;
		19'b0001100000110000110: color_data = Z;
		19'b0001100000110000111: color_data = Z;
		19'b0001100000110001000: color_data = Z;
		19'b0001100000110001001: color_data = Z;
		19'b0001100000110001010: color_data = Z;
		19'b0001100000110001011: color_data = Z;
		19'b0001100000110001100: color_data = Z;
		19'b0001100000110001101: color_data = Z;
		19'b0001100000110001110: color_data = Z;
		19'b0001100000110001111: color_data = Z;
		19'b0001100000110010000: color_data = Z;
		19'b0001100000110010001: color_data = Z;
		19'b0001100000110010010: color_data = Z;
		19'b0001100000110010011: color_data = Z;
		19'b0001100000110010100: color_data = Z;
		19'b0001100000110010101: color_data = Z;
		19'b0001100000110010110: color_data = Z;
		19'b0001100000110010111: color_data = Z;
		19'b0001100000110011000: color_data = Z;
		19'b0001100000110011001: color_data = Z;
		19'b0001100000110011010: color_data = Z;
		19'b0001100000110011011: color_data = Z;
		19'b0001100000110011100: color_data = Z;
		19'b0001100000110100010: color_data = Z;
		19'b0001100000110100011: color_data = Z;
		19'b0001100000110100100: color_data = Z;
		19'b0001100000110100101: color_data = Z;
		19'b0001100000110100110: color_data = Z;
		19'b0001100000110100111: color_data = Z;
		19'b0001100000110101100: color_data = Z;
		19'b0001100000110101101: color_data = Z;
		19'b0001100000110101110: color_data = Z;
		19'b0001100000110101111: color_data = Z;
		19'b0001100000110110000: color_data = Z;
		19'b0001100000110110001: color_data = Z;
		19'b0001100010011011101: color_data = Z;
		19'b0001100010011011110: color_data = Z;
		19'b0001100010011011111: color_data = Z;
		19'b0001100010011100000: color_data = Z;
		19'b0001100010011100001: color_data = Z;
		19'b0001100010011100010: color_data = Z;
		19'b0001100010011100011: color_data = Z;
		19'b0001100010011100100: color_data = Z;
		19'b0001100010011100101: color_data = Z;
		19'b0001100010011100110: color_data = Z;
		19'b0001100010011100111: color_data = Z;
		19'b0001100010011101000: color_data = Z;
		19'b0001100010011101001: color_data = Z;
		19'b0001100010011101010: color_data = Z;
		19'b0001100010011101011: color_data = Z;
		19'b0001100010011101100: color_data = Z;
		19'b0001100010011101101: color_data = Z;
		19'b0001100010011101110: color_data = Z;
		19'b0001100010011101111: color_data = Z;
		19'b0001100010011110000: color_data = Z;
		19'b0001100010011110001: color_data = Z;
		19'b0001100010011110010: color_data = Z;
		19'b0001100010011110011: color_data = Z;
		19'b0001100010011110100: color_data = Z;
		19'b0001100010011110101: color_data = Z;
		19'b0001100010011110110: color_data = Z;
		19'b0001100010011110111: color_data = Z;
		19'b0001100010011111000: color_data = Z;
		19'b0001100010011111001: color_data = Z;
		19'b0001100010011111010: color_data = Z;
		19'b0001100010011111011: color_data = Z;
		19'b0001100010011111100: color_data = Z;
		19'b0001100010011111101: color_data = Z;
		19'b0001100010011111110: color_data = Z;
		19'b0001100010011111111: color_data = Z;
		19'b0001100010100000000: color_data = Z;
		19'b0001100010100000001: color_data = Z;
		19'b0001100010100000010: color_data = Z;
		19'b0001100010100000011: color_data = Z;
		19'b0001100010100000100: color_data = Z;
		19'b0001100010100000101: color_data = Z;
		19'b0001100010100000110: color_data = Z;
		19'b0001100010100000111: color_data = Z;
		19'b0001100010100001000: color_data = Z;
		19'b0001100010100001001: color_data = Z;
		19'b0001100010100001010: color_data = Z;
		19'b0001100010100001011: color_data = Z;
		19'b0001100010100001100: color_data = Z;
		19'b0001100010100001101: color_data = Z;
		19'b0001100010100001110: color_data = Z;
		19'b0001100010100001111: color_data = Z;
		19'b0001100010100010000: color_data = Z;
		19'b0001100010100010001: color_data = Z;
		19'b0001100010100010010: color_data = Z;
		19'b0001100010100010011: color_data = Z;
		19'b0001100010100010100: color_data = Z;
		19'b0001100010100010101: color_data = Z;
		19'b0001100010100010110: color_data = Z;
		19'b0001100010100010111: color_data = Z;
		19'b0001100010100011000: color_data = Z;
		19'b0001100010100011001: color_data = Z;
		19'b0001100010100011010: color_data = Z;
		19'b0001100010100011011: color_data = Z;
		19'b0001100010100011100: color_data = Z;
		19'b0001100010100011101: color_data = Z;
		19'b0001100010100011110: color_data = Z;
		19'b0001100010100011111: color_data = Z;
		19'b0001100010100100000: color_data = Z;
		19'b0001100010100100001: color_data = Z;
		19'b0001100010100100010: color_data = Z;
		19'b0001100010100100011: color_data = Z;
		19'b0001100010100100100: color_data = Z;
		19'b0001100010100100101: color_data = Z;
		19'b0001100010100100110: color_data = Z;
		19'b0001100010100100111: color_data = Z;
		19'b0001100010100101000: color_data = Z;
		19'b0001100010100101001: color_data = Z;
		19'b0001100010100101010: color_data = Z;
		19'b0001100010100101011: color_data = Z;
		19'b0001100010100101100: color_data = Z;
		19'b0001100010100101101: color_data = Z;
		19'b0001100010100101110: color_data = Z;
		19'b0001100010100101111: color_data = Z;
		19'b0001100010100110000: color_data = Z;
		19'b0001100010100110001: color_data = Z;
		19'b0001100010100110010: color_data = Z;
		19'b0001100010100110011: color_data = Z;
		19'b0001100010100110100: color_data = Z;
		19'b0001100010100110101: color_data = Z;
		19'b0001100010100110110: color_data = Z;
		19'b0001100010100110111: color_data = Z;
		19'b0001100010100111000: color_data = Z;
		19'b0001100010100111001: color_data = Z;
		19'b0001100010100111010: color_data = Z;
		19'b0001100010100111011: color_data = Z;
		19'b0001100010100111100: color_data = Z;
		19'b0001100010100111101: color_data = Z;
		19'b0001100010100111110: color_data = Z;
		19'b0001100010100111111: color_data = Z;
		19'b0001100010101000000: color_data = Z;
		19'b0001100010101000001: color_data = Z;
		19'b0001100010101000010: color_data = Z;
		19'b0001100010101000011: color_data = Z;
		19'b0001100010101000100: color_data = Z;
		19'b0001100010101000101: color_data = Z;
		19'b0001100010101000110: color_data = Z;
		19'b0001100010101000111: color_data = Z;
		19'b0001100010101001000: color_data = Z;
		19'b0001100010101001001: color_data = Z;
		19'b0001100010101001010: color_data = Z;
		19'b0001100010101001011: color_data = Z;
		19'b0001100010101001100: color_data = Z;
		19'b0001100010101001101: color_data = Z;
		19'b0001100010101001110: color_data = Z;
		19'b0001100010101001111: color_data = Z;
		19'b0001100010101010000: color_data = Z;
		19'b0001100010101010001: color_data = Z;
		19'b0001100010101010010: color_data = Z;
		19'b0001100010101010011: color_data = Z;
		19'b0001100010101010100: color_data = Z;
		19'b0001100010101010101: color_data = Z;
		19'b0001100010101010110: color_data = Z;
		19'b0001100010101010111: color_data = Z;
		19'b0001100010101011000: color_data = Z;
		19'b0001100010101011001: color_data = Z;
		19'b0001100010101011010: color_data = Z;
		19'b0001100010101011011: color_data = Z;
		19'b0001100010101011100: color_data = Z;
		19'b0001100010101011101: color_data = Z;
		19'b0001100010101011110: color_data = Z;
		19'b0001100010101011111: color_data = Z;
		19'b0001100010101100000: color_data = Z;
		19'b0001100010101100001: color_data = Z;
		19'b0001100010101100010: color_data = Z;
		19'b0001100010101100011: color_data = Z;
		19'b0001100010101100100: color_data = Z;
		19'b0001100010101100101: color_data = Z;
		19'b0001100010101100110: color_data = Z;
		19'b0001100010101100111: color_data = Z;
		19'b0001100010101101000: color_data = Z;
		19'b0001100010101101001: color_data = Z;
		19'b0001100010101101010: color_data = Z;
		19'b0001100010101101011: color_data = Z;
		19'b0001100010101101100: color_data = Z;
		19'b0001100010101101101: color_data = Z;
		19'b0001100010101101110: color_data = Z;
		19'b0001100010101101111: color_data = Z;
		19'b0001100010101110000: color_data = Z;
		19'b0001100010101110001: color_data = Z;
		19'b0001100010101110010: color_data = Z;
		19'b0001100010101110011: color_data = Z;
		19'b0001100010101110100: color_data = Z;
		19'b0001100010101110101: color_data = Z;
		19'b0001100010101110110: color_data = Z;
		19'b0001100010101110111: color_data = Z;
		19'b0001100010101111000: color_data = Z;
		19'b0001100010101111001: color_data = Z;
		19'b0001100010101111010: color_data = Z;
		19'b0001100010101111011: color_data = Z;
		19'b0001100010101111100: color_data = Z;
		19'b0001100010101111101: color_data = Z;
		19'b0001100010101111110: color_data = Z;
		19'b0001100010101111111: color_data = Z;
		19'b0001100010110000000: color_data = Z;
		19'b0001100010110000001: color_data = Z;
		19'b0001100010110000010: color_data = Z;
		19'b0001100010110000011: color_data = Z;
		19'b0001100010110000100: color_data = Z;
		19'b0001100010110000101: color_data = Z;
		19'b0001100010110000110: color_data = Z;
		19'b0001100010110000111: color_data = Z;
		19'b0001100010110001000: color_data = Z;
		19'b0001100010110001001: color_data = Z;
		19'b0001100010110001010: color_data = Z;
		19'b0001100010110001011: color_data = Z;
		19'b0001100010110001100: color_data = Z;
		19'b0001100010110001101: color_data = Z;
		19'b0001100010110001110: color_data = Z;
		19'b0001100010110001111: color_data = Z;
		19'b0001100010110010000: color_data = Z;
		19'b0001100010110010001: color_data = Z;
		19'b0001100010110010010: color_data = Z;
		19'b0001100010110010011: color_data = Z;
		19'b0001100010110010100: color_data = Z;
		19'b0001100010110010101: color_data = Z;
		19'b0001100010110010110: color_data = Z;
		19'b0001100010110010111: color_data = Z;
		19'b0001100010110011000: color_data = Z;
		19'b0001100010110011001: color_data = Z;
		19'b0001100010110011010: color_data = Z;
		19'b0001100010110011011: color_data = Z;
		19'b0001100010110011100: color_data = Z;
		19'b0001100010110011101: color_data = Z;
		19'b0001100010110100010: color_data = Z;
		19'b0001100010110100011: color_data = Z;
		19'b0001100010110100100: color_data = Z;
		19'b0001100010110100101: color_data = Z;
		19'b0001100010110100110: color_data = Z;
		19'b0001100010110100111: color_data = Z;
		19'b0001100010110101101: color_data = Z;
		19'b0001100010110101110: color_data = Z;
		19'b0001100010110101111: color_data = Z;
		19'b0001100010110110000: color_data = Z;
		19'b0001100010110110001: color_data = Z;
		19'b0001100010110110010: color_data = Z;
		19'b0001100100011011100: color_data = Z;
		19'b0001100100011011101: color_data = Z;
		19'b0001100100011011110: color_data = Z;
		19'b0001100100011011111: color_data = Z;
		19'b0001100100011100000: color_data = Z;
		19'b0001100100011100001: color_data = Z;
		19'b0001100100011100010: color_data = Z;
		19'b0001100100011100011: color_data = Z;
		19'b0001100100011100100: color_data = Z;
		19'b0001100100011100101: color_data = Z;
		19'b0001100100011100110: color_data = Z;
		19'b0001100100011100111: color_data = Z;
		19'b0001100100011101000: color_data = Z;
		19'b0001100100011101001: color_data = Z;
		19'b0001100100011101010: color_data = Z;
		19'b0001100100011101011: color_data = Z;
		19'b0001100100011101100: color_data = Z;
		19'b0001100100011101101: color_data = Z;
		19'b0001100100011101110: color_data = Z;
		19'b0001100100011101111: color_data = Z;
		19'b0001100100011110000: color_data = Z;
		19'b0001100100011110001: color_data = Z;
		19'b0001100100011110010: color_data = Z;
		19'b0001100100011110011: color_data = Z;
		19'b0001100100011110100: color_data = Z;
		19'b0001100100011110101: color_data = Z;
		19'b0001100100011110110: color_data = Z;
		19'b0001100100011110111: color_data = Z;
		19'b0001100100011111000: color_data = Z;
		19'b0001100100011111001: color_data = Z;
		19'b0001100100011111010: color_data = Z;
		19'b0001100100011111011: color_data = Z;
		19'b0001100100011111100: color_data = Z;
		19'b0001100100011111101: color_data = Z;
		19'b0001100100011111110: color_data = Z;
		19'b0001100100011111111: color_data = Z;
		19'b0001100100100000000: color_data = Z;
		19'b0001100100100000001: color_data = Z;
		19'b0001100100100000010: color_data = Z;
		19'b0001100100100000011: color_data = Z;
		19'b0001100100100000100: color_data = Z;
		19'b0001100100100000101: color_data = Z;
		19'b0001100100100000110: color_data = Z;
		19'b0001100100100000111: color_data = Z;
		19'b0001100100100001000: color_data = Z;
		19'b0001100100100001001: color_data = Z;
		19'b0001100100100001010: color_data = Z;
		19'b0001100100100001011: color_data = Z;
		19'b0001100100100001100: color_data = Z;
		19'b0001100100100001101: color_data = Z;
		19'b0001100100100001110: color_data = Z;
		19'b0001100100100001111: color_data = Z;
		19'b0001100100100010000: color_data = Z;
		19'b0001100100100010001: color_data = Z;
		19'b0001100100100010010: color_data = Z;
		19'b0001100100100010011: color_data = Z;
		19'b0001100100100010100: color_data = Z;
		19'b0001100100100010101: color_data = Z;
		19'b0001100100100010110: color_data = Z;
		19'b0001100100100010111: color_data = Z;
		19'b0001100100100011000: color_data = Z;
		19'b0001100100100011001: color_data = Z;
		19'b0001100100100011010: color_data = Z;
		19'b0001100100100011011: color_data = Z;
		19'b0001100100100011100: color_data = Z;
		19'b0001100100100011101: color_data = Z;
		19'b0001100100100011110: color_data = Z;
		19'b0001100100100011111: color_data = Z;
		19'b0001100100100100000: color_data = Z;
		19'b0001100100100100001: color_data = Z;
		19'b0001100100100100010: color_data = Z;
		19'b0001100100100100011: color_data = Z;
		19'b0001100100100100100: color_data = Z;
		19'b0001100100100100101: color_data = Z;
		19'b0001100100100100110: color_data = Z;
		19'b0001100100100100111: color_data = Z;
		19'b0001100100100101000: color_data = Z;
		19'b0001100100100101001: color_data = Z;
		19'b0001100100100101010: color_data = Z;
		19'b0001100100100101011: color_data = Z;
		19'b0001100100100101100: color_data = Z;
		19'b0001100100100101101: color_data = Z;
		19'b0001100100100101110: color_data = Z;
		19'b0001100100100101111: color_data = Z;
		19'b0001100100100110000: color_data = Z;
		19'b0001100100100110001: color_data = Z;
		19'b0001100100100110010: color_data = Z;
		19'b0001100100100110011: color_data = Z;
		19'b0001100100100110100: color_data = Z;
		19'b0001100100100110101: color_data = Z;
		19'b0001100100100110110: color_data = Z;
		19'b0001100100100110111: color_data = Z;
		19'b0001100100100111000: color_data = Z;
		19'b0001100100100111001: color_data = Z;
		19'b0001100100100111010: color_data = Z;
		19'b0001100100100111011: color_data = Z;
		19'b0001100100100111100: color_data = Z;
		19'b0001100100100111101: color_data = Z;
		19'b0001100100100111110: color_data = Z;
		19'b0001100100100111111: color_data = Z;
		19'b0001100100101000000: color_data = Z;
		19'b0001100100101000001: color_data = Z;
		19'b0001100100101000010: color_data = Z;
		19'b0001100100101000011: color_data = Z;
		19'b0001100100101000100: color_data = Z;
		19'b0001100100101000101: color_data = Z;
		19'b0001100100101000110: color_data = Z;
		19'b0001100100101000111: color_data = Z;
		19'b0001100100101001000: color_data = Z;
		19'b0001100100101001001: color_data = Z;
		19'b0001100100101001010: color_data = Z;
		19'b0001100100101001011: color_data = Z;
		19'b0001100100101001100: color_data = Z;
		19'b0001100100101001101: color_data = Z;
		19'b0001100100101001110: color_data = Z;
		19'b0001100100101001111: color_data = Z;
		19'b0001100100101010000: color_data = Z;
		19'b0001100100101010001: color_data = Z;
		19'b0001100100101010010: color_data = Z;
		19'b0001100100101010011: color_data = Z;
		19'b0001100100101010100: color_data = Z;
		19'b0001100100101010101: color_data = Z;
		19'b0001100100101010110: color_data = Z;
		19'b0001100100101010111: color_data = Z;
		19'b0001100100101011000: color_data = Z;
		19'b0001100100101011001: color_data = Z;
		19'b0001100100101011010: color_data = Z;
		19'b0001100100101011011: color_data = Z;
		19'b0001100100101011100: color_data = Z;
		19'b0001100100101011101: color_data = Z;
		19'b0001100100101011110: color_data = Z;
		19'b0001100100101011111: color_data = Z;
		19'b0001100100101100000: color_data = Z;
		19'b0001100100101100001: color_data = Z;
		19'b0001100100101100010: color_data = Z;
		19'b0001100100101100011: color_data = Z;
		19'b0001100100101100100: color_data = Z;
		19'b0001100100101100101: color_data = Z;
		19'b0001100100101100110: color_data = Z;
		19'b0001100100101100111: color_data = Z;
		19'b0001100100101101000: color_data = Z;
		19'b0001100100101101001: color_data = Z;
		19'b0001100100101101010: color_data = Z;
		19'b0001100100101101011: color_data = Z;
		19'b0001100100101101100: color_data = Z;
		19'b0001100100101101101: color_data = Z;
		19'b0001100100101101110: color_data = Z;
		19'b0001100100101101111: color_data = Z;
		19'b0001100100101110000: color_data = Z;
		19'b0001100100101110001: color_data = Z;
		19'b0001100100101110010: color_data = Z;
		19'b0001100100101110011: color_data = Z;
		19'b0001100100101110100: color_data = Z;
		19'b0001100100101110101: color_data = Z;
		19'b0001100100101110110: color_data = Z;
		19'b0001100100101110111: color_data = Z;
		19'b0001100100101111000: color_data = Z;
		19'b0001100100101111001: color_data = Z;
		19'b0001100100101111010: color_data = Z;
		19'b0001100100101111011: color_data = Z;
		19'b0001100100101111100: color_data = Z;
		19'b0001100100101111101: color_data = Z;
		19'b0001100100101111110: color_data = Z;
		19'b0001100100101111111: color_data = Z;
		19'b0001100100110000000: color_data = Z;
		19'b0001100100110000001: color_data = Z;
		19'b0001100100110000010: color_data = Z;
		19'b0001100100110000011: color_data = Z;
		19'b0001100100110000100: color_data = Z;
		19'b0001100100110000101: color_data = Z;
		19'b0001100100110000110: color_data = Z;
		19'b0001100100110000111: color_data = Z;
		19'b0001100100110001000: color_data = Z;
		19'b0001100100110001001: color_data = Z;
		19'b0001100100110001010: color_data = Z;
		19'b0001100100110001011: color_data = Z;
		19'b0001100100110001100: color_data = Z;
		19'b0001100100110001101: color_data = Z;
		19'b0001100100110001110: color_data = Z;
		19'b0001100100110001111: color_data = Z;
		19'b0001100100110010000: color_data = Z;
		19'b0001100100110010001: color_data = Z;
		19'b0001100100110010010: color_data = Z;
		19'b0001100100110010011: color_data = Z;
		19'b0001100100110010100: color_data = Z;
		19'b0001100100110010101: color_data = Z;
		19'b0001100100110010110: color_data = Z;
		19'b0001100100110010111: color_data = Z;
		19'b0001100100110011000: color_data = Z;
		19'b0001100100110011001: color_data = Z;
		19'b0001100100110011010: color_data = Z;
		19'b0001100100110011011: color_data = Z;
		19'b0001100100110011100: color_data = Z;
		19'b0001100100110011101: color_data = Z;
		19'b0001100100110100011: color_data = Z;
		19'b0001100100110100100: color_data = Z;
		19'b0001100100110100101: color_data = Z;
		19'b0001100100110100110: color_data = Z;
		19'b0001100100110100111: color_data = Z;
		19'b0001100100110101000: color_data = Z;
		19'b0001100100110101110: color_data = Z;
		19'b0001100100110101111: color_data = Z;
		19'b0001100100110110000: color_data = Z;
		19'b0001100100110110001: color_data = Z;
		19'b0001100100110110010: color_data = Z;
		19'b0001100100110110011: color_data = Z;
		19'b0001100110011011011: color_data = Z;
		19'b0001100110011011100: color_data = Z;
		19'b0001100110011011101: color_data = Z;
		19'b0001100110011011110: color_data = Z;
		19'b0001100110011011111: color_data = Z;
		19'b0001100110011100000: color_data = Z;
		19'b0001100110011100001: color_data = Z;
		19'b0001100110011100010: color_data = Z;
		19'b0001100110011100011: color_data = Z;
		19'b0001100110011100100: color_data = Z;
		19'b0001100110011100101: color_data = Z;
		19'b0001100110011100110: color_data = Z;
		19'b0001100110011100111: color_data = Z;
		19'b0001100110011101000: color_data = Z;
		19'b0001100110011101001: color_data = Z;
		19'b0001100110011101010: color_data = Z;
		19'b0001100110011101011: color_data = Z;
		19'b0001100110011101100: color_data = Z;
		19'b0001100110011101101: color_data = Z;
		19'b0001100110011101110: color_data = Z;
		19'b0001100110011101111: color_data = Z;
		19'b0001100110011110000: color_data = Z;
		19'b0001100110011110001: color_data = Z;
		19'b0001100110011110010: color_data = Z;
		19'b0001100110011110011: color_data = Z;
		19'b0001100110011110100: color_data = Z;
		19'b0001100110011110101: color_data = Z;
		19'b0001100110011110110: color_data = Z;
		19'b0001100110011110111: color_data = Z;
		19'b0001100110011111000: color_data = Z;
		19'b0001100110011111001: color_data = Z;
		19'b0001100110011111010: color_data = Z;
		19'b0001100110011111011: color_data = Z;
		19'b0001100110011111100: color_data = Z;
		19'b0001100110011111101: color_data = Z;
		19'b0001100110011111110: color_data = Z;
		19'b0001100110011111111: color_data = Z;
		19'b0001100110100000000: color_data = Z;
		19'b0001100110100000001: color_data = Z;
		19'b0001100110100000010: color_data = Z;
		19'b0001100110100000011: color_data = Z;
		19'b0001100110100000100: color_data = Z;
		19'b0001100110100000101: color_data = Z;
		19'b0001100110100000110: color_data = Z;
		19'b0001100110100000111: color_data = Z;
		19'b0001100110100001000: color_data = Z;
		19'b0001100110100001001: color_data = Z;
		19'b0001100110100001010: color_data = Z;
		19'b0001100110100001011: color_data = Z;
		19'b0001100110100001100: color_data = Z;
		19'b0001100110100001101: color_data = Z;
		19'b0001100110100001110: color_data = Z;
		19'b0001100110100001111: color_data = Z;
		19'b0001100110100010000: color_data = Z;
		19'b0001100110100010001: color_data = Z;
		19'b0001100110100010010: color_data = Z;
		19'b0001100110100010011: color_data = Z;
		19'b0001100110100010100: color_data = Z;
		19'b0001100110100010101: color_data = Z;
		19'b0001100110100010110: color_data = Z;
		19'b0001100110100010111: color_data = Z;
		19'b0001100110100011000: color_data = Z;
		19'b0001100110100011001: color_data = Z;
		19'b0001100110100011010: color_data = Z;
		19'b0001100110100011011: color_data = Z;
		19'b0001100110100011100: color_data = Z;
		19'b0001100110100011101: color_data = Z;
		19'b0001100110100011110: color_data = Z;
		19'b0001100110100011111: color_data = Z;
		19'b0001100110100100000: color_data = Z;
		19'b0001100110100100001: color_data = Z;
		19'b0001100110100100010: color_data = Z;
		19'b0001100110100100011: color_data = Z;
		19'b0001100110100100100: color_data = Z;
		19'b0001100110100100101: color_data = Z;
		19'b0001100110100100110: color_data = Z;
		19'b0001100110100100111: color_data = Z;
		19'b0001100110100101000: color_data = Z;
		19'b0001100110100101001: color_data = Z;
		19'b0001100110100101010: color_data = Z;
		19'b0001100110100101011: color_data = Z;
		19'b0001100110100101100: color_data = Z;
		19'b0001100110100101101: color_data = Z;
		19'b0001100110100101110: color_data = Z;
		19'b0001100110100101111: color_data = Z;
		19'b0001100110100110000: color_data = Z;
		19'b0001100110100110001: color_data = Z;
		19'b0001100110100110010: color_data = Z;
		19'b0001100110100110011: color_data = Z;
		19'b0001100110100110100: color_data = Z;
		19'b0001100110100110101: color_data = Z;
		19'b0001100110100110110: color_data = Z;
		19'b0001100110100110111: color_data = Z;
		19'b0001100110100111000: color_data = Z;
		19'b0001100110100111001: color_data = Z;
		19'b0001100110100111010: color_data = Z;
		19'b0001100110100111011: color_data = Z;
		19'b0001100110100111100: color_data = Z;
		19'b0001100110100111101: color_data = Z;
		19'b0001100110100111110: color_data = Z;
		19'b0001100110100111111: color_data = Z;
		19'b0001100110101000000: color_data = Z;
		19'b0001100110101000001: color_data = Z;
		19'b0001100110101000010: color_data = Z;
		19'b0001100110101000011: color_data = Z;
		19'b0001100110101000100: color_data = Z;
		19'b0001100110101000101: color_data = Z;
		19'b0001100110101000110: color_data = Z;
		19'b0001100110101000111: color_data = Z;
		19'b0001100110101001000: color_data = Z;
		19'b0001100110101001001: color_data = Z;
		19'b0001100110101001010: color_data = Z;
		19'b0001100110101001011: color_data = Z;
		19'b0001100110101001100: color_data = Z;
		19'b0001100110101001101: color_data = Z;
		19'b0001100110101001110: color_data = Z;
		19'b0001100110101001111: color_data = Z;
		19'b0001100110101010000: color_data = Z;
		19'b0001100110101010001: color_data = Z;
		19'b0001100110101010010: color_data = Z;
		19'b0001100110101010011: color_data = Z;
		19'b0001100110101010100: color_data = Z;
		19'b0001100110101010101: color_data = Z;
		19'b0001100110101010110: color_data = Z;
		19'b0001100110101010111: color_data = Z;
		19'b0001100110101011000: color_data = Z;
		19'b0001100110101011001: color_data = Z;
		19'b0001100110101011010: color_data = Z;
		19'b0001100110101011011: color_data = Z;
		19'b0001100110101011100: color_data = Z;
		19'b0001100110101011101: color_data = Z;
		19'b0001100110101011110: color_data = Z;
		19'b0001100110101011111: color_data = Z;
		19'b0001100110101100000: color_data = Z;
		19'b0001100110101100001: color_data = Z;
		19'b0001100110101100010: color_data = Z;
		19'b0001100110101100011: color_data = Z;
		19'b0001100110101100100: color_data = Z;
		19'b0001100110101100101: color_data = Z;
		19'b0001100110101100110: color_data = Z;
		19'b0001100110101100111: color_data = Z;
		19'b0001100110101101000: color_data = Z;
		19'b0001100110101101001: color_data = Z;
		19'b0001100110101101010: color_data = Z;
		19'b0001100110101101011: color_data = Z;
		19'b0001100110101101100: color_data = Z;
		19'b0001100110101101101: color_data = Z;
		19'b0001100110101101110: color_data = Z;
		19'b0001100110101101111: color_data = Z;
		19'b0001100110101110000: color_data = Z;
		19'b0001100110101110001: color_data = Z;
		19'b0001100110101110010: color_data = Z;
		19'b0001100110101110011: color_data = Z;
		19'b0001100110101110100: color_data = Z;
		19'b0001100110101110101: color_data = Z;
		19'b0001100110101110110: color_data = Z;
		19'b0001100110101110111: color_data = Z;
		19'b0001100110101111000: color_data = Z;
		19'b0001100110101111001: color_data = Z;
		19'b0001100110101111010: color_data = Z;
		19'b0001100110101111011: color_data = Z;
		19'b0001100110101111100: color_data = Z;
		19'b0001100110101111101: color_data = Z;
		19'b0001100110101111110: color_data = Z;
		19'b0001100110101111111: color_data = Z;
		19'b0001100110110000000: color_data = Z;
		19'b0001100110110000001: color_data = Z;
		19'b0001100110110000010: color_data = Z;
		19'b0001100110110000011: color_data = Z;
		19'b0001100110110000100: color_data = Z;
		19'b0001100110110000101: color_data = Z;
		19'b0001100110110000110: color_data = Z;
		19'b0001100110110000111: color_data = Z;
		19'b0001100110110001000: color_data = Z;
		19'b0001100110110001001: color_data = Z;
		19'b0001100110110001010: color_data = Z;
		19'b0001100110110001011: color_data = Z;
		19'b0001100110110001100: color_data = Z;
		19'b0001100110110001101: color_data = Z;
		19'b0001100110110001110: color_data = Z;
		19'b0001100110110001111: color_data = Z;
		19'b0001100110110010000: color_data = Z;
		19'b0001100110110010001: color_data = Z;
		19'b0001100110110010010: color_data = Z;
		19'b0001100110110010011: color_data = Z;
		19'b0001100110110010100: color_data = Z;
		19'b0001100110110010101: color_data = Z;
		19'b0001100110110010110: color_data = Z;
		19'b0001100110110010111: color_data = Z;
		19'b0001100110110011000: color_data = Z;
		19'b0001100110110011001: color_data = Z;
		19'b0001100110110011010: color_data = Z;
		19'b0001100110110011011: color_data = Z;
		19'b0001100110110011100: color_data = Z;
		19'b0001100110110011101: color_data = Z;
		19'b0001100110110011110: color_data = Z;
		19'b0001100110110100011: color_data = Z;
		19'b0001100110110100100: color_data = Z;
		19'b0001100110110100101: color_data = Z;
		19'b0001100110110100110: color_data = Z;
		19'b0001100110110100111: color_data = Z;
		19'b0001100110110101000: color_data = Z;
		19'b0001100110110101111: color_data = Z;
		19'b0001100110110110000: color_data = Z;
		19'b0001100110110110001: color_data = Z;
		19'b0001100110110110010: color_data = Z;
		19'b0001100110110110011: color_data = Z;
		19'b0001100110110110100: color_data = Z;
		19'b0001101000011011011: color_data = Z;
		19'b0001101000011011100: color_data = Z;
		19'b0001101000011011101: color_data = Z;
		19'b0001101000011011110: color_data = Z;
		19'b0001101000011011111: color_data = Z;
		19'b0001101000011100000: color_data = Z;
		19'b0001101000011100001: color_data = Z;
		19'b0001101000011100010: color_data = Z;
		19'b0001101000011100011: color_data = Z;
		19'b0001101000011100100: color_data = Z;
		19'b0001101000011100101: color_data = Z;
		19'b0001101000011100110: color_data = Z;
		19'b0001101000011100111: color_data = Z;
		19'b0001101000011101000: color_data = Z;
		19'b0001101000011101001: color_data = Z;
		19'b0001101000011101010: color_data = Z;
		19'b0001101000011101011: color_data = Z;
		19'b0001101000011101100: color_data = Z;
		19'b0001101000011101101: color_data = Z;
		19'b0001101000011101110: color_data = Z;
		19'b0001101000011101111: color_data = Z;
		19'b0001101000011110000: color_data = Z;
		19'b0001101000011110001: color_data = Z;
		19'b0001101000011110010: color_data = Z;
		19'b0001101000011110011: color_data = Z;
		19'b0001101000011110100: color_data = Z;
		19'b0001101000011110101: color_data = Z;
		19'b0001101000011110110: color_data = Z;
		19'b0001101000011110111: color_data = Z;
		19'b0001101000011111000: color_data = Z;
		19'b0001101000011111001: color_data = Z;
		19'b0001101000011111010: color_data = Z;
		19'b0001101000011111011: color_data = Z;
		19'b0001101000011111100: color_data = Z;
		19'b0001101000011111101: color_data = Z;
		19'b0001101000011111110: color_data = Z;
		19'b0001101000011111111: color_data = Z;
		19'b0001101000100000000: color_data = Z;
		19'b0001101000100000001: color_data = Z;
		19'b0001101000100000010: color_data = Z;
		19'b0001101000100000011: color_data = Z;
		19'b0001101000100000100: color_data = Z;
		19'b0001101000100000101: color_data = Z;
		19'b0001101000100000110: color_data = Z;
		19'b0001101000100000111: color_data = Z;
		19'b0001101000100001000: color_data = Z;
		19'b0001101000100001001: color_data = Z;
		19'b0001101000100001010: color_data = Z;
		19'b0001101000100001011: color_data = Z;
		19'b0001101000100001100: color_data = Z;
		19'b0001101000100001101: color_data = Z;
		19'b0001101000100001110: color_data = Z;
		19'b0001101000100001111: color_data = Z;
		19'b0001101000100010000: color_data = Z;
		19'b0001101000100010001: color_data = Z;
		19'b0001101000100010010: color_data = Z;
		19'b0001101000100010011: color_data = Z;
		19'b0001101000100010100: color_data = Z;
		19'b0001101000100010101: color_data = Z;
		19'b0001101000100010110: color_data = Z;
		19'b0001101000100010111: color_data = Z;
		19'b0001101000100011000: color_data = Z;
		19'b0001101000100011001: color_data = Z;
		19'b0001101000100011010: color_data = Z;
		19'b0001101000100011011: color_data = Z;
		19'b0001101000100011100: color_data = Z;
		19'b0001101000100011101: color_data = Z;
		19'b0001101000100011110: color_data = Z;
		19'b0001101000100011111: color_data = Z;
		19'b0001101000100100000: color_data = Z;
		19'b0001101000100100001: color_data = Z;
		19'b0001101000100100010: color_data = Z;
		19'b0001101000100100011: color_data = Z;
		19'b0001101000100100100: color_data = Z;
		19'b0001101000100100101: color_data = Z;
		19'b0001101000100100110: color_data = Z;
		19'b0001101000100100111: color_data = Z;
		19'b0001101000100101000: color_data = Z;
		19'b0001101000100101001: color_data = Z;
		19'b0001101000100101010: color_data = Z;
		19'b0001101000100101011: color_data = Z;
		19'b0001101000100101100: color_data = Z;
		19'b0001101000100101101: color_data = Z;
		19'b0001101000100101110: color_data = Z;
		19'b0001101000100101111: color_data = Z;
		19'b0001101000100110000: color_data = Z;
		19'b0001101000100110001: color_data = Z;
		19'b0001101000100110010: color_data = Z;
		19'b0001101000100110011: color_data = Z;
		19'b0001101000100110100: color_data = Z;
		19'b0001101000100110101: color_data = Z;
		19'b0001101000100110110: color_data = Z;
		19'b0001101000100110111: color_data = Z;
		19'b0001101000100111000: color_data = Z;
		19'b0001101000100111001: color_data = Z;
		19'b0001101000100111010: color_data = Z;
		19'b0001101000100111011: color_data = Z;
		19'b0001101000100111100: color_data = Z;
		19'b0001101000100111101: color_data = Z;
		19'b0001101000100111110: color_data = Z;
		19'b0001101000100111111: color_data = Z;
		19'b0001101000101000000: color_data = Z;
		19'b0001101000101000001: color_data = Z;
		19'b0001101000101000010: color_data = Z;
		19'b0001101000101000011: color_data = Z;
		19'b0001101000101000100: color_data = Z;
		19'b0001101000101000101: color_data = Z;
		19'b0001101000101000110: color_data = Z;
		19'b0001101000101000111: color_data = Z;
		19'b0001101000101001000: color_data = Z;
		19'b0001101000101001001: color_data = Z;
		19'b0001101000101001010: color_data = Z;
		19'b0001101000101001011: color_data = Z;
		19'b0001101000101001100: color_data = Z;
		19'b0001101000101001101: color_data = Z;
		19'b0001101000101001110: color_data = Z;
		19'b0001101000101001111: color_data = Z;
		19'b0001101000101010000: color_data = Z;
		19'b0001101000101010001: color_data = Z;
		19'b0001101000101010010: color_data = Z;
		19'b0001101000101010011: color_data = Z;
		19'b0001101000101010100: color_data = Z;
		19'b0001101000101010101: color_data = Z;
		19'b0001101000101010110: color_data = Z;
		19'b0001101000101010111: color_data = Z;
		19'b0001101000101011000: color_data = Z;
		19'b0001101000101011001: color_data = Z;
		19'b0001101000101011010: color_data = Z;
		19'b0001101000101011011: color_data = Z;
		19'b0001101000101011100: color_data = Z;
		19'b0001101000101011101: color_data = Z;
		19'b0001101000101011110: color_data = Z;
		19'b0001101000101011111: color_data = Z;
		19'b0001101000101100000: color_data = Z;
		19'b0001101000101100001: color_data = Z;
		19'b0001101000101100010: color_data = Z;
		19'b0001101000101100011: color_data = Z;
		19'b0001101000101100100: color_data = Z;
		19'b0001101000101100101: color_data = Z;
		19'b0001101000101100110: color_data = Z;
		19'b0001101000101100111: color_data = Z;
		19'b0001101000101101000: color_data = Z;
		19'b0001101000101101001: color_data = Z;
		19'b0001101000101101010: color_data = Z;
		19'b0001101000101101011: color_data = Z;
		19'b0001101000101101100: color_data = Z;
		19'b0001101000101101101: color_data = Z;
		19'b0001101000101101110: color_data = Z;
		19'b0001101000101101111: color_data = Z;
		19'b0001101000101110000: color_data = Z;
		19'b0001101000101110001: color_data = Z;
		19'b0001101000101110010: color_data = Z;
		19'b0001101000101110011: color_data = Z;
		19'b0001101000101110100: color_data = Z;
		19'b0001101000101110101: color_data = Z;
		19'b0001101000101110110: color_data = Z;
		19'b0001101000101110111: color_data = Z;
		19'b0001101000101111000: color_data = Z;
		19'b0001101000101111001: color_data = Z;
		19'b0001101000101111010: color_data = Z;
		19'b0001101000101111011: color_data = Z;
		19'b0001101000101111100: color_data = Z;
		19'b0001101000101111101: color_data = Z;
		19'b0001101000101111110: color_data = Z;
		19'b0001101000101111111: color_data = Z;
		19'b0001101000110000000: color_data = Z;
		19'b0001101000110000001: color_data = Z;
		19'b0001101000110000010: color_data = Z;
		19'b0001101000110000011: color_data = Z;
		19'b0001101000110000100: color_data = Z;
		19'b0001101000110000101: color_data = Z;
		19'b0001101000110000110: color_data = Z;
		19'b0001101000110000111: color_data = Z;
		19'b0001101000110001000: color_data = Z;
		19'b0001101000110001001: color_data = Z;
		19'b0001101000110001010: color_data = Z;
		19'b0001101000110001011: color_data = Z;
		19'b0001101000110001100: color_data = Z;
		19'b0001101000110001101: color_data = Z;
		19'b0001101000110001110: color_data = Z;
		19'b0001101000110001111: color_data = Z;
		19'b0001101000110010000: color_data = Z;
		19'b0001101000110010001: color_data = Z;
		19'b0001101000110010010: color_data = Z;
		19'b0001101000110010011: color_data = Z;
		19'b0001101000110010100: color_data = Z;
		19'b0001101000110010101: color_data = Z;
		19'b0001101000110010110: color_data = Z;
		19'b0001101000110010111: color_data = Z;
		19'b0001101000110011000: color_data = Z;
		19'b0001101000110011001: color_data = Z;
		19'b0001101000110011010: color_data = Z;
		19'b0001101000110011011: color_data = Z;
		19'b0001101000110011100: color_data = Z;
		19'b0001101000110011101: color_data = Z;
		19'b0001101000110011110: color_data = Z;
		19'b0001101000110100100: color_data = Z;
		19'b0001101000110100101: color_data = Z;
		19'b0001101000110100110: color_data = Z;
		19'b0001101000110100111: color_data = Z;
		19'b0001101000110101000: color_data = Z;
		19'b0001101000110101001: color_data = Z;
		19'b0001101000110110000: color_data = Z;
		19'b0001101000110110001: color_data = Z;
		19'b0001101000110110010: color_data = Z;
		19'b0001101000110110011: color_data = Z;
		19'b0001101000110110100: color_data = Z;
		19'b0001101000110110101: color_data = Z;
		19'b0001101000110110110: color_data = Z;
		19'b0001101010011011010: color_data = Z;
		19'b0001101010011011011: color_data = Z;
		19'b0001101010011011100: color_data = Z;
		19'b0001101010011011101: color_data = Z;
		19'b0001101010011011110: color_data = Z;
		19'b0001101010011011111: color_data = Z;
		19'b0001101010011100000: color_data = Z;
		19'b0001101010011100001: color_data = Z;
		19'b0001101010011100010: color_data = Z;
		19'b0001101010011100011: color_data = Z;
		19'b0001101010011100100: color_data = Z;
		19'b0001101010011100101: color_data = Z;
		19'b0001101010011100110: color_data = Z;
		19'b0001101010011100111: color_data = Z;
		19'b0001101010011101000: color_data = Z;
		19'b0001101010011101001: color_data = Z;
		19'b0001101010011101010: color_data = Z;
		19'b0001101010011101011: color_data = Z;
		19'b0001101010011101100: color_data = Z;
		19'b0001101010011101101: color_data = Z;
		19'b0001101010011101110: color_data = Z;
		19'b0001101010011101111: color_data = Z;
		19'b0001101010011110000: color_data = Z;
		19'b0001101010011110001: color_data = Z;
		19'b0001101010011110010: color_data = Z;
		19'b0001101010011110011: color_data = Z;
		19'b0001101010011110100: color_data = Z;
		19'b0001101010011110101: color_data = Z;
		19'b0001101010011110110: color_data = Z;
		19'b0001101010011110111: color_data = Z;
		19'b0001101010011111000: color_data = Z;
		19'b0001101010011111001: color_data = Z;
		19'b0001101010011111010: color_data = Z;
		19'b0001101010011111011: color_data = Z;
		19'b0001101010011111100: color_data = Z;
		19'b0001101010011111101: color_data = Z;
		19'b0001101010011111110: color_data = Z;
		19'b0001101010011111111: color_data = Z;
		19'b0001101010100000000: color_data = Z;
		19'b0001101010100000001: color_data = Z;
		19'b0001101010100000010: color_data = Z;
		19'b0001101010100000011: color_data = Z;
		19'b0001101010100000100: color_data = Z;
		19'b0001101010100000101: color_data = Z;
		19'b0001101010100000110: color_data = Z;
		19'b0001101010100000111: color_data = Z;
		19'b0001101010100001000: color_data = Z;
		19'b0001101010100001001: color_data = Z;
		19'b0001101010100001010: color_data = Z;
		19'b0001101010100001011: color_data = Z;
		19'b0001101010100001100: color_data = Z;
		19'b0001101010100001101: color_data = Z;
		19'b0001101010100001110: color_data = Z;
		19'b0001101010100001111: color_data = Z;
		19'b0001101010100010000: color_data = Z;
		19'b0001101010100010001: color_data = Z;
		19'b0001101010100010010: color_data = Z;
		19'b0001101010100010011: color_data = Z;
		19'b0001101010100010100: color_data = Z;
		19'b0001101010100010101: color_data = Z;
		19'b0001101010100010110: color_data = Z;
		19'b0001101010100010111: color_data = Z;
		19'b0001101010100011000: color_data = Z;
		19'b0001101010100011001: color_data = Z;
		19'b0001101010100011010: color_data = Z;
		19'b0001101010100011011: color_data = Z;
		19'b0001101010100011100: color_data = Z;
		19'b0001101010100011101: color_data = Z;
		19'b0001101010100011110: color_data = Z;
		19'b0001101010100011111: color_data = Z;
		19'b0001101010100100000: color_data = Z;
		19'b0001101010100100001: color_data = Z;
		19'b0001101010100100010: color_data = Z;
		19'b0001101010100100011: color_data = Z;
		19'b0001101010100100100: color_data = Z;
		19'b0001101010100100101: color_data = Z;
		19'b0001101010100100110: color_data = Z;
		19'b0001101010100100111: color_data = Z;
		19'b0001101010100101000: color_data = Z;
		19'b0001101010100101001: color_data = Z;
		19'b0001101010100101010: color_data = Z;
		19'b0001101010100101011: color_data = Z;
		19'b0001101010100101100: color_data = Z;
		19'b0001101010100101101: color_data = Z;
		19'b0001101010100101110: color_data = Z;
		19'b0001101010100101111: color_data = Z;
		19'b0001101010100110000: color_data = Z;
		19'b0001101010100110001: color_data = Z;
		19'b0001101010100110010: color_data = Z;
		19'b0001101010100110011: color_data = Z;
		19'b0001101010100110100: color_data = Z;
		19'b0001101010100110101: color_data = Z;
		19'b0001101010100110110: color_data = Z;
		19'b0001101010100110111: color_data = Z;
		19'b0001101010100111000: color_data = Z;
		19'b0001101010100111001: color_data = Z;
		19'b0001101010100111010: color_data = Z;
		19'b0001101010100111011: color_data = Z;
		19'b0001101010100111100: color_data = Z;
		19'b0001101010100111101: color_data = Z;
		19'b0001101010100111110: color_data = Z;
		19'b0001101010100111111: color_data = Z;
		19'b0001101010101000000: color_data = Z;
		19'b0001101010101000001: color_data = Z;
		19'b0001101010101000010: color_data = Z;
		19'b0001101010101000011: color_data = Z;
		19'b0001101010101000100: color_data = Z;
		19'b0001101010101000101: color_data = Z;
		19'b0001101010101000110: color_data = Z;
		19'b0001101010101000111: color_data = Z;
		19'b0001101010101001000: color_data = Z;
		19'b0001101010101001001: color_data = Z;
		19'b0001101010101001010: color_data = Z;
		19'b0001101010101001011: color_data = Z;
		19'b0001101010101001100: color_data = Z;
		19'b0001101010101001101: color_data = Z;
		19'b0001101010101001110: color_data = Z;
		19'b0001101010101001111: color_data = Z;
		19'b0001101010101010000: color_data = Z;
		19'b0001101010101010001: color_data = Z;
		19'b0001101010101010010: color_data = Z;
		19'b0001101010101010011: color_data = Z;
		19'b0001101010101010100: color_data = Z;
		19'b0001101010101010101: color_data = Z;
		19'b0001101010101010110: color_data = Z;
		19'b0001101010101010111: color_data = Z;
		19'b0001101010101011000: color_data = Z;
		19'b0001101010101011001: color_data = Z;
		19'b0001101010101011010: color_data = Z;
		19'b0001101010101011011: color_data = Z;
		19'b0001101010101011100: color_data = Z;
		19'b0001101010101011101: color_data = Z;
		19'b0001101010101011110: color_data = Z;
		19'b0001101010101011111: color_data = Z;
		19'b0001101010101100000: color_data = Z;
		19'b0001101010101100001: color_data = Z;
		19'b0001101010101100010: color_data = Z;
		19'b0001101010101100011: color_data = Z;
		19'b0001101010101100100: color_data = Z;
		19'b0001101010101100101: color_data = Z;
		19'b0001101010101100110: color_data = Z;
		19'b0001101010101100111: color_data = Z;
		19'b0001101010101101000: color_data = Z;
		19'b0001101010101101001: color_data = Z;
		19'b0001101010101101010: color_data = Z;
		19'b0001101010101101011: color_data = Z;
		19'b0001101010101101100: color_data = Z;
		19'b0001101010101101101: color_data = Z;
		19'b0001101010101101110: color_data = Z;
		19'b0001101010101101111: color_data = Z;
		19'b0001101010101110000: color_data = Z;
		19'b0001101010101110001: color_data = Z;
		19'b0001101010101110010: color_data = Z;
		19'b0001101010101110011: color_data = Z;
		19'b0001101010101110100: color_data = Z;
		19'b0001101010101110101: color_data = Z;
		19'b0001101010101110110: color_data = Z;
		19'b0001101010101110111: color_data = Z;
		19'b0001101010101111000: color_data = Z;
		19'b0001101010101111001: color_data = Z;
		19'b0001101010101111010: color_data = Z;
		19'b0001101010101111011: color_data = Z;
		19'b0001101010101111100: color_data = Z;
		19'b0001101010101111101: color_data = Z;
		19'b0001101010101111110: color_data = Z;
		19'b0001101010101111111: color_data = Z;
		19'b0001101010110000000: color_data = Z;
		19'b0001101010110000001: color_data = Z;
		19'b0001101010110000010: color_data = Z;
		19'b0001101010110000011: color_data = Z;
		19'b0001101010110000100: color_data = Z;
		19'b0001101010110000101: color_data = Z;
		19'b0001101010110000110: color_data = Z;
		19'b0001101010110000111: color_data = Z;
		19'b0001101010110001000: color_data = Z;
		19'b0001101010110001001: color_data = Z;
		19'b0001101010110001010: color_data = Z;
		19'b0001101010110001011: color_data = Z;
		19'b0001101010110001100: color_data = Z;
		19'b0001101010110001101: color_data = Z;
		19'b0001101010110001110: color_data = Z;
		19'b0001101010110001111: color_data = Z;
		19'b0001101010110010000: color_data = Z;
		19'b0001101010110010001: color_data = Z;
		19'b0001101010110010010: color_data = Z;
		19'b0001101010110010011: color_data = Z;
		19'b0001101010110010100: color_data = Z;
		19'b0001101010110010101: color_data = Z;
		19'b0001101010110010110: color_data = Z;
		19'b0001101010110010111: color_data = Z;
		19'b0001101010110011000: color_data = Z;
		19'b0001101010110011001: color_data = Z;
		19'b0001101010110011010: color_data = Z;
		19'b0001101010110011011: color_data = Z;
		19'b0001101010110011100: color_data = Z;
		19'b0001101010110011101: color_data = Z;
		19'b0001101010110011110: color_data = Z;
		19'b0001101010110011111: color_data = Z;
		19'b0001101010110100101: color_data = Z;
		19'b0001101010110100110: color_data = Z;
		19'b0001101010110100111: color_data = Z;
		19'b0001101010110101000: color_data = Z;
		19'b0001101010110101001: color_data = Z;
		19'b0001101010110101010: color_data = Z;
		19'b0001101010110110001: color_data = Z;
		19'b0001101010110110010: color_data = Z;
		19'b0001101010110110011: color_data = Z;
		19'b0001101010110110100: color_data = Z;
		19'b0001101010110110101: color_data = Z;
		19'b0001101010110110110: color_data = Z;
		19'b0001101010110110111: color_data = Z;
		19'b0001101100011011001: color_data = Z;
		19'b0001101100011011010: color_data = Z;
		19'b0001101100011011011: color_data = Z;
		19'b0001101100011011100: color_data = Z;
		19'b0001101100011011101: color_data = Z;
		19'b0001101100011011110: color_data = Z;
		19'b0001101100011011111: color_data = Z;
		19'b0001101100011100000: color_data = Z;
		19'b0001101100011100001: color_data = Z;
		19'b0001101100011100010: color_data = Z;
		19'b0001101100011100011: color_data = Z;
		19'b0001101100011100100: color_data = Z;
		19'b0001101100011100101: color_data = Z;
		19'b0001101100011100110: color_data = Z;
		19'b0001101100011100111: color_data = Z;
		19'b0001101100011101000: color_data = Z;
		19'b0001101100011101001: color_data = Z;
		19'b0001101100011101010: color_data = Z;
		19'b0001101100011101011: color_data = Z;
		19'b0001101100011101100: color_data = Z;
		19'b0001101100011101101: color_data = Z;
		19'b0001101100011101110: color_data = Z;
		19'b0001101100011101111: color_data = Z;
		19'b0001101100011110000: color_data = Z;
		19'b0001101100011110001: color_data = Z;
		19'b0001101100011110010: color_data = Z;
		19'b0001101100011110011: color_data = Z;
		19'b0001101100011110100: color_data = Z;
		19'b0001101100011110101: color_data = Z;
		19'b0001101100011110110: color_data = Z;
		19'b0001101100011110111: color_data = Z;
		19'b0001101100011111000: color_data = Z;
		19'b0001101100011111001: color_data = Z;
		19'b0001101100011111010: color_data = Z;
		19'b0001101100011111011: color_data = Z;
		19'b0001101100011111100: color_data = Z;
		19'b0001101100011111101: color_data = Z;
		19'b0001101100011111110: color_data = Z;
		19'b0001101100011111111: color_data = Z;
		19'b0001101100100000000: color_data = Z;
		19'b0001101100100000001: color_data = Z;
		19'b0001101100100000010: color_data = Z;
		19'b0001101100100000011: color_data = Z;
		19'b0001101100100000100: color_data = Z;
		19'b0001101100100000101: color_data = Z;
		19'b0001101100100000110: color_data = Z;
		19'b0001101100100000111: color_data = Z;
		19'b0001101100100001000: color_data = Z;
		19'b0001101100100001001: color_data = Z;
		19'b0001101100100001010: color_data = Z;
		19'b0001101100100001011: color_data = Z;
		19'b0001101100100001100: color_data = Z;
		19'b0001101100100001101: color_data = Z;
		19'b0001101100100001110: color_data = Z;
		19'b0001101100100001111: color_data = Z;
		19'b0001101100100010000: color_data = Z;
		19'b0001101100100010001: color_data = Z;
		19'b0001101100100010010: color_data = Z;
		19'b0001101100100010011: color_data = Z;
		19'b0001101100100010100: color_data = Z;
		19'b0001101100100010101: color_data = Z;
		19'b0001101100100010110: color_data = Z;
		19'b0001101100100010111: color_data = Z;
		19'b0001101100100011000: color_data = Z;
		19'b0001101100100011001: color_data = Z;
		19'b0001101100100011010: color_data = Z;
		19'b0001101100100011011: color_data = Z;
		19'b0001101100100011100: color_data = Z;
		19'b0001101100100011101: color_data = Z;
		19'b0001101100100011110: color_data = Z;
		19'b0001101100100011111: color_data = Z;
		19'b0001101100100100000: color_data = Z;
		19'b0001101100100100001: color_data = Z;
		19'b0001101100100100010: color_data = Z;
		19'b0001101100100100011: color_data = Z;
		19'b0001101100100100100: color_data = Z;
		19'b0001101100100100101: color_data = Z;
		19'b0001101100100100110: color_data = Z;
		19'b0001101100100100111: color_data = Z;
		19'b0001101100100101000: color_data = Z;
		19'b0001101100100101001: color_data = Z;
		19'b0001101100100101010: color_data = Z;
		19'b0001101100100101011: color_data = Z;
		19'b0001101100100101100: color_data = Z;
		19'b0001101100100101101: color_data = Z;
		19'b0001101100100101110: color_data = Z;
		19'b0001101100100101111: color_data = Z;
		19'b0001101100100110000: color_data = Z;
		19'b0001101100100110001: color_data = Z;
		19'b0001101100100110010: color_data = Z;
		19'b0001101100100110011: color_data = Z;
		19'b0001101100100110100: color_data = Z;
		19'b0001101100100110101: color_data = Z;
		19'b0001101100100110110: color_data = Z;
		19'b0001101100100110111: color_data = Z;
		19'b0001101100100111000: color_data = Z;
		19'b0001101100100111001: color_data = Z;
		19'b0001101100100111010: color_data = Z;
		19'b0001101100100111011: color_data = Z;
		19'b0001101100100111100: color_data = Z;
		19'b0001101100100111101: color_data = Z;
		19'b0001101100100111110: color_data = Z;
		19'b0001101100100111111: color_data = Z;
		19'b0001101100101000000: color_data = Z;
		19'b0001101100101000001: color_data = Z;
		19'b0001101100101000010: color_data = Z;
		19'b0001101100101000011: color_data = Z;
		19'b0001101100101000100: color_data = Z;
		19'b0001101100101000101: color_data = Z;
		19'b0001101100101000110: color_data = Z;
		19'b0001101100101000111: color_data = Z;
		19'b0001101100101001000: color_data = Z;
		19'b0001101100101001001: color_data = Z;
		19'b0001101100101001010: color_data = Z;
		19'b0001101100101001011: color_data = Z;
		19'b0001101100101001100: color_data = Z;
		19'b0001101100101001101: color_data = Z;
		19'b0001101100101001110: color_data = Z;
		19'b0001101100101001111: color_data = Z;
		19'b0001101100101010000: color_data = Z;
		19'b0001101100101010001: color_data = Z;
		19'b0001101100101010010: color_data = Z;
		19'b0001101100101010011: color_data = Z;
		19'b0001101100101010100: color_data = Z;
		19'b0001101100101010101: color_data = Z;
		19'b0001101100101010110: color_data = Z;
		19'b0001101100101010111: color_data = Z;
		19'b0001101100101011000: color_data = Z;
		19'b0001101100101011001: color_data = Z;
		19'b0001101100101011010: color_data = Z;
		19'b0001101100101011011: color_data = Z;
		19'b0001101100101011100: color_data = Z;
		19'b0001101100101011101: color_data = Z;
		19'b0001101100101011110: color_data = Z;
		19'b0001101100101011111: color_data = Z;
		19'b0001101100101100000: color_data = Z;
		19'b0001101100101100001: color_data = Z;
		19'b0001101100101100010: color_data = Z;
		19'b0001101100101100011: color_data = Z;
		19'b0001101100101100100: color_data = Z;
		19'b0001101100101100101: color_data = Z;
		19'b0001101100101100110: color_data = Z;
		19'b0001101100101100111: color_data = Z;
		19'b0001101100101101000: color_data = Z;
		19'b0001101100101101001: color_data = Z;
		19'b0001101100101101010: color_data = Z;
		19'b0001101100101101011: color_data = Z;
		19'b0001101100101101100: color_data = Z;
		19'b0001101100101101101: color_data = Z;
		19'b0001101100101101110: color_data = Z;
		19'b0001101100101101111: color_data = Z;
		19'b0001101100101110000: color_data = Z;
		19'b0001101100101110001: color_data = Z;
		19'b0001101100101110010: color_data = Z;
		19'b0001101100101110011: color_data = Z;
		19'b0001101100101110100: color_data = Z;
		19'b0001101100101110101: color_data = Z;
		19'b0001101100101110110: color_data = Z;
		19'b0001101100101110111: color_data = Z;
		19'b0001101100101111000: color_data = Z;
		19'b0001101100101111001: color_data = Z;
		19'b0001101100101111010: color_data = Z;
		19'b0001101100101111011: color_data = Z;
		19'b0001101100101111100: color_data = Z;
		19'b0001101100101111101: color_data = Z;
		19'b0001101100101111110: color_data = Z;
		19'b0001101100101111111: color_data = Z;
		19'b0001101100110000000: color_data = Z;
		19'b0001101100110000001: color_data = Z;
		19'b0001101100110000010: color_data = Z;
		19'b0001101100110000011: color_data = Z;
		19'b0001101100110000100: color_data = Z;
		19'b0001101100110000101: color_data = Z;
		19'b0001101100110000110: color_data = Z;
		19'b0001101100110000111: color_data = Z;
		19'b0001101100110001000: color_data = Z;
		19'b0001101100110001001: color_data = Z;
		19'b0001101100110001010: color_data = Z;
		19'b0001101100110001011: color_data = Z;
		19'b0001101100110001100: color_data = Z;
		19'b0001101100110001101: color_data = Z;
		19'b0001101100110001110: color_data = Z;
		19'b0001101100110001111: color_data = Z;
		19'b0001101100110010000: color_data = Z;
		19'b0001101100110010001: color_data = Z;
		19'b0001101100110010010: color_data = Z;
		19'b0001101100110010011: color_data = Z;
		19'b0001101100110010100: color_data = Z;
		19'b0001101100110010101: color_data = Z;
		19'b0001101100110010110: color_data = Z;
		19'b0001101100110010111: color_data = Z;
		19'b0001101100110011000: color_data = Z;
		19'b0001101100110011001: color_data = Z;
		19'b0001101100110011010: color_data = Z;
		19'b0001101100110011011: color_data = Z;
		19'b0001101100110011100: color_data = Z;
		19'b0001101100110011101: color_data = Z;
		19'b0001101100110011110: color_data = Z;
		19'b0001101100110011111: color_data = Z;
		19'b0001101100110100110: color_data = Z;
		19'b0001101100110100111: color_data = Z;
		19'b0001101100110101000: color_data = Z;
		19'b0001101100110101001: color_data = Z;
		19'b0001101100110101010: color_data = Z;
		19'b0001101100110101011: color_data = Z;
		19'b0001101100110110010: color_data = Z;
		19'b0001101100110110011: color_data = Z;
		19'b0001101100110110100: color_data = Z;
		19'b0001101100110110101: color_data = Z;
		19'b0001101100110110110: color_data = Z;
		19'b0001101100110110111: color_data = Z;
		19'b0001101100110111000: color_data = Z;
		19'b0001101110011011000: color_data = Z;
		19'b0001101110011011001: color_data = Z;
		19'b0001101110011011010: color_data = Z;
		19'b0001101110011011011: color_data = Z;
		19'b0001101110011011100: color_data = Z;
		19'b0001101110011011101: color_data = Z;
		19'b0001101110011011110: color_data = Z;
		19'b0001101110011011111: color_data = Z;
		19'b0001101110011100000: color_data = Z;
		19'b0001101110011100001: color_data = Z;
		19'b0001101110011100010: color_data = Z;
		19'b0001101110011100011: color_data = Z;
		19'b0001101110011100100: color_data = Z;
		19'b0001101110011100101: color_data = Z;
		19'b0001101110011100110: color_data = Z;
		19'b0001101110011100111: color_data = Z;
		19'b0001101110011101000: color_data = Z;
		19'b0001101110011101001: color_data = Z;
		19'b0001101110011101010: color_data = Z;
		19'b0001101110011101011: color_data = Z;
		19'b0001101110011101100: color_data = Z;
		19'b0001101110011101101: color_data = Z;
		19'b0001101110011101110: color_data = Z;
		19'b0001101110011101111: color_data = Z;
		19'b0001101110011110000: color_data = Z;
		19'b0001101110011110001: color_data = Z;
		19'b0001101110011110010: color_data = Z;
		19'b0001101110011110011: color_data = Z;
		19'b0001101110011110100: color_data = Z;
		19'b0001101110011110101: color_data = Z;
		19'b0001101110011110110: color_data = Z;
		19'b0001101110011110111: color_data = Z;
		19'b0001101110011111000: color_data = Z;
		19'b0001101110011111001: color_data = Z;
		19'b0001101110011111010: color_data = Z;
		19'b0001101110011111011: color_data = Z;
		19'b0001101110011111100: color_data = Z;
		19'b0001101110011111101: color_data = Z;
		19'b0001101110011111110: color_data = Z;
		19'b0001101110011111111: color_data = Z;
		19'b0001101110100000000: color_data = Z;
		19'b0001101110100000001: color_data = Z;
		19'b0001101110100000010: color_data = Z;
		19'b0001101110100000011: color_data = Z;
		19'b0001101110100000100: color_data = Z;
		19'b0001101110100000101: color_data = Z;
		19'b0001101110100000110: color_data = Z;
		19'b0001101110100000111: color_data = Z;
		19'b0001101110100001000: color_data = Z;
		19'b0001101110100001001: color_data = Z;
		19'b0001101110100001010: color_data = Z;
		19'b0001101110100001011: color_data = Z;
		19'b0001101110100001100: color_data = Z;
		19'b0001101110100001101: color_data = Z;
		19'b0001101110100001110: color_data = Z;
		19'b0001101110100001111: color_data = Z;
		19'b0001101110100010000: color_data = Z;
		19'b0001101110100010001: color_data = Z;
		19'b0001101110100010010: color_data = Z;
		19'b0001101110100010011: color_data = Z;
		19'b0001101110100010100: color_data = Z;
		19'b0001101110100010101: color_data = Z;
		19'b0001101110100010110: color_data = Z;
		19'b0001101110100010111: color_data = Z;
		19'b0001101110100011000: color_data = Z;
		19'b0001101110100011001: color_data = Z;
		19'b0001101110100011010: color_data = Z;
		19'b0001101110100011011: color_data = Z;
		19'b0001101110100011100: color_data = Z;
		19'b0001101110100011101: color_data = Z;
		19'b0001101110100011110: color_data = Z;
		19'b0001101110100011111: color_data = Z;
		19'b0001101110100100000: color_data = Z;
		19'b0001101110100100001: color_data = Z;
		19'b0001101110100100010: color_data = Z;
		19'b0001101110100100011: color_data = Z;
		19'b0001101110100100100: color_data = Z;
		19'b0001101110100100101: color_data = Z;
		19'b0001101110100100110: color_data = Z;
		19'b0001101110100100111: color_data = Z;
		19'b0001101110100101000: color_data = Z;
		19'b0001101110100101001: color_data = Z;
		19'b0001101110100101010: color_data = Z;
		19'b0001101110100101011: color_data = Z;
		19'b0001101110100101100: color_data = Z;
		19'b0001101110100101101: color_data = Z;
		19'b0001101110100101110: color_data = Z;
		19'b0001101110100101111: color_data = Z;
		19'b0001101110100110000: color_data = Z;
		19'b0001101110100110001: color_data = Z;
		19'b0001101110100110010: color_data = Z;
		19'b0001101110100110011: color_data = Z;
		19'b0001101110100110100: color_data = Z;
		19'b0001101110100110101: color_data = Z;
		19'b0001101110100110110: color_data = Z;
		19'b0001101110100110111: color_data = Z;
		19'b0001101110100111000: color_data = Z;
		19'b0001101110100111001: color_data = Z;
		19'b0001101110100111010: color_data = Z;
		19'b0001101110100111011: color_data = Z;
		19'b0001101110100111100: color_data = Z;
		19'b0001101110100111101: color_data = Z;
		19'b0001101110100111110: color_data = Z;
		19'b0001101110100111111: color_data = Z;
		19'b0001101110101000000: color_data = Z;
		19'b0001101110101000001: color_data = Z;
		19'b0001101110101000010: color_data = Z;
		19'b0001101110101000011: color_data = Z;
		19'b0001101110101000100: color_data = Z;
		19'b0001101110101000101: color_data = Z;
		19'b0001101110101000110: color_data = Z;
		19'b0001101110101000111: color_data = Z;
		19'b0001101110101001000: color_data = Z;
		19'b0001101110101001001: color_data = Z;
		19'b0001101110101001010: color_data = Z;
		19'b0001101110101001011: color_data = Z;
		19'b0001101110101001100: color_data = Z;
		19'b0001101110101001101: color_data = Z;
		19'b0001101110101001110: color_data = Z;
		19'b0001101110101001111: color_data = Z;
		19'b0001101110101010000: color_data = Z;
		19'b0001101110101010001: color_data = Z;
		19'b0001101110101010010: color_data = Z;
		19'b0001101110101010011: color_data = Z;
		19'b0001101110101010100: color_data = Z;
		19'b0001101110101010101: color_data = Z;
		19'b0001101110101010110: color_data = Z;
		19'b0001101110101010111: color_data = Z;
		19'b0001101110101011000: color_data = Z;
		19'b0001101110101011001: color_data = Z;
		19'b0001101110101011010: color_data = Z;
		19'b0001101110101011011: color_data = Z;
		19'b0001101110101011100: color_data = Z;
		19'b0001101110101011101: color_data = Z;
		19'b0001101110101011110: color_data = Z;
		19'b0001101110101011111: color_data = Z;
		19'b0001101110101100000: color_data = Z;
		19'b0001101110101100001: color_data = Z;
		19'b0001101110101100010: color_data = Z;
		19'b0001101110101100011: color_data = Z;
		19'b0001101110101100100: color_data = Z;
		19'b0001101110101100101: color_data = Z;
		19'b0001101110101100110: color_data = Z;
		19'b0001101110101100111: color_data = Z;
		19'b0001101110101101000: color_data = Z;
		19'b0001101110101101001: color_data = Z;
		19'b0001101110101101010: color_data = Z;
		19'b0001101110101101011: color_data = Z;
		19'b0001101110101101100: color_data = Z;
		19'b0001101110101101101: color_data = Z;
		19'b0001101110101101110: color_data = Z;
		19'b0001101110101101111: color_data = Z;
		19'b0001101110101110000: color_data = Z;
		19'b0001101110101110001: color_data = Z;
		19'b0001101110101110010: color_data = Z;
		19'b0001101110101110011: color_data = Z;
		19'b0001101110101110100: color_data = Z;
		19'b0001101110101110101: color_data = Z;
		19'b0001101110101110110: color_data = Z;
		19'b0001101110101110111: color_data = Z;
		19'b0001101110101111000: color_data = Z;
		19'b0001101110101111001: color_data = Z;
		19'b0001101110101111010: color_data = Z;
		19'b0001101110101111011: color_data = Z;
		19'b0001101110101111100: color_data = Z;
		19'b0001101110101111101: color_data = Z;
		19'b0001101110101111110: color_data = Z;
		19'b0001101110101111111: color_data = Z;
		19'b0001101110110000000: color_data = Z;
		19'b0001101110110000001: color_data = Z;
		19'b0001101110110000010: color_data = Z;
		19'b0001101110110000011: color_data = Z;
		19'b0001101110110000100: color_data = Z;
		19'b0001101110110000101: color_data = Z;
		19'b0001101110110000110: color_data = Z;
		19'b0001101110110000111: color_data = Z;
		19'b0001101110110001000: color_data = Z;
		19'b0001101110110001001: color_data = Z;
		19'b0001101110110001010: color_data = Z;
		19'b0001101110110001011: color_data = Z;
		19'b0001101110110001100: color_data = Z;
		19'b0001101110110001101: color_data = Z;
		19'b0001101110110001110: color_data = Z;
		19'b0001101110110001111: color_data = Z;
		19'b0001101110110010000: color_data = Z;
		19'b0001101110110010001: color_data = Z;
		19'b0001101110110010010: color_data = Z;
		19'b0001101110110010011: color_data = Z;
		19'b0001101110110010100: color_data = Z;
		19'b0001101110110010101: color_data = Z;
		19'b0001101110110010110: color_data = Z;
		19'b0001101110110010111: color_data = Z;
		19'b0001101110110011000: color_data = Z;
		19'b0001101110110011001: color_data = Z;
		19'b0001101110110011010: color_data = Z;
		19'b0001101110110011011: color_data = Z;
		19'b0001101110110011100: color_data = Z;
		19'b0001101110110011101: color_data = Z;
		19'b0001101110110011110: color_data = Z;
		19'b0001101110110011111: color_data = Z;
		19'b0001101110110100000: color_data = Z;
		19'b0001101110110100111: color_data = Z;
		19'b0001101110110101000: color_data = Z;
		19'b0001101110110101001: color_data = Z;
		19'b0001101110110101010: color_data = Z;
		19'b0001101110110101011: color_data = Z;
		19'b0001101110110110011: color_data = Z;
		19'b0001101110110110100: color_data = Z;
		19'b0001101110110110101: color_data = Z;
		19'b0001101110110110110: color_data = Z;
		19'b0001101110110110111: color_data = Z;
		19'b0001101110110111000: color_data = Z;
		19'b0001101110110111001: color_data = Z;
		19'b0001110000011010111: color_data = Z;
		19'b0001110000011011000: color_data = Z;
		19'b0001110000011011001: color_data = Z;
		19'b0001110000011011010: color_data = Z;
		19'b0001110000011011011: color_data = Z;
		19'b0001110000011011100: color_data = Z;
		19'b0001110000011011101: color_data = Z;
		19'b0001110000011011110: color_data = Z;
		19'b0001110000011011111: color_data = Z;
		19'b0001110000011100000: color_data = Z;
		19'b0001110000011100001: color_data = Z;
		19'b0001110000011100010: color_data = Z;
		19'b0001110000011100011: color_data = Z;
		19'b0001110000011100100: color_data = Z;
		19'b0001110000011100101: color_data = Z;
		19'b0001110000011100110: color_data = Z;
		19'b0001110000011100111: color_data = Z;
		19'b0001110000011101000: color_data = Z;
		19'b0001110000011101001: color_data = Z;
		19'b0001110000011101010: color_data = Z;
		19'b0001110000011101011: color_data = Z;
		19'b0001110000011101100: color_data = Z;
		19'b0001110000011101101: color_data = Z;
		19'b0001110000011101110: color_data = Z;
		19'b0001110000011101111: color_data = Z;
		19'b0001110000011110000: color_data = Z;
		19'b0001110000011110001: color_data = Z;
		19'b0001110000011110010: color_data = Z;
		19'b0001110000011110011: color_data = Z;
		19'b0001110000011110100: color_data = Z;
		19'b0001110000011110101: color_data = Z;
		19'b0001110000011110110: color_data = Z;
		19'b0001110000011110111: color_data = Z;
		19'b0001110000011111000: color_data = Z;
		19'b0001110000011111001: color_data = Z;
		19'b0001110000011111010: color_data = Z;
		19'b0001110000011111011: color_data = Z;
		19'b0001110000011111100: color_data = Z;
		19'b0001110000011111101: color_data = Z;
		19'b0001110000011111110: color_data = Z;
		19'b0001110000011111111: color_data = Z;
		19'b0001110000100000000: color_data = Z;
		19'b0001110000100000001: color_data = Z;
		19'b0001110000100000010: color_data = Z;
		19'b0001110000100000011: color_data = Z;
		19'b0001110000100000100: color_data = Z;
		19'b0001110000100000101: color_data = Z;
		19'b0001110000100000110: color_data = Z;
		19'b0001110000100000111: color_data = Z;
		19'b0001110000100001000: color_data = Z;
		19'b0001110000100001001: color_data = Z;
		19'b0001110000100001010: color_data = Z;
		19'b0001110000100001011: color_data = Z;
		19'b0001110000100001100: color_data = Z;
		19'b0001110000100001101: color_data = Z;
		19'b0001110000100001110: color_data = Z;
		19'b0001110000100001111: color_data = Z;
		19'b0001110000100010000: color_data = Z;
		19'b0001110000100010001: color_data = Z;
		19'b0001110000100010010: color_data = Z;
		19'b0001110000100010011: color_data = Z;
		19'b0001110000100010100: color_data = Z;
		19'b0001110000100010101: color_data = Z;
		19'b0001110000100010110: color_data = Z;
		19'b0001110000100010111: color_data = Z;
		19'b0001110000100011000: color_data = Z;
		19'b0001110000100011001: color_data = Z;
		19'b0001110000100011010: color_data = Z;
		19'b0001110000100011011: color_data = Z;
		19'b0001110000100011100: color_data = Z;
		19'b0001110000100011101: color_data = Z;
		19'b0001110000100011110: color_data = Z;
		19'b0001110000100011111: color_data = Z;
		19'b0001110000100100000: color_data = Z;
		19'b0001110000100100001: color_data = Z;
		19'b0001110000100100010: color_data = Z;
		19'b0001110000100100011: color_data = Z;
		19'b0001110000100100100: color_data = Z;
		19'b0001110000100100101: color_data = Z;
		19'b0001110000100100110: color_data = Z;
		19'b0001110000100100111: color_data = Z;
		19'b0001110000100101000: color_data = Z;
		19'b0001110000100101001: color_data = Z;
		19'b0001110000100101010: color_data = Z;
		19'b0001110000100101011: color_data = Z;
		19'b0001110000100101100: color_data = Z;
		19'b0001110000100101101: color_data = Z;
		19'b0001110000100101110: color_data = Z;
		19'b0001110000100101111: color_data = Z;
		19'b0001110000100110000: color_data = Z;
		19'b0001110000100110001: color_data = Z;
		19'b0001110000100110010: color_data = Z;
		19'b0001110000100110011: color_data = Z;
		19'b0001110000100110100: color_data = Z;
		19'b0001110000100110101: color_data = Z;
		19'b0001110000100110110: color_data = Z;
		19'b0001110000100110111: color_data = Z;
		19'b0001110000100111000: color_data = Z;
		19'b0001110000100111001: color_data = Z;
		19'b0001110000100111010: color_data = Z;
		19'b0001110000100111011: color_data = Z;
		19'b0001110000100111100: color_data = Z;
		19'b0001110000100111101: color_data = Z;
		19'b0001110000100111110: color_data = Z;
		19'b0001110000100111111: color_data = Z;
		19'b0001110000101000000: color_data = Z;
		19'b0001110000101000001: color_data = Z;
		19'b0001110000101000010: color_data = Z;
		19'b0001110000101000011: color_data = Z;
		19'b0001110000101000100: color_data = Z;
		19'b0001110000101000101: color_data = Z;
		19'b0001110000101000110: color_data = Z;
		19'b0001110000101000111: color_data = Z;
		19'b0001110000101001000: color_data = Z;
		19'b0001110000101001001: color_data = Z;
		19'b0001110000101001010: color_data = Z;
		19'b0001110000101001011: color_data = Z;
		19'b0001110000101001100: color_data = Z;
		19'b0001110000101001101: color_data = Z;
		19'b0001110000101001110: color_data = Z;
		19'b0001110000101001111: color_data = Z;
		19'b0001110000101010000: color_data = Z;
		19'b0001110000101010001: color_data = Z;
		19'b0001110000101010010: color_data = Z;
		19'b0001110000101010011: color_data = Z;
		19'b0001110000101010100: color_data = Z;
		19'b0001110000101010101: color_data = Z;
		19'b0001110000101010110: color_data = Z;
		19'b0001110000101010111: color_data = Z;
		19'b0001110000101011000: color_data = Z;
		19'b0001110000101011001: color_data = Z;
		19'b0001110000101011010: color_data = Z;
		19'b0001110000101011011: color_data = Z;
		19'b0001110000101011100: color_data = Z;
		19'b0001110000101011101: color_data = Z;
		19'b0001110000101011110: color_data = Z;
		19'b0001110000101011111: color_data = Z;
		19'b0001110000101100000: color_data = Z;
		19'b0001110000101100001: color_data = Z;
		19'b0001110000101100010: color_data = Z;
		19'b0001110000101100011: color_data = Z;
		19'b0001110000101100100: color_data = Z;
		19'b0001110000101100101: color_data = Z;
		19'b0001110000101100110: color_data = Z;
		19'b0001110000101100111: color_data = Z;
		19'b0001110000101101000: color_data = Z;
		19'b0001110000101101001: color_data = Z;
		19'b0001110000101101010: color_data = Z;
		19'b0001110000101101011: color_data = Z;
		19'b0001110000101101100: color_data = Z;
		19'b0001110000101101101: color_data = Z;
		19'b0001110000101101110: color_data = Z;
		19'b0001110000101101111: color_data = Z;
		19'b0001110000101110000: color_data = Z;
		19'b0001110000101110001: color_data = Z;
		19'b0001110000101110010: color_data = Z;
		19'b0001110000101110011: color_data = Z;
		19'b0001110000101110100: color_data = Z;
		19'b0001110000101110101: color_data = Z;
		19'b0001110000101110110: color_data = Z;
		19'b0001110000101110111: color_data = Z;
		19'b0001110000101111000: color_data = Z;
		19'b0001110000101111001: color_data = Z;
		19'b0001110000101111010: color_data = Z;
		19'b0001110000101111011: color_data = Z;
		19'b0001110000101111100: color_data = Z;
		19'b0001110000101111101: color_data = Z;
		19'b0001110000101111110: color_data = Z;
		19'b0001110000101111111: color_data = Z;
		19'b0001110000110000000: color_data = Z;
		19'b0001110000110000001: color_data = Z;
		19'b0001110000110000010: color_data = Z;
		19'b0001110000110000011: color_data = Z;
		19'b0001110000110000100: color_data = Z;
		19'b0001110000110000101: color_data = Z;
		19'b0001110000110000110: color_data = Z;
		19'b0001110000110000111: color_data = Z;
		19'b0001110000110001000: color_data = Z;
		19'b0001110000110001001: color_data = Z;
		19'b0001110000110001010: color_data = Z;
		19'b0001110000110001011: color_data = Z;
		19'b0001110000110001100: color_data = Z;
		19'b0001110000110001101: color_data = Z;
		19'b0001110000110001110: color_data = Z;
		19'b0001110000110001111: color_data = Z;
		19'b0001110000110010000: color_data = Z;
		19'b0001110000110010001: color_data = Z;
		19'b0001110000110010010: color_data = Z;
		19'b0001110000110010011: color_data = Z;
		19'b0001110000110010100: color_data = Z;
		19'b0001110000110010101: color_data = Z;
		19'b0001110000110010110: color_data = Z;
		19'b0001110000110010111: color_data = Z;
		19'b0001110000110011000: color_data = Z;
		19'b0001110000110011001: color_data = Z;
		19'b0001110000110011010: color_data = Z;
		19'b0001110000110011011: color_data = Z;
		19'b0001110000110011100: color_data = Z;
		19'b0001110000110011101: color_data = Z;
		19'b0001110000110011110: color_data = Z;
		19'b0001110000110011111: color_data = Z;
		19'b0001110000110100000: color_data = Z;
		19'b0001110000110101000: color_data = Z;
		19'b0001110000110101001: color_data = Z;
		19'b0001110000110101010: color_data = Z;
		19'b0001110000110101011: color_data = Z;
		19'b0001110000110101100: color_data = Z;
		19'b0001110000110110011: color_data = Z;
		19'b0001110000110110100: color_data = Z;
		19'b0001110000110110101: color_data = Z;
		19'b0001110000110110110: color_data = Z;
		19'b0001110000110110111: color_data = Z;
		19'b0001110000110111000: color_data = Z;
		19'b0001110000110111001: color_data = Z;
		19'b0001110000110111010: color_data = Z;
		19'b0001110010011010111: color_data = Z;
		19'b0001110010011011000: color_data = Z;
		19'b0001110010011011001: color_data = Z;
		19'b0001110010011011010: color_data = Z;
		19'b0001110010011011011: color_data = Z;
		19'b0001110010011011100: color_data = Z;
		19'b0001110010011011101: color_data = Z;
		19'b0001110010011011110: color_data = Z;
		19'b0001110010011011111: color_data = Z;
		19'b0001110010011100000: color_data = Z;
		19'b0001110010011100001: color_data = Z;
		19'b0001110010011100010: color_data = Z;
		19'b0001110010011100011: color_data = Z;
		19'b0001110010011100100: color_data = Z;
		19'b0001110010011100101: color_data = Z;
		19'b0001110010011100110: color_data = Z;
		19'b0001110010011100111: color_data = Z;
		19'b0001110010011101000: color_data = Z;
		19'b0001110010011101001: color_data = Z;
		19'b0001110010011101010: color_data = Z;
		19'b0001110010011101011: color_data = Z;
		19'b0001110010011101100: color_data = Z;
		19'b0001110010011101101: color_data = Z;
		19'b0001110010011101110: color_data = Z;
		19'b0001110010011101111: color_data = Z;
		19'b0001110010011110000: color_data = Z;
		19'b0001110010011110001: color_data = Z;
		19'b0001110010011110010: color_data = Z;
		19'b0001110010011110011: color_data = Z;
		19'b0001110010011110100: color_data = Z;
		19'b0001110010011110101: color_data = Z;
		19'b0001110010011110110: color_data = Z;
		19'b0001110010011110111: color_data = Z;
		19'b0001110010011111000: color_data = Z;
		19'b0001110010011111001: color_data = Z;
		19'b0001110010011111010: color_data = Z;
		19'b0001110010011111011: color_data = Z;
		19'b0001110010011111100: color_data = Z;
		19'b0001110010011111101: color_data = Z;
		19'b0001110010011111110: color_data = Z;
		19'b0001110010011111111: color_data = Z;
		19'b0001110010100000000: color_data = Z;
		19'b0001110010100000001: color_data = Z;
		19'b0001110010100000010: color_data = Z;
		19'b0001110010100000011: color_data = Z;
		19'b0001110010100000100: color_data = Z;
		19'b0001110010100000101: color_data = Z;
		19'b0001110010100000110: color_data = Z;
		19'b0001110010100000111: color_data = Z;
		19'b0001110010100001000: color_data = Z;
		19'b0001110010100001001: color_data = Z;
		19'b0001110010100001010: color_data = Z;
		19'b0001110010100001011: color_data = Z;
		19'b0001110010100001100: color_data = Z;
		19'b0001110010100001101: color_data = Z;
		19'b0001110010100001110: color_data = Z;
		19'b0001110010100001111: color_data = Z;
		19'b0001110010100010000: color_data = Z;
		19'b0001110010100010001: color_data = Z;
		19'b0001110010100010010: color_data = Z;
		19'b0001110010100010011: color_data = Z;
		19'b0001110010100010100: color_data = Z;
		19'b0001110010100010101: color_data = Z;
		19'b0001110010100010110: color_data = Z;
		19'b0001110010100010111: color_data = Z;
		19'b0001110010100011000: color_data = Z;
		19'b0001110010100011001: color_data = Z;
		19'b0001110010100011010: color_data = Z;
		19'b0001110010100011011: color_data = Z;
		19'b0001110010100011100: color_data = Z;
		19'b0001110010100011101: color_data = Z;
		19'b0001110010100011110: color_data = Z;
		19'b0001110010100011111: color_data = Z;
		19'b0001110010100100000: color_data = Z;
		19'b0001110010100100001: color_data = Z;
		19'b0001110010100100010: color_data = Z;
		19'b0001110010100100011: color_data = Z;
		19'b0001110010100100100: color_data = Z;
		19'b0001110010100100101: color_data = Z;
		19'b0001110010100100110: color_data = Z;
		19'b0001110010100100111: color_data = Z;
		19'b0001110010100101000: color_data = Z;
		19'b0001110010100101001: color_data = Z;
		19'b0001110010100101010: color_data = Z;
		19'b0001110010100101011: color_data = Z;
		19'b0001110010100101100: color_data = Z;
		19'b0001110010100101101: color_data = Z;
		19'b0001110010100101110: color_data = Z;
		19'b0001110010100101111: color_data = Z;
		19'b0001110010100110000: color_data = Z;
		19'b0001110010100110001: color_data = Z;
		19'b0001110010100110010: color_data = Z;
		19'b0001110010100110011: color_data = Z;
		19'b0001110010100110100: color_data = Z;
		19'b0001110010100110101: color_data = Z;
		19'b0001110010100110110: color_data = Z;
		19'b0001110010100110111: color_data = Z;
		19'b0001110010100111000: color_data = Z;
		19'b0001110010100111001: color_data = Z;
		19'b0001110010100111010: color_data = Z;
		19'b0001110010100111011: color_data = Z;
		19'b0001110010100111100: color_data = Z;
		19'b0001110010100111101: color_data = Z;
		19'b0001110010100111110: color_data = Z;
		19'b0001110010100111111: color_data = Z;
		19'b0001110010101000000: color_data = Z;
		19'b0001110010101000001: color_data = Z;
		19'b0001110010101000010: color_data = Z;
		19'b0001110010101000011: color_data = Z;
		19'b0001110010101000100: color_data = Z;
		19'b0001110010101000101: color_data = Z;
		19'b0001110010101000110: color_data = Z;
		19'b0001110010101000111: color_data = Z;
		19'b0001110010101001000: color_data = Z;
		19'b0001110010101001001: color_data = Z;
		19'b0001110010101001010: color_data = Z;
		19'b0001110010101001011: color_data = Z;
		19'b0001110010101001100: color_data = Z;
		19'b0001110010101001101: color_data = Z;
		19'b0001110010101001110: color_data = Z;
		19'b0001110010101001111: color_data = Z;
		19'b0001110010101010000: color_data = Z;
		19'b0001110010101010001: color_data = Z;
		19'b0001110010101010010: color_data = Z;
		19'b0001110010101010011: color_data = Z;
		19'b0001110010101010100: color_data = Z;
		19'b0001110010101010101: color_data = Z;
		19'b0001110010101010110: color_data = Z;
		19'b0001110010101010111: color_data = Z;
		19'b0001110010101011000: color_data = Z;
		19'b0001110010101011001: color_data = Z;
		19'b0001110010101011010: color_data = Z;
		19'b0001110010101011011: color_data = Z;
		19'b0001110010101011100: color_data = Z;
		19'b0001110010101011101: color_data = Z;
		19'b0001110010101011110: color_data = Z;
		19'b0001110010101011111: color_data = Z;
		19'b0001110010101100000: color_data = Z;
		19'b0001110010101100001: color_data = Z;
		19'b0001110010101100010: color_data = Z;
		19'b0001110010101100011: color_data = Z;
		19'b0001110010101100100: color_data = Z;
		19'b0001110010101100101: color_data = Z;
		19'b0001110010101100110: color_data = Z;
		19'b0001110010101100111: color_data = Z;
		19'b0001110010101101000: color_data = Z;
		19'b0001110010101101001: color_data = Z;
		19'b0001110010101101010: color_data = Z;
		19'b0001110010101101011: color_data = Z;
		19'b0001110010101101100: color_data = Z;
		19'b0001110010101101101: color_data = Z;
		19'b0001110010101101110: color_data = Z;
		19'b0001110010101101111: color_data = Z;
		19'b0001110010101110000: color_data = Z;
		19'b0001110010101110001: color_data = Z;
		19'b0001110010101110010: color_data = Z;
		19'b0001110010101110011: color_data = Z;
		19'b0001110010101110100: color_data = Z;
		19'b0001110010101110101: color_data = Z;
		19'b0001110010101110110: color_data = Z;
		19'b0001110010101110111: color_data = Z;
		19'b0001110010101111000: color_data = Z;
		19'b0001110010101111001: color_data = Z;
		19'b0001110010101111010: color_data = Z;
		19'b0001110010101111011: color_data = Z;
		19'b0001110010101111100: color_data = Z;
		19'b0001110010101111101: color_data = Z;
		19'b0001110010101111110: color_data = Z;
		19'b0001110010101111111: color_data = Z;
		19'b0001110010110000000: color_data = Z;
		19'b0001110010110000001: color_data = Z;
		19'b0001110010110000010: color_data = Z;
		19'b0001110010110000011: color_data = Z;
		19'b0001110010110000100: color_data = Z;
		19'b0001110010110000101: color_data = Z;
		19'b0001110010110000110: color_data = Z;
		19'b0001110010110000111: color_data = Z;
		19'b0001110010110001000: color_data = Z;
		19'b0001110010110001001: color_data = Z;
		19'b0001110010110001010: color_data = Z;
		19'b0001110010110001011: color_data = Z;
		19'b0001110010110001100: color_data = Z;
		19'b0001110010110001101: color_data = Z;
		19'b0001110010110001110: color_data = Z;
		19'b0001110010110001111: color_data = Z;
		19'b0001110010110010000: color_data = Z;
		19'b0001110010110010001: color_data = Z;
		19'b0001110010110010010: color_data = Z;
		19'b0001110010110010011: color_data = Z;
		19'b0001110010110010100: color_data = Z;
		19'b0001110010110010101: color_data = Z;
		19'b0001110010110010110: color_data = Z;
		19'b0001110010110010111: color_data = Z;
		19'b0001110010110011000: color_data = Z;
		19'b0001110010110011001: color_data = Z;
		19'b0001110010110011010: color_data = Z;
		19'b0001110010110011011: color_data = Z;
		19'b0001110010110011100: color_data = Z;
		19'b0001110010110011101: color_data = Z;
		19'b0001110010110011110: color_data = Z;
		19'b0001110010110011111: color_data = Z;
		19'b0001110010110100000: color_data = Z;
		19'b0001110010110100001: color_data = Z;
		19'b0001110010110101001: color_data = Z;
		19'b0001110010110101010: color_data = Z;
		19'b0001110010110101011: color_data = Z;
		19'b0001110010110101100: color_data = Z;
		19'b0001110010110101101: color_data = Z;
		19'b0001110010110110100: color_data = Z;
		19'b0001110010110110101: color_data = Z;
		19'b0001110010110110110: color_data = Z;
		19'b0001110010110110111: color_data = Z;
		19'b0001110010110111000: color_data = Z;
		19'b0001110010110111001: color_data = Z;
		19'b0001110010110111010: color_data = Z;
		19'b0001110010110111011: color_data = Z;
		19'b0001110100011010110: color_data = Z;
		19'b0001110100011010111: color_data = Z;
		19'b0001110100011011000: color_data = Z;
		19'b0001110100011011001: color_data = Z;
		19'b0001110100011011010: color_data = Z;
		19'b0001110100011011011: color_data = Z;
		19'b0001110100011011100: color_data = Z;
		19'b0001110100011011101: color_data = Z;
		19'b0001110100011011110: color_data = Z;
		19'b0001110100011011111: color_data = Z;
		19'b0001110100011100000: color_data = Z;
		19'b0001110100011100001: color_data = Z;
		19'b0001110100011100010: color_data = Z;
		19'b0001110100011100011: color_data = Z;
		19'b0001110100011100100: color_data = Z;
		19'b0001110100011100101: color_data = Z;
		19'b0001110100011100110: color_data = Z;
		19'b0001110100011100111: color_data = Z;
		19'b0001110100011101000: color_data = Z;
		19'b0001110100011101001: color_data = Z;
		19'b0001110100011101010: color_data = Z;
		19'b0001110100011101011: color_data = Z;
		19'b0001110100011101100: color_data = Z;
		19'b0001110100011101101: color_data = Z;
		19'b0001110100011101110: color_data = Z;
		19'b0001110100011101111: color_data = Z;
		19'b0001110100011110000: color_data = Z;
		19'b0001110100011110001: color_data = Z;
		19'b0001110100011110010: color_data = Z;
		19'b0001110100011110011: color_data = Z;
		19'b0001110100011110100: color_data = Z;
		19'b0001110100011110101: color_data = Z;
		19'b0001110100011110110: color_data = Z;
		19'b0001110100011110111: color_data = Z;
		19'b0001110100011111000: color_data = Z;
		19'b0001110100011111001: color_data = Z;
		19'b0001110100011111010: color_data = Z;
		19'b0001110100011111011: color_data = Z;
		19'b0001110100011111100: color_data = Z;
		19'b0001110100011111101: color_data = Z;
		19'b0001110100011111110: color_data = Z;
		19'b0001110100011111111: color_data = Z;
		19'b0001110100100000000: color_data = Z;
		19'b0001110100100000001: color_data = Z;
		19'b0001110100100000010: color_data = Z;
		19'b0001110100100000011: color_data = Z;
		19'b0001110100100000100: color_data = Z;
		19'b0001110100100000101: color_data = Z;
		19'b0001110100100000110: color_data = Z;
		19'b0001110100100000111: color_data = Z;
		19'b0001110100100001000: color_data = Z;
		19'b0001110100100001001: color_data = Z;
		19'b0001110100100001010: color_data = Z;
		19'b0001110100100001011: color_data = Z;
		19'b0001110100100001100: color_data = Z;
		19'b0001110100100001101: color_data = Z;
		19'b0001110100100001110: color_data = Z;
		19'b0001110100100001111: color_data = Z;
		19'b0001110100100010000: color_data = Z;
		19'b0001110100100010001: color_data = Z;
		19'b0001110100100010010: color_data = Z;
		19'b0001110100100010011: color_data = Z;
		19'b0001110100100010100: color_data = Z;
		19'b0001110100100010101: color_data = Z;
		19'b0001110100100010110: color_data = Z;
		19'b0001110100100010111: color_data = Z;
		19'b0001110100100011000: color_data = Z;
		19'b0001110100100011001: color_data = Z;
		19'b0001110100100011010: color_data = Z;
		19'b0001110100100011011: color_data = Z;
		19'b0001110100100011100: color_data = Z;
		19'b0001110100100011101: color_data = Z;
		19'b0001110100100011110: color_data = Z;
		19'b0001110100100011111: color_data = Z;
		19'b0001110100100100000: color_data = Z;
		19'b0001110100100100001: color_data = Z;
		19'b0001110100100100010: color_data = Z;
		19'b0001110100100100011: color_data = Z;
		19'b0001110100100100100: color_data = Z;
		19'b0001110100100100101: color_data = Z;
		19'b0001110100100100110: color_data = Z;
		19'b0001110100100100111: color_data = Z;
		19'b0001110100100101000: color_data = Z;
		19'b0001110100100101001: color_data = Z;
		19'b0001110100100101010: color_data = Z;
		19'b0001110100100101011: color_data = Z;
		19'b0001110100100101100: color_data = Z;
		19'b0001110100100101101: color_data = Z;
		19'b0001110100100101110: color_data = Z;
		19'b0001110100100101111: color_data = Z;
		19'b0001110100100110000: color_data = Z;
		19'b0001110100100110001: color_data = Z;
		19'b0001110100100110010: color_data = Z;
		19'b0001110100100110011: color_data = Z;
		19'b0001110100100110100: color_data = Z;
		19'b0001110100100110101: color_data = Z;
		19'b0001110100100110110: color_data = Z;
		19'b0001110100100110111: color_data = Z;
		19'b0001110100100111000: color_data = Z;
		19'b0001110100100111001: color_data = Z;
		19'b0001110100100111010: color_data = Z;
		19'b0001110100100111011: color_data = Z;
		19'b0001110100100111100: color_data = Z;
		19'b0001110100100111101: color_data = Z;
		19'b0001110100100111110: color_data = Z;
		19'b0001110100100111111: color_data = Z;
		19'b0001110100101000000: color_data = Z;
		19'b0001110100101000001: color_data = Z;
		19'b0001110100101000010: color_data = Z;
		19'b0001110100101000011: color_data = Z;
		19'b0001110100101000100: color_data = Z;
		19'b0001110100101000101: color_data = Z;
		19'b0001110100101000110: color_data = Z;
		19'b0001110100101000111: color_data = Z;
		19'b0001110100101001000: color_data = Z;
		19'b0001110100101001001: color_data = Z;
		19'b0001110100101001010: color_data = Z;
		19'b0001110100101001011: color_data = Z;
		19'b0001110100101001100: color_data = Z;
		19'b0001110100101001101: color_data = Z;
		19'b0001110100101001110: color_data = Z;
		19'b0001110100101001111: color_data = Z;
		19'b0001110100101010000: color_data = Z;
		19'b0001110100101010001: color_data = Z;
		19'b0001110100101010010: color_data = Z;
		19'b0001110100101010011: color_data = Z;
		19'b0001110100101010100: color_data = Z;
		19'b0001110100101010101: color_data = Z;
		19'b0001110100101010110: color_data = Z;
		19'b0001110100101010111: color_data = Z;
		19'b0001110100101011000: color_data = Z;
		19'b0001110100101011001: color_data = Z;
		19'b0001110100101011010: color_data = Z;
		19'b0001110100101011011: color_data = Z;
		19'b0001110100101011100: color_data = Z;
		19'b0001110100101011101: color_data = Z;
		19'b0001110100101011110: color_data = Z;
		19'b0001110100101011111: color_data = Z;
		19'b0001110100101100000: color_data = Z;
		19'b0001110100101100001: color_data = Z;
		19'b0001110100101100010: color_data = Z;
		19'b0001110100101100011: color_data = Z;
		19'b0001110100101100100: color_data = Z;
		19'b0001110100101100101: color_data = Z;
		19'b0001110100101100110: color_data = Z;
		19'b0001110100101100111: color_data = Z;
		19'b0001110100101101000: color_data = Z;
		19'b0001110100101101001: color_data = Z;
		19'b0001110100101101010: color_data = Z;
		19'b0001110100101101011: color_data = Z;
		19'b0001110100101101100: color_data = Z;
		19'b0001110100101101101: color_data = Z;
		19'b0001110100101101110: color_data = Z;
		19'b0001110100101101111: color_data = Z;
		19'b0001110100101110000: color_data = Z;
		19'b0001110100101110001: color_data = Z;
		19'b0001110100101110010: color_data = Z;
		19'b0001110100101110011: color_data = Z;
		19'b0001110100101110100: color_data = Z;
		19'b0001110100101110101: color_data = Z;
		19'b0001110100101110110: color_data = Z;
		19'b0001110100101110111: color_data = Z;
		19'b0001110100101111000: color_data = Z;
		19'b0001110100101111001: color_data = Z;
		19'b0001110100101111010: color_data = Z;
		19'b0001110100101111011: color_data = Z;
		19'b0001110100101111100: color_data = Z;
		19'b0001110100101111101: color_data = Z;
		19'b0001110100101111110: color_data = Z;
		19'b0001110100101111111: color_data = Z;
		19'b0001110100110000000: color_data = Z;
		19'b0001110100110000001: color_data = Z;
		19'b0001110100110000010: color_data = Z;
		19'b0001110100110000011: color_data = Z;
		19'b0001110100110000100: color_data = Z;
		19'b0001110100110000101: color_data = Z;
		19'b0001110100110000110: color_data = Z;
		19'b0001110100110000111: color_data = Z;
		19'b0001110100110001000: color_data = Z;
		19'b0001110100110001001: color_data = Z;
		19'b0001110100110001010: color_data = Z;
		19'b0001110100110001011: color_data = Z;
		19'b0001110100110001100: color_data = Z;
		19'b0001110100110001101: color_data = Z;
		19'b0001110100110001110: color_data = Z;
		19'b0001110100110001111: color_data = Z;
		19'b0001110100110010000: color_data = Z;
		19'b0001110100110010001: color_data = Z;
		19'b0001110100110010010: color_data = Z;
		19'b0001110100110010011: color_data = Z;
		19'b0001110100110010100: color_data = Z;
		19'b0001110100110010101: color_data = Z;
		19'b0001110100110010110: color_data = Z;
		19'b0001110100110010111: color_data = Z;
		19'b0001110100110011000: color_data = Z;
		19'b0001110100110011001: color_data = Z;
		19'b0001110100110011010: color_data = Z;
		19'b0001110100110011011: color_data = Z;
		19'b0001110100110011100: color_data = Z;
		19'b0001110100110011101: color_data = Z;
		19'b0001110100110011110: color_data = Z;
		19'b0001110100110011111: color_data = Z;
		19'b0001110100110100000: color_data = Z;
		19'b0001110100110100001: color_data = Z;
		19'b0001110100110100010: color_data = Z;
		19'b0001110100110101001: color_data = Z;
		19'b0001110100110101010: color_data = Z;
		19'b0001110100110101011: color_data = Z;
		19'b0001110100110101100: color_data = Z;
		19'b0001110100110101101: color_data = Z;
		19'b0001110100110110100: color_data = Z;
		19'b0001110100110110101: color_data = Z;
		19'b0001110100110110110: color_data = Z;
		19'b0001110100110110111: color_data = Z;
		19'b0001110100110111000: color_data = Z;
		19'b0001110100110111001: color_data = Z;
		19'b0001110100110111010: color_data = Z;
		19'b0001110100110111011: color_data = Z;
		19'b0001110100110111100: color_data = Z;
		19'b0001110110011010101: color_data = Z;
		19'b0001110110011010110: color_data = Z;
		19'b0001110110011010111: color_data = Z;
		19'b0001110110011011000: color_data = Z;
		19'b0001110110011011001: color_data = Z;
		19'b0001110110011011010: color_data = Z;
		19'b0001110110011011011: color_data = Z;
		19'b0001110110011011100: color_data = Z;
		19'b0001110110011011101: color_data = Z;
		19'b0001110110011011110: color_data = Z;
		19'b0001110110011011111: color_data = Z;
		19'b0001110110011100000: color_data = Z;
		19'b0001110110011100001: color_data = Z;
		19'b0001110110011100010: color_data = Z;
		19'b0001110110011100011: color_data = Z;
		19'b0001110110011100100: color_data = Z;
		19'b0001110110011100101: color_data = Z;
		19'b0001110110011100110: color_data = Z;
		19'b0001110110011100111: color_data = Z;
		19'b0001110110011101000: color_data = Z;
		19'b0001110110011101001: color_data = Z;
		19'b0001110110011101010: color_data = Z;
		19'b0001110110011101011: color_data = Z;
		19'b0001110110011101100: color_data = Z;
		19'b0001110110011101101: color_data = Z;
		19'b0001110110011101110: color_data = Z;
		19'b0001110110011101111: color_data = Z;
		19'b0001110110011110000: color_data = Z;
		19'b0001110110011110001: color_data = Z;
		19'b0001110110011110010: color_data = Z;
		19'b0001110110011110011: color_data = Z;
		19'b0001110110011110100: color_data = Z;
		19'b0001110110011110101: color_data = Z;
		19'b0001110110011110110: color_data = Z;
		19'b0001110110011110111: color_data = Z;
		19'b0001110110011111000: color_data = Z;
		19'b0001110110011111001: color_data = Z;
		19'b0001110110011111010: color_data = Z;
		19'b0001110110011111011: color_data = Z;
		19'b0001110110011111100: color_data = Z;
		19'b0001110110011111101: color_data = Z;
		19'b0001110110011111110: color_data = Z;
		19'b0001110110011111111: color_data = Z;
		19'b0001110110100000000: color_data = Z;
		19'b0001110110100000001: color_data = Z;
		19'b0001110110100000010: color_data = Z;
		19'b0001110110100000011: color_data = Z;
		19'b0001110110100000100: color_data = Z;
		19'b0001110110100000101: color_data = Z;
		19'b0001110110100000110: color_data = Z;
		19'b0001110110100000111: color_data = Z;
		19'b0001110110100001000: color_data = Z;
		19'b0001110110100001001: color_data = Z;
		19'b0001110110100001010: color_data = Z;
		19'b0001110110100001011: color_data = Z;
		19'b0001110110100001100: color_data = Z;
		19'b0001110110100001101: color_data = Z;
		19'b0001110110100001110: color_data = Z;
		19'b0001110110100001111: color_data = Z;
		19'b0001110110100010000: color_data = Z;
		19'b0001110110100010001: color_data = Z;
		19'b0001110110100010010: color_data = Z;
		19'b0001110110100010011: color_data = Z;
		19'b0001110110100010100: color_data = Z;
		19'b0001110110100010101: color_data = Z;
		19'b0001110110100010110: color_data = Z;
		19'b0001110110100010111: color_data = Z;
		19'b0001110110100011000: color_data = Z;
		19'b0001110110100011001: color_data = Z;
		19'b0001110110100011010: color_data = Z;
		19'b0001110110100011011: color_data = Z;
		19'b0001110110100011100: color_data = Z;
		19'b0001110110100011101: color_data = Z;
		19'b0001110110100011110: color_data = Z;
		19'b0001110110100011111: color_data = Z;
		19'b0001110110100100000: color_data = Z;
		19'b0001110110100100001: color_data = Z;
		19'b0001110110100100010: color_data = Z;
		19'b0001110110100100011: color_data = Z;
		19'b0001110110100100100: color_data = Z;
		19'b0001110110100100101: color_data = Z;
		19'b0001110110100100110: color_data = Z;
		19'b0001110110100100111: color_data = Z;
		19'b0001110110100101000: color_data = Z;
		19'b0001110110100101001: color_data = Z;
		19'b0001110110100101010: color_data = Z;
		19'b0001110110100101011: color_data = Z;
		19'b0001110110100101100: color_data = Z;
		19'b0001110110100101101: color_data = Z;
		19'b0001110110100101110: color_data = Z;
		19'b0001110110100101111: color_data = Z;
		19'b0001110110100110000: color_data = Z;
		19'b0001110110100110001: color_data = Z;
		19'b0001110110100110010: color_data = Z;
		19'b0001110110100110011: color_data = Z;
		19'b0001110110100110100: color_data = Z;
		19'b0001110110100110101: color_data = Z;
		19'b0001110110100110110: color_data = Z;
		19'b0001110110100110111: color_data = Z;
		19'b0001110110100111000: color_data = Z;
		19'b0001110110100111001: color_data = Z;
		19'b0001110110100111010: color_data = Z;
		19'b0001110110100111011: color_data = Z;
		19'b0001110110100111100: color_data = Z;
		19'b0001110110100111101: color_data = Z;
		19'b0001110110100111110: color_data = Z;
		19'b0001110110100111111: color_data = Z;
		19'b0001110110101000000: color_data = Z;
		19'b0001110110101000001: color_data = Z;
		19'b0001110110101000010: color_data = Z;
		19'b0001110110101000011: color_data = Z;
		19'b0001110110101000100: color_data = Z;
		19'b0001110110101000101: color_data = Z;
		19'b0001110110101000110: color_data = Z;
		19'b0001110110101000111: color_data = Z;
		19'b0001110110101001000: color_data = Z;
		19'b0001110110101001001: color_data = Z;
		19'b0001110110101001010: color_data = Z;
		19'b0001110110101001011: color_data = Z;
		19'b0001110110101001100: color_data = Z;
		19'b0001110110101001101: color_data = Z;
		19'b0001110110101001110: color_data = Z;
		19'b0001110110101001111: color_data = Z;
		19'b0001110110101010000: color_data = Z;
		19'b0001110110101010001: color_data = Z;
		19'b0001110110101010010: color_data = Z;
		19'b0001110110101010011: color_data = Z;
		19'b0001110110101010100: color_data = Z;
		19'b0001110110101010101: color_data = Z;
		19'b0001110110101010110: color_data = Z;
		19'b0001110110101010111: color_data = Z;
		19'b0001110110101011000: color_data = Z;
		19'b0001110110101011001: color_data = Z;
		19'b0001110110101011010: color_data = Z;
		19'b0001110110101011011: color_data = Z;
		19'b0001110110101011100: color_data = Z;
		19'b0001110110101011101: color_data = Z;
		19'b0001110110101011110: color_data = Z;
		19'b0001110110101011111: color_data = Z;
		19'b0001110110101100000: color_data = Z;
		19'b0001110110101100001: color_data = Z;
		19'b0001110110101100010: color_data = Z;
		19'b0001110110101100011: color_data = Z;
		19'b0001110110101100100: color_data = Z;
		19'b0001110110101100101: color_data = Z;
		19'b0001110110101100110: color_data = Z;
		19'b0001110110101100111: color_data = Z;
		19'b0001110110101101000: color_data = Z;
		19'b0001110110101101001: color_data = Z;
		19'b0001110110101101010: color_data = Z;
		19'b0001110110101101011: color_data = Z;
		19'b0001110110101101100: color_data = Z;
		19'b0001110110101101101: color_data = Z;
		19'b0001110110101101110: color_data = Z;
		19'b0001110110101101111: color_data = Z;
		19'b0001110110101110000: color_data = Z;
		19'b0001110110101110001: color_data = Z;
		19'b0001110110101110010: color_data = Z;
		19'b0001110110101110011: color_data = Z;
		19'b0001110110101110100: color_data = Z;
		19'b0001110110101110101: color_data = Z;
		19'b0001110110101110110: color_data = Z;
		19'b0001110110101110111: color_data = Z;
		19'b0001110110101111000: color_data = Z;
		19'b0001110110101111001: color_data = Z;
		19'b0001110110101111010: color_data = Z;
		19'b0001110110101111011: color_data = Z;
		19'b0001110110101111100: color_data = Z;
		19'b0001110110101111101: color_data = Z;
		19'b0001110110101111110: color_data = Z;
		19'b0001110110101111111: color_data = Z;
		19'b0001110110110000000: color_data = Z;
		19'b0001110110110000001: color_data = Z;
		19'b0001110110110000010: color_data = Z;
		19'b0001110110110000011: color_data = Z;
		19'b0001110110110000100: color_data = Z;
		19'b0001110110110000101: color_data = Z;
		19'b0001110110110000110: color_data = Z;
		19'b0001110110110000111: color_data = Z;
		19'b0001110110110001000: color_data = Z;
		19'b0001110110110001001: color_data = Z;
		19'b0001110110110001010: color_data = Z;
		19'b0001110110110001011: color_data = Z;
		19'b0001110110110001100: color_data = Z;
		19'b0001110110110001101: color_data = Z;
		19'b0001110110110001110: color_data = Z;
		19'b0001110110110001111: color_data = Z;
		19'b0001110110110010000: color_data = Z;
		19'b0001110110110010001: color_data = Z;
		19'b0001110110110010010: color_data = Z;
		19'b0001110110110010011: color_data = Z;
		19'b0001110110110010100: color_data = Z;
		19'b0001110110110010101: color_data = Z;
		19'b0001110110110010110: color_data = Z;
		19'b0001110110110010111: color_data = Z;
		19'b0001110110110011000: color_data = Z;
		19'b0001110110110011001: color_data = Z;
		19'b0001110110110011010: color_data = Z;
		19'b0001110110110011011: color_data = Z;
		19'b0001110110110011100: color_data = Z;
		19'b0001110110110011101: color_data = Z;
		19'b0001110110110011110: color_data = Z;
		19'b0001110110110011111: color_data = Z;
		19'b0001110110110100000: color_data = Z;
		19'b0001110110110100001: color_data = Z;
		19'b0001110110110100010: color_data = Z;
		19'b0001110110110100011: color_data = Z;
		19'b0001110110110101010: color_data = Z;
		19'b0001110110110101011: color_data = Z;
		19'b0001110110110101100: color_data = Z;
		19'b0001110110110101101: color_data = Z;
		19'b0001110110110101110: color_data = Z;
		19'b0001110110110110101: color_data = Z;
		19'b0001110110110110110: color_data = Z;
		19'b0001110110110110111: color_data = Z;
		19'b0001110110110111000: color_data = Z;
		19'b0001110110110111001: color_data = Z;
		19'b0001110110110111010: color_data = Z;
		19'b0001110110110111011: color_data = Z;
		19'b0001110110110111100: color_data = Z;
		19'b0001110110110111101: color_data = Z;
		19'b0001111000011010100: color_data = Z;
		19'b0001111000011010101: color_data = Z;
		19'b0001111000011010110: color_data = Z;
		19'b0001111000011010111: color_data = Z;
		19'b0001111000011011000: color_data = Z;
		19'b0001111000011011001: color_data = Z;
		19'b0001111000011011010: color_data = Z;
		19'b0001111000011011011: color_data = Z;
		19'b0001111000011011100: color_data = Z;
		19'b0001111000011011101: color_data = Z;
		19'b0001111000011011110: color_data = Z;
		19'b0001111000011011111: color_data = Z;
		19'b0001111000011100000: color_data = Z;
		19'b0001111000011100001: color_data = Z;
		19'b0001111000011100010: color_data = Z;
		19'b0001111000011100011: color_data = Z;
		19'b0001111000011100100: color_data = Z;
		19'b0001111000011100101: color_data = Z;
		19'b0001111000011100110: color_data = Z;
		19'b0001111000011100111: color_data = Z;
		19'b0001111000011101000: color_data = Z;
		19'b0001111000011101001: color_data = Z;
		19'b0001111000011101010: color_data = Z;
		19'b0001111000011101011: color_data = Z;
		19'b0001111000011101100: color_data = Z;
		19'b0001111000011101101: color_data = Z;
		19'b0001111000011101110: color_data = Z;
		19'b0001111000011101111: color_data = Z;
		19'b0001111000011110000: color_data = Z;
		19'b0001111000011110001: color_data = Z;
		19'b0001111000011110010: color_data = Z;
		19'b0001111000011110011: color_data = Z;
		19'b0001111000011110100: color_data = Z;
		19'b0001111000011110101: color_data = Z;
		19'b0001111000011110110: color_data = Z;
		19'b0001111000011110111: color_data = Z;
		19'b0001111000011111000: color_data = Z;
		19'b0001111000011111001: color_data = Z;
		19'b0001111000011111010: color_data = Z;
		19'b0001111000011111011: color_data = Z;
		19'b0001111000011111100: color_data = Z;
		19'b0001111000011111101: color_data = Z;
		19'b0001111000011111110: color_data = Z;
		19'b0001111000011111111: color_data = Z;
		19'b0001111000100000000: color_data = Z;
		19'b0001111000100000001: color_data = Z;
		19'b0001111000100000010: color_data = Z;
		19'b0001111000100000011: color_data = Z;
		19'b0001111000100000100: color_data = Z;
		19'b0001111000100000101: color_data = Z;
		19'b0001111000100000110: color_data = Z;
		19'b0001111000100000111: color_data = Z;
		19'b0001111000100001000: color_data = Z;
		19'b0001111000100001001: color_data = Z;
		19'b0001111000100001010: color_data = Z;
		19'b0001111000100001011: color_data = Z;
		19'b0001111000100001100: color_data = Z;
		19'b0001111000100001101: color_data = Z;
		19'b0001111000100001110: color_data = Z;
		19'b0001111000100001111: color_data = Z;
		19'b0001111000100010000: color_data = Z;
		19'b0001111000100010001: color_data = Z;
		19'b0001111000100010010: color_data = Z;
		19'b0001111000100010011: color_data = Z;
		19'b0001111000100010100: color_data = Z;
		19'b0001111000100010101: color_data = Z;
		19'b0001111000100010110: color_data = Z;
		19'b0001111000100010111: color_data = Z;
		19'b0001111000100011000: color_data = Z;
		19'b0001111000100011001: color_data = Z;
		19'b0001111000100011010: color_data = Z;
		19'b0001111000100011011: color_data = Z;
		19'b0001111000100011100: color_data = Z;
		19'b0001111000100011101: color_data = Z;
		19'b0001111000100011110: color_data = Z;
		19'b0001111000100011111: color_data = Z;
		19'b0001111000100100000: color_data = Z;
		19'b0001111000100100001: color_data = Z;
		19'b0001111000100100010: color_data = Z;
		19'b0001111000100100011: color_data = Z;
		19'b0001111000100100100: color_data = Z;
		19'b0001111000100100101: color_data = Z;
		19'b0001111000100100110: color_data = Z;
		19'b0001111000100100111: color_data = Z;
		19'b0001111000100101000: color_data = Z;
		19'b0001111000100101001: color_data = Z;
		19'b0001111000100101010: color_data = Z;
		19'b0001111000100101011: color_data = Z;
		19'b0001111000100101100: color_data = Z;
		19'b0001111000100101101: color_data = Z;
		19'b0001111000100101110: color_data = Z;
		19'b0001111000100101111: color_data = Z;
		19'b0001111000100110000: color_data = Z;
		19'b0001111000100110001: color_data = Z;
		19'b0001111000100110010: color_data = Z;
		19'b0001111000100110011: color_data = Z;
		19'b0001111000100110100: color_data = Z;
		19'b0001111000100110101: color_data = Z;
		19'b0001111000100110110: color_data = Z;
		19'b0001111000100110111: color_data = Z;
		19'b0001111000100111000: color_data = Z;
		19'b0001111000100111001: color_data = Z;
		19'b0001111000100111010: color_data = Z;
		19'b0001111000100111011: color_data = Z;
		19'b0001111000100111100: color_data = Z;
		19'b0001111000100111101: color_data = Z;
		19'b0001111000100111110: color_data = Z;
		19'b0001111000100111111: color_data = Z;
		19'b0001111000101000000: color_data = Z;
		19'b0001111000101000001: color_data = Z;
		19'b0001111000101000010: color_data = Z;
		19'b0001111000101000011: color_data = Z;
		19'b0001111000101000100: color_data = Z;
		19'b0001111000101000101: color_data = Z;
		19'b0001111000101000110: color_data = Z;
		19'b0001111000101000111: color_data = Z;
		19'b0001111000101001000: color_data = Z;
		19'b0001111000101001001: color_data = Z;
		19'b0001111000101001010: color_data = Z;
		19'b0001111000101001011: color_data = Z;
		19'b0001111000101001100: color_data = Z;
		19'b0001111000101001101: color_data = Z;
		19'b0001111000101001110: color_data = Z;
		19'b0001111000101001111: color_data = Z;
		19'b0001111000101010000: color_data = Z;
		19'b0001111000101010001: color_data = Z;
		19'b0001111000101010010: color_data = Z;
		19'b0001111000101010011: color_data = Z;
		19'b0001111000101010100: color_data = Z;
		19'b0001111000101010101: color_data = Z;
		19'b0001111000101010110: color_data = Z;
		19'b0001111000101010111: color_data = Z;
		19'b0001111000101011000: color_data = Z;
		19'b0001111000101011001: color_data = Z;
		19'b0001111000101011010: color_data = Z;
		19'b0001111000101011011: color_data = Z;
		19'b0001111000101011100: color_data = Z;
		19'b0001111000101011101: color_data = Z;
		19'b0001111000101011110: color_data = Z;
		19'b0001111000101011111: color_data = Z;
		19'b0001111000101100000: color_data = Z;
		19'b0001111000101100001: color_data = Z;
		19'b0001111000101100010: color_data = Z;
		19'b0001111000101100011: color_data = Z;
		19'b0001111000101100100: color_data = Z;
		19'b0001111000101100101: color_data = Z;
		19'b0001111000101100110: color_data = Z;
		19'b0001111000101100111: color_data = Z;
		19'b0001111000101101000: color_data = Z;
		19'b0001111000101101001: color_data = Z;
		19'b0001111000101101010: color_data = Z;
		19'b0001111000101101011: color_data = Z;
		19'b0001111000101101100: color_data = Z;
		19'b0001111000101101101: color_data = Z;
		19'b0001111000101101110: color_data = Z;
		19'b0001111000101101111: color_data = Z;
		19'b0001111000101110000: color_data = Z;
		19'b0001111000101110001: color_data = Z;
		19'b0001111000101110010: color_data = Z;
		19'b0001111000101110011: color_data = Z;
		19'b0001111000101110100: color_data = Z;
		19'b0001111000101110101: color_data = Z;
		19'b0001111000101110110: color_data = Z;
		19'b0001111000101110111: color_data = Z;
		19'b0001111000101111000: color_data = Z;
		19'b0001111000101111001: color_data = Z;
		19'b0001111000101111010: color_data = Z;
		19'b0001111000101111011: color_data = Z;
		19'b0001111000101111100: color_data = Z;
		19'b0001111000101111101: color_data = Z;
		19'b0001111000101111110: color_data = Z;
		19'b0001111000101111111: color_data = Z;
		19'b0001111000110000000: color_data = Z;
		19'b0001111000110000001: color_data = Z;
		19'b0001111000110000010: color_data = Z;
		19'b0001111000110000011: color_data = Z;
		19'b0001111000110000100: color_data = Z;
		19'b0001111000110000101: color_data = Z;
		19'b0001111000110000110: color_data = Z;
		19'b0001111000110000111: color_data = Z;
		19'b0001111000110001000: color_data = Z;
		19'b0001111000110001001: color_data = Z;
		19'b0001111000110001010: color_data = Z;
		19'b0001111000110001011: color_data = Z;
		19'b0001111000110001100: color_data = Z;
		19'b0001111000110001101: color_data = Z;
		19'b0001111000110001110: color_data = Z;
		19'b0001111000110001111: color_data = Z;
		19'b0001111000110010000: color_data = Z;
		19'b0001111000110010001: color_data = Z;
		19'b0001111000110010010: color_data = Z;
		19'b0001111000110010011: color_data = Z;
		19'b0001111000110010100: color_data = Z;
		19'b0001111000110010101: color_data = Z;
		19'b0001111000110010110: color_data = Z;
		19'b0001111000110010111: color_data = Z;
		19'b0001111000110011000: color_data = Z;
		19'b0001111000110011001: color_data = Z;
		19'b0001111000110011010: color_data = Z;
		19'b0001111000110011011: color_data = Z;
		19'b0001111000110011100: color_data = Z;
		19'b0001111000110011101: color_data = Z;
		19'b0001111000110011110: color_data = Z;
		19'b0001111000110011111: color_data = Z;
		19'b0001111000110100000: color_data = Z;
		19'b0001111000110100001: color_data = Z;
		19'b0001111000110100010: color_data = Z;
		19'b0001111000110100011: color_data = Z;
		19'b0001111000110100100: color_data = Z;
		19'b0001111000110101010: color_data = Z;
		19'b0001111000110101011: color_data = Z;
		19'b0001111000110101100: color_data = Z;
		19'b0001111000110101101: color_data = Z;
		19'b0001111000110101110: color_data = Z;
		19'b0001111000110101111: color_data = Z;
		19'b0001111000110110101: color_data = Z;
		19'b0001111000110110110: color_data = Z;
		19'b0001111000110110111: color_data = Z;
		19'b0001111000110111000: color_data = Z;
		19'b0001111000110111001: color_data = Z;
		19'b0001111000110111010: color_data = Z;
		19'b0001111000110111011: color_data = Z;
		19'b0001111000110111100: color_data = Z;
		19'b0001111000110111101: color_data = Z;
		19'b0001111000110111110: color_data = Z;
		19'b0001111010011010011: color_data = Z;
		19'b0001111010011010100: color_data = Z;
		19'b0001111010011010101: color_data = Z;
		19'b0001111010011010110: color_data = Z;
		19'b0001111010011010111: color_data = Z;
		19'b0001111010011011000: color_data = Z;
		19'b0001111010011011001: color_data = Z;
		19'b0001111010011011010: color_data = Z;
		19'b0001111010011011011: color_data = Z;
		19'b0001111010011011100: color_data = Z;
		19'b0001111010011011101: color_data = Z;
		19'b0001111010011011110: color_data = Z;
		19'b0001111010011011111: color_data = Z;
		19'b0001111010011100000: color_data = Z;
		19'b0001111010011100001: color_data = Z;
		19'b0001111010011100010: color_data = Z;
		19'b0001111010011100011: color_data = Z;
		19'b0001111010011100100: color_data = Z;
		19'b0001111010011100101: color_data = Z;
		19'b0001111010011100110: color_data = Z;
		19'b0001111010011100111: color_data = Z;
		19'b0001111010011101000: color_data = Z;
		19'b0001111010011101001: color_data = Z;
		19'b0001111010011101010: color_data = Z;
		19'b0001111010011101011: color_data = Z;
		19'b0001111010011101100: color_data = Z;
		19'b0001111010011101101: color_data = Z;
		19'b0001111010011101110: color_data = Z;
		19'b0001111010011101111: color_data = Z;
		19'b0001111010011110000: color_data = Z;
		19'b0001111010011110001: color_data = Z;
		19'b0001111010011110010: color_data = Z;
		19'b0001111010011110011: color_data = Z;
		19'b0001111010011110100: color_data = Z;
		19'b0001111010011110101: color_data = Z;
		19'b0001111010011110110: color_data = Z;
		19'b0001111010011110111: color_data = Z;
		19'b0001111010011111000: color_data = Z;
		19'b0001111010011111001: color_data = Z;
		19'b0001111010011111010: color_data = Z;
		19'b0001111010011111011: color_data = Z;
		19'b0001111010011111100: color_data = Z;
		19'b0001111010011111101: color_data = Z;
		19'b0001111010011111110: color_data = Z;
		19'b0001111010011111111: color_data = Z;
		19'b0001111010100000000: color_data = Z;
		19'b0001111010100000001: color_data = Z;
		19'b0001111010100000010: color_data = Z;
		19'b0001111010100000011: color_data = Z;
		19'b0001111010100000100: color_data = Z;
		19'b0001111010100000101: color_data = Z;
		19'b0001111010100000110: color_data = Z;
		19'b0001111010100000111: color_data = Z;
		19'b0001111010100001000: color_data = Z;
		19'b0001111010100001001: color_data = Z;
		19'b0001111010100001010: color_data = Z;
		19'b0001111010100001011: color_data = Z;
		19'b0001111010100001100: color_data = Z;
		19'b0001111010100001101: color_data = Z;
		19'b0001111010100001110: color_data = Z;
		19'b0001111010100001111: color_data = Z;
		19'b0001111010100010000: color_data = Z;
		19'b0001111010100010001: color_data = Z;
		19'b0001111010100010010: color_data = Z;
		19'b0001111010100010011: color_data = Z;
		19'b0001111010100010100: color_data = Z;
		19'b0001111010100010101: color_data = Z;
		19'b0001111010100010110: color_data = Z;
		19'b0001111010100010111: color_data = Z;
		19'b0001111010100011000: color_data = Z;
		19'b0001111010100011001: color_data = Z;
		19'b0001111010100011010: color_data = Z;
		19'b0001111010100011011: color_data = Z;
		19'b0001111010100011100: color_data = Z;
		19'b0001111010100011101: color_data = Z;
		19'b0001111010100011110: color_data = Z;
		19'b0001111010100011111: color_data = Z;
		19'b0001111010100100000: color_data = Z;
		19'b0001111010100100001: color_data = Z;
		19'b0001111010100100010: color_data = Z;
		19'b0001111010100100011: color_data = Z;
		19'b0001111010100100100: color_data = Z;
		19'b0001111010100100101: color_data = Z;
		19'b0001111010100100110: color_data = Z;
		19'b0001111010100100111: color_data = Z;
		19'b0001111010100101000: color_data = Z;
		19'b0001111010100101001: color_data = Z;
		19'b0001111010100101010: color_data = Z;
		19'b0001111010100101011: color_data = Z;
		19'b0001111010100101100: color_data = Z;
		19'b0001111010100101101: color_data = Z;
		19'b0001111010100101110: color_data = Z;
		19'b0001111010100101111: color_data = Z;
		19'b0001111010100110000: color_data = Z;
		19'b0001111010100110001: color_data = Z;
		19'b0001111010100110010: color_data = Z;
		19'b0001111010100110011: color_data = Z;
		19'b0001111010100110100: color_data = Z;
		19'b0001111010100110101: color_data = Z;
		19'b0001111010100110110: color_data = Z;
		19'b0001111010100110111: color_data = Z;
		19'b0001111010100111000: color_data = Z;
		19'b0001111010100111001: color_data = Z;
		19'b0001111010100111010: color_data = Z;
		19'b0001111010100111011: color_data = Z;
		19'b0001111010100111100: color_data = Z;
		19'b0001111010100111101: color_data = Z;
		19'b0001111010100111110: color_data = Z;
		19'b0001111010100111111: color_data = Z;
		19'b0001111010101000000: color_data = Z;
		19'b0001111010101000001: color_data = Z;
		19'b0001111010101000010: color_data = Z;
		19'b0001111010101000011: color_data = Z;
		19'b0001111010101000100: color_data = Z;
		19'b0001111010101000101: color_data = Z;
		19'b0001111010101000110: color_data = Z;
		19'b0001111010101000111: color_data = Z;
		19'b0001111010101001000: color_data = Z;
		19'b0001111010101001001: color_data = Z;
		19'b0001111010101001010: color_data = Z;
		19'b0001111010101001011: color_data = Z;
		19'b0001111010101001100: color_data = Z;
		19'b0001111010101001101: color_data = Z;
		19'b0001111010101001110: color_data = Z;
		19'b0001111010101001111: color_data = Z;
		19'b0001111010101010000: color_data = Z;
		19'b0001111010101010001: color_data = Z;
		19'b0001111010101010010: color_data = Z;
		19'b0001111010101010011: color_data = Z;
		19'b0001111010101010100: color_data = Z;
		19'b0001111010101010101: color_data = Z;
		19'b0001111010101010110: color_data = Z;
		19'b0001111010101010111: color_data = Z;
		19'b0001111010101011000: color_data = Z;
		19'b0001111010101011001: color_data = Z;
		19'b0001111010101011010: color_data = Z;
		19'b0001111010101011011: color_data = Z;
		19'b0001111010101011100: color_data = Z;
		19'b0001111010101011101: color_data = Z;
		19'b0001111010101011110: color_data = Z;
		19'b0001111010101011111: color_data = Z;
		19'b0001111010101100000: color_data = Z;
		19'b0001111010101100001: color_data = Z;
		19'b0001111010101100010: color_data = Z;
		19'b0001111010101100011: color_data = Z;
		19'b0001111010101100100: color_data = Z;
		19'b0001111010101100101: color_data = Z;
		19'b0001111010101100110: color_data = Z;
		19'b0001111010101100111: color_data = Z;
		19'b0001111010101101000: color_data = Z;
		19'b0001111010101101001: color_data = Z;
		19'b0001111010101101010: color_data = Z;
		19'b0001111010101101011: color_data = Z;
		19'b0001111010101101100: color_data = Z;
		19'b0001111010101101101: color_data = Z;
		19'b0001111010101101110: color_data = Z;
		19'b0001111010101101111: color_data = Z;
		19'b0001111010101110000: color_data = Z;
		19'b0001111010101110001: color_data = Z;
		19'b0001111010101110010: color_data = Z;
		19'b0001111010101110011: color_data = Z;
		19'b0001111010101110100: color_data = Z;
		19'b0001111010101110101: color_data = Z;
		19'b0001111010101110110: color_data = Z;
		19'b0001111010101110111: color_data = Z;
		19'b0001111010101111000: color_data = Z;
		19'b0001111010101111001: color_data = Z;
		19'b0001111010101111010: color_data = Z;
		19'b0001111010101111011: color_data = Z;
		19'b0001111010101111100: color_data = Z;
		19'b0001111010101111101: color_data = Z;
		19'b0001111010101111110: color_data = Z;
		19'b0001111010101111111: color_data = Z;
		19'b0001111010110000000: color_data = Z;
		19'b0001111010110000001: color_data = Z;
		19'b0001111010110000010: color_data = Z;
		19'b0001111010110000011: color_data = Z;
		19'b0001111010110000100: color_data = Z;
		19'b0001111010110000101: color_data = Z;
		19'b0001111010110000110: color_data = Z;
		19'b0001111010110000111: color_data = Z;
		19'b0001111010110001000: color_data = Z;
		19'b0001111010110001001: color_data = Z;
		19'b0001111010110001010: color_data = Z;
		19'b0001111010110001011: color_data = Z;
		19'b0001111010110001100: color_data = Z;
		19'b0001111010110001101: color_data = Z;
		19'b0001111010110001110: color_data = Z;
		19'b0001111010110001111: color_data = Z;
		19'b0001111010110010000: color_data = Z;
		19'b0001111010110010001: color_data = Z;
		19'b0001111010110010010: color_data = Z;
		19'b0001111010110010011: color_data = Z;
		19'b0001111010110010100: color_data = Z;
		19'b0001111010110010101: color_data = Z;
		19'b0001111010110010110: color_data = Z;
		19'b0001111010110010111: color_data = Z;
		19'b0001111010110011000: color_data = Z;
		19'b0001111010110011001: color_data = Z;
		19'b0001111010110011010: color_data = Z;
		19'b0001111010110011011: color_data = Z;
		19'b0001111010110011100: color_data = Z;
		19'b0001111010110011101: color_data = Z;
		19'b0001111010110011110: color_data = Z;
		19'b0001111010110011111: color_data = Z;
		19'b0001111010110100000: color_data = Z;
		19'b0001111010110100001: color_data = Z;
		19'b0001111010110100010: color_data = Z;
		19'b0001111010110100011: color_data = Z;
		19'b0001111010110100100: color_data = Z;
		19'b0001111010110100101: color_data = Z;
		19'b0001111010110101010: color_data = Z;
		19'b0001111010110101011: color_data = Z;
		19'b0001111010110101100: color_data = Z;
		19'b0001111010110101101: color_data = Z;
		19'b0001111010110101110: color_data = Z;
		19'b0001111010110101111: color_data = Z;
		19'b0001111010110110101: color_data = Z;
		19'b0001111010110110110: color_data = Z;
		19'b0001111010110110111: color_data = Z;
		19'b0001111010110111000: color_data = Z;
		19'b0001111010110111001: color_data = Z;
		19'b0001111010110111010: color_data = Z;
		19'b0001111010110111011: color_data = Z;
		19'b0001111010110111100: color_data = Z;
		19'b0001111010110111101: color_data = Z;
		19'b0001111010110111110: color_data = Z;
		19'b0001111010110111111: color_data = Z;
		19'b0001111100011010010: color_data = Z;
		19'b0001111100011010011: color_data = Z;
		19'b0001111100011010100: color_data = Z;
		19'b0001111100011010101: color_data = Z;
		19'b0001111100011010110: color_data = Z;
		19'b0001111100011010111: color_data = Z;
		19'b0001111100011011000: color_data = Z;
		19'b0001111100011011001: color_data = Z;
		19'b0001111100011011010: color_data = Z;
		19'b0001111100011011011: color_data = Z;
		19'b0001111100011011100: color_data = Z;
		19'b0001111100011011101: color_data = Z;
		19'b0001111100011011110: color_data = Z;
		19'b0001111100011011111: color_data = Z;
		19'b0001111100011100000: color_data = Z;
		19'b0001111100011100001: color_data = Z;
		19'b0001111100011100010: color_data = Z;
		19'b0001111100011100011: color_data = Z;
		19'b0001111100011100100: color_data = Z;
		19'b0001111100011100101: color_data = Z;
		19'b0001111100011100110: color_data = Z;
		19'b0001111100011100111: color_data = Z;
		19'b0001111100011101000: color_data = Z;
		19'b0001111100011101001: color_data = Z;
		19'b0001111100011101010: color_data = Z;
		19'b0001111100011101011: color_data = Z;
		19'b0001111100011101100: color_data = Z;
		19'b0001111100011101101: color_data = Z;
		19'b0001111100011101110: color_data = Z;
		19'b0001111100011101111: color_data = Z;
		19'b0001111100011110000: color_data = Z;
		19'b0001111100011110001: color_data = Z;
		19'b0001111100011110010: color_data = Z;
		19'b0001111100011110011: color_data = Z;
		19'b0001111100011110100: color_data = Z;
		19'b0001111100011110101: color_data = Z;
		19'b0001111100011110110: color_data = Z;
		19'b0001111100011110111: color_data = Z;
		19'b0001111100011111000: color_data = Z;
		19'b0001111100011111001: color_data = Z;
		19'b0001111100011111010: color_data = Z;
		19'b0001111100011111011: color_data = Z;
		19'b0001111100011111100: color_data = Z;
		19'b0001111100011111101: color_data = Z;
		19'b0001111100011111110: color_data = Z;
		19'b0001111100011111111: color_data = Z;
		19'b0001111100100000000: color_data = Z;
		19'b0001111100100000001: color_data = Z;
		19'b0001111100100000010: color_data = Z;
		19'b0001111100100000011: color_data = Z;
		19'b0001111100100000100: color_data = Z;
		19'b0001111100100000101: color_data = Z;
		19'b0001111100100000110: color_data = Z;
		19'b0001111100100000111: color_data = Z;
		19'b0001111100100001000: color_data = Z;
		19'b0001111100100001001: color_data = Z;
		19'b0001111100100001010: color_data = Z;
		19'b0001111100100001011: color_data = Z;
		19'b0001111100100001100: color_data = Z;
		19'b0001111100100001101: color_data = Z;
		19'b0001111100100001110: color_data = Z;
		19'b0001111100100001111: color_data = Z;
		19'b0001111100100010000: color_data = Z;
		19'b0001111100100010001: color_data = Z;
		19'b0001111100100010010: color_data = Z;
		19'b0001111100100010011: color_data = Z;
		19'b0001111100100010100: color_data = Z;
		19'b0001111100100010101: color_data = Z;
		19'b0001111100100010110: color_data = Z;
		19'b0001111100100010111: color_data = Z;
		19'b0001111100100011000: color_data = Z;
		19'b0001111100100011001: color_data = Z;
		19'b0001111100100011010: color_data = Z;
		19'b0001111100100011011: color_data = Z;
		19'b0001111100100011100: color_data = Z;
		19'b0001111100100011101: color_data = Z;
		19'b0001111100100011110: color_data = Z;
		19'b0001111100100011111: color_data = Z;
		19'b0001111100100100000: color_data = Z;
		19'b0001111100100100001: color_data = Z;
		19'b0001111100100100010: color_data = Z;
		19'b0001111100100100011: color_data = Z;
		19'b0001111100100100100: color_data = Z;
		19'b0001111100100100101: color_data = Z;
		19'b0001111100100100110: color_data = Z;
		19'b0001111100100100111: color_data = Z;
		19'b0001111100100101000: color_data = Z;
		19'b0001111100100101001: color_data = Z;
		19'b0001111100100101010: color_data = Z;
		19'b0001111100100101011: color_data = Z;
		19'b0001111100100101100: color_data = Z;
		19'b0001111100100101101: color_data = Z;
		19'b0001111100100101110: color_data = Z;
		19'b0001111100100101111: color_data = Z;
		19'b0001111100100110000: color_data = Z;
		19'b0001111100100110001: color_data = Z;
		19'b0001111100100110010: color_data = Z;
		19'b0001111100100110011: color_data = Z;
		19'b0001111100100110100: color_data = Z;
		19'b0001111100100110101: color_data = Z;
		19'b0001111100100110110: color_data = Z;
		19'b0001111100100110111: color_data = Z;
		19'b0001111100100111000: color_data = Z;
		19'b0001111100100111001: color_data = Z;
		19'b0001111100100111010: color_data = Z;
		19'b0001111100100111011: color_data = Z;
		19'b0001111100100111100: color_data = Z;
		19'b0001111100100111101: color_data = Z;
		19'b0001111100100111110: color_data = Z;
		19'b0001111100100111111: color_data = Z;
		19'b0001111100101000000: color_data = Z;
		19'b0001111100101000001: color_data = Z;
		19'b0001111100101000010: color_data = Z;
		19'b0001111100101000011: color_data = Z;
		19'b0001111100101000100: color_data = Z;
		19'b0001111100101000101: color_data = Z;
		19'b0001111100101000110: color_data = Z;
		19'b0001111100101000111: color_data = Z;
		19'b0001111100101001000: color_data = Z;
		19'b0001111100101001001: color_data = Z;
		19'b0001111100101001010: color_data = Z;
		19'b0001111100101001011: color_data = Z;
		19'b0001111100101001100: color_data = Z;
		19'b0001111100101001101: color_data = Z;
		19'b0001111100101001110: color_data = Z;
		19'b0001111100101001111: color_data = Z;
		19'b0001111100101010000: color_data = Z;
		19'b0001111100101010001: color_data = Z;
		19'b0001111100101010010: color_data = Z;
		19'b0001111100101010011: color_data = Z;
		19'b0001111100101010100: color_data = Z;
		19'b0001111100101010101: color_data = Z;
		19'b0001111100101010110: color_data = Z;
		19'b0001111100101010111: color_data = Z;
		19'b0001111100101011000: color_data = Z;
		19'b0001111100101011001: color_data = Z;
		19'b0001111100101011010: color_data = Z;
		19'b0001111100101011011: color_data = Z;
		19'b0001111100101011100: color_data = Z;
		19'b0001111100101011101: color_data = Z;
		19'b0001111100101011110: color_data = Z;
		19'b0001111100101011111: color_data = Z;
		19'b0001111100101100000: color_data = Z;
		19'b0001111100101100001: color_data = Z;
		19'b0001111100101100010: color_data = Z;
		19'b0001111100101100011: color_data = Z;
		19'b0001111100101100100: color_data = Z;
		19'b0001111100101100101: color_data = Z;
		19'b0001111100101100110: color_data = Z;
		19'b0001111100101100111: color_data = Z;
		19'b0001111100101101000: color_data = Z;
		19'b0001111100101101001: color_data = Z;
		19'b0001111100101101010: color_data = Z;
		19'b0001111100101101011: color_data = Z;
		19'b0001111100101101100: color_data = Z;
		19'b0001111100101101101: color_data = Z;
		19'b0001111100101101110: color_data = Z;
		19'b0001111100101101111: color_data = Z;
		19'b0001111100101110000: color_data = Z;
		19'b0001111100101110001: color_data = Z;
		19'b0001111100101110010: color_data = Z;
		19'b0001111100101110011: color_data = Z;
		19'b0001111100101110100: color_data = Z;
		19'b0001111100101110101: color_data = Z;
		19'b0001111100101110110: color_data = Z;
		19'b0001111100101110111: color_data = Z;
		19'b0001111100101111000: color_data = Z;
		19'b0001111100101111001: color_data = Z;
		19'b0001111100101111010: color_data = Z;
		19'b0001111100101111011: color_data = Z;
		19'b0001111100101111100: color_data = Z;
		19'b0001111100101111101: color_data = Z;
		19'b0001111100101111110: color_data = Z;
		19'b0001111100101111111: color_data = Z;
		19'b0001111100110000000: color_data = Z;
		19'b0001111100110000001: color_data = Z;
		19'b0001111100110000010: color_data = Z;
		19'b0001111100110000011: color_data = Z;
		19'b0001111100110000100: color_data = Z;
		19'b0001111100110000101: color_data = Z;
		19'b0001111100110000110: color_data = Z;
		19'b0001111100110000111: color_data = Z;
		19'b0001111100110001000: color_data = Z;
		19'b0001111100110001001: color_data = Z;
		19'b0001111100110001010: color_data = Z;
		19'b0001111100110001011: color_data = Z;
		19'b0001111100110001100: color_data = Z;
		19'b0001111100110001101: color_data = Z;
		19'b0001111100110001110: color_data = Z;
		19'b0001111100110001111: color_data = Z;
		19'b0001111100110010000: color_data = Z;
		19'b0001111100110010001: color_data = Z;
		19'b0001111100110010010: color_data = Z;
		19'b0001111100110010011: color_data = Z;
		19'b0001111100110010100: color_data = Z;
		19'b0001111100110010101: color_data = Z;
		19'b0001111100110010110: color_data = Z;
		19'b0001111100110010111: color_data = Z;
		19'b0001111100110011000: color_data = Z;
		19'b0001111100110011001: color_data = Z;
		19'b0001111100110011010: color_data = Z;
		19'b0001111100110011011: color_data = Z;
		19'b0001111100110011100: color_data = Z;
		19'b0001111100110011101: color_data = Z;
		19'b0001111100110011110: color_data = Z;
		19'b0001111100110011111: color_data = Z;
		19'b0001111100110100000: color_data = Z;
		19'b0001111100110100001: color_data = Z;
		19'b0001111100110100010: color_data = Z;
		19'b0001111100110100011: color_data = Z;
		19'b0001111100110100100: color_data = Z;
		19'b0001111100110100101: color_data = Z;
		19'b0001111100110100110: color_data = Z;
		19'b0001111100110101011: color_data = Z;
		19'b0001111100110101100: color_data = Z;
		19'b0001111100110101101: color_data = Z;
		19'b0001111100110101110: color_data = Z;
		19'b0001111100110101111: color_data = Z;
		19'b0001111100110110110: color_data = Z;
		19'b0001111100110110111: color_data = Z;
		19'b0001111100110111000: color_data = Z;
		19'b0001111100110111001: color_data = Z;
		19'b0001111100110111010: color_data = Z;
		19'b0001111100110111011: color_data = Z;
		19'b0001111100110111100: color_data = Z;
		19'b0001111100110111101: color_data = Z;
		19'b0001111100110111110: color_data = Z;
		19'b0001111100110111111: color_data = Z;
		19'b0001111100111000000: color_data = Z;
		19'b0001111110011010001: color_data = Z;
		19'b0001111110011010010: color_data = Z;
		19'b0001111110011010011: color_data = Z;
		19'b0001111110011010100: color_data = Z;
		19'b0001111110011010101: color_data = Z;
		19'b0001111110011010110: color_data = Z;
		19'b0001111110011010111: color_data = Z;
		19'b0001111110011011000: color_data = Z;
		19'b0001111110011011001: color_data = Z;
		19'b0001111110011011010: color_data = Z;
		19'b0001111110011011011: color_data = Z;
		19'b0001111110011011100: color_data = Z;
		19'b0001111110011011101: color_data = Z;
		19'b0001111110011011110: color_data = Z;
		19'b0001111110011011111: color_data = Z;
		19'b0001111110011100000: color_data = Z;
		19'b0001111110011100001: color_data = Z;
		19'b0001111110011100010: color_data = Z;
		19'b0001111110011100011: color_data = Z;
		19'b0001111110011100100: color_data = Z;
		19'b0001111110011100101: color_data = Z;
		19'b0001111110011100110: color_data = Z;
		19'b0001111110011100111: color_data = Z;
		19'b0001111110011101000: color_data = Z;
		19'b0001111110011101001: color_data = Z;
		19'b0001111110011101010: color_data = Z;
		19'b0001111110011101011: color_data = Z;
		19'b0001111110011101100: color_data = Z;
		19'b0001111110011101101: color_data = Z;
		19'b0001111110011101110: color_data = Z;
		19'b0001111110011101111: color_data = Z;
		19'b0001111110011110000: color_data = Z;
		19'b0001111110011110001: color_data = Z;
		19'b0001111110011110010: color_data = Z;
		19'b0001111110011110011: color_data = Z;
		19'b0001111110011110100: color_data = Z;
		19'b0001111110011110101: color_data = Z;
		19'b0001111110011110110: color_data = Z;
		19'b0001111110011110111: color_data = Z;
		19'b0001111110011111000: color_data = Z;
		19'b0001111110011111001: color_data = Z;
		19'b0001111110011111010: color_data = Z;
		19'b0001111110011111011: color_data = Z;
		19'b0001111110011111100: color_data = Z;
		19'b0001111110011111101: color_data = Z;
		19'b0001111110011111110: color_data = Z;
		19'b0001111110011111111: color_data = Z;
		19'b0001111110100000000: color_data = Z;
		19'b0001111110100000001: color_data = Z;
		19'b0001111110100000010: color_data = Z;
		19'b0001111110100000011: color_data = Z;
		19'b0001111110100000100: color_data = Z;
		19'b0001111110100000101: color_data = Z;
		19'b0001111110100000110: color_data = Z;
		19'b0001111110100000111: color_data = Z;
		19'b0001111110100001000: color_data = Z;
		19'b0001111110100001001: color_data = Z;
		19'b0001111110100001010: color_data = Z;
		19'b0001111110100001011: color_data = Z;
		19'b0001111110100001100: color_data = Z;
		19'b0001111110100001101: color_data = Z;
		19'b0001111110100001110: color_data = Z;
		19'b0001111110100001111: color_data = Z;
		19'b0001111110100010000: color_data = Z;
		19'b0001111110100010001: color_data = Z;
		19'b0001111110100010010: color_data = Z;
		19'b0001111110100010011: color_data = Z;
		19'b0001111110100010100: color_data = Z;
		19'b0001111110100010101: color_data = Z;
		19'b0001111110100010110: color_data = Z;
		19'b0001111110100010111: color_data = Z;
		19'b0001111110100011000: color_data = Z;
		19'b0001111110100011001: color_data = Z;
		19'b0001111110100011010: color_data = Z;
		19'b0001111110100011011: color_data = Z;
		19'b0001111110100011100: color_data = Z;
		19'b0001111110100011101: color_data = Z;
		19'b0001111110100011110: color_data = Z;
		19'b0001111110100011111: color_data = Z;
		19'b0001111110100100000: color_data = Z;
		19'b0001111110100100001: color_data = Z;
		19'b0001111110100100010: color_data = Z;
		19'b0001111110100100011: color_data = Z;
		19'b0001111110100100100: color_data = Z;
		19'b0001111110100100101: color_data = Z;
		19'b0001111110100100110: color_data = Z;
		19'b0001111110100100111: color_data = Z;
		19'b0001111110100101000: color_data = Z;
		19'b0001111110100101001: color_data = Z;
		19'b0001111110100101010: color_data = Z;
		19'b0001111110100101011: color_data = Z;
		19'b0001111110100101100: color_data = Z;
		19'b0001111110100101101: color_data = Z;
		19'b0001111110100101110: color_data = Z;
		19'b0001111110100101111: color_data = Z;
		19'b0001111110100110000: color_data = Z;
		19'b0001111110100110001: color_data = Z;
		19'b0001111110100110010: color_data = Z;
		19'b0001111110100110011: color_data = Z;
		19'b0001111110100110100: color_data = Z;
		19'b0001111110100110101: color_data = Z;
		19'b0001111110100110110: color_data = Z;
		19'b0001111110100110111: color_data = Z;
		19'b0001111110100111000: color_data = Z;
		19'b0001111110100111001: color_data = Z;
		19'b0001111110100111010: color_data = Z;
		19'b0001111110100111011: color_data = Z;
		19'b0001111110100111100: color_data = Z;
		19'b0001111110100111101: color_data = Z;
		19'b0001111110100111110: color_data = Z;
		19'b0001111110100111111: color_data = Z;
		19'b0001111110101000000: color_data = Z;
		19'b0001111110101000001: color_data = Z;
		19'b0001111110101000010: color_data = Z;
		19'b0001111110101000011: color_data = Z;
		19'b0001111110101000100: color_data = Z;
		19'b0001111110101000101: color_data = Z;
		19'b0001111110101000110: color_data = Z;
		19'b0001111110101000111: color_data = Z;
		19'b0001111110101001000: color_data = Z;
		19'b0001111110101001001: color_data = Z;
		19'b0001111110101001010: color_data = Z;
		19'b0001111110101001011: color_data = Z;
		19'b0001111110101001100: color_data = Z;
		19'b0001111110101001101: color_data = Z;
		19'b0001111110101001110: color_data = Z;
		19'b0001111110101001111: color_data = Z;
		19'b0001111110101010000: color_data = Z;
		19'b0001111110101010001: color_data = Z;
		19'b0001111110101010010: color_data = Z;
		19'b0001111110101010011: color_data = Z;
		19'b0001111110101010100: color_data = Z;
		19'b0001111110101010101: color_data = Z;
		19'b0001111110101010110: color_data = Z;
		19'b0001111110101010111: color_data = Z;
		19'b0001111110101011000: color_data = Z;
		19'b0001111110101011001: color_data = Z;
		19'b0001111110101011010: color_data = Z;
		19'b0001111110101011011: color_data = Z;
		19'b0001111110101011100: color_data = Z;
		19'b0001111110101011101: color_data = Z;
		19'b0001111110101011110: color_data = Z;
		19'b0001111110101011111: color_data = Z;
		19'b0001111110101100000: color_data = Z;
		19'b0001111110101100001: color_data = Z;
		19'b0001111110101100010: color_data = Z;
		19'b0001111110101100011: color_data = Z;
		19'b0001111110101100100: color_data = Z;
		19'b0001111110101100101: color_data = Z;
		19'b0001111110101100110: color_data = Z;
		19'b0001111110101100111: color_data = Z;
		19'b0001111110101101000: color_data = Z;
		19'b0001111110101101001: color_data = Z;
		19'b0001111110101101010: color_data = Z;
		19'b0001111110101101011: color_data = Z;
		19'b0001111110101101100: color_data = Z;
		19'b0001111110101101101: color_data = Z;
		19'b0001111110101101110: color_data = Z;
		19'b0001111110101101111: color_data = Z;
		19'b0001111110101110000: color_data = Z;
		19'b0001111110101110001: color_data = Z;
		19'b0001111110101110010: color_data = Z;
		19'b0001111110101110011: color_data = Z;
		19'b0001111110101110100: color_data = Z;
		19'b0001111110101110101: color_data = Z;
		19'b0001111110101110110: color_data = Z;
		19'b0001111110101110111: color_data = Z;
		19'b0001111110101111000: color_data = Z;
		19'b0001111110101111001: color_data = Z;
		19'b0001111110101111010: color_data = Z;
		19'b0001111110101111011: color_data = Z;
		19'b0001111110101111100: color_data = Z;
		19'b0001111110101111101: color_data = Z;
		19'b0001111110101111110: color_data = Z;
		19'b0001111110101111111: color_data = Z;
		19'b0001111110110000000: color_data = Z;
		19'b0001111110110000001: color_data = Z;
		19'b0001111110110000010: color_data = Z;
		19'b0001111110110000011: color_data = Z;
		19'b0001111110110000100: color_data = Z;
		19'b0001111110110000101: color_data = Z;
		19'b0001111110110000110: color_data = Z;
		19'b0001111110110000111: color_data = Z;
		19'b0001111110110001000: color_data = Z;
		19'b0001111110110001001: color_data = Z;
		19'b0001111110110001010: color_data = Z;
		19'b0001111110110001011: color_data = Z;
		19'b0001111110110001100: color_data = Z;
		19'b0001111110110001101: color_data = Z;
		19'b0001111110110001110: color_data = Z;
		19'b0001111110110001111: color_data = Z;
		19'b0001111110110010000: color_data = Z;
		19'b0001111110110010001: color_data = Z;
		19'b0001111110110010010: color_data = Z;
		19'b0001111110110010011: color_data = Z;
		19'b0001111110110010100: color_data = Z;
		19'b0001111110110010101: color_data = Z;
		19'b0001111110110010110: color_data = Z;
		19'b0001111110110010111: color_data = Z;
		19'b0001111110110011000: color_data = Z;
		19'b0001111110110011001: color_data = Z;
		19'b0001111110110011010: color_data = Z;
		19'b0001111110110011011: color_data = Z;
		19'b0001111110110011100: color_data = Z;
		19'b0001111110110011101: color_data = Z;
		19'b0001111110110011110: color_data = Z;
		19'b0001111110110011111: color_data = Z;
		19'b0001111110110100000: color_data = Z;
		19'b0001111110110100001: color_data = Z;
		19'b0001111110110100010: color_data = Z;
		19'b0001111110110100011: color_data = Z;
		19'b0001111110110100100: color_data = Z;
		19'b0001111110110100101: color_data = Z;
		19'b0001111110110100110: color_data = Z;
		19'b0001111110110100111: color_data = Z;
		19'b0001111110110101011: color_data = Z;
		19'b0001111110110101100: color_data = Z;
		19'b0001111110110101101: color_data = Z;
		19'b0001111110110101110: color_data = Z;
		19'b0001111110110101111: color_data = Z;
		19'b0001111110110110000: color_data = Z;
		19'b0001111110110110110: color_data = Z;
		19'b0001111110110110111: color_data = Z;
		19'b0001111110110111000: color_data = Z;
		19'b0001111110110111001: color_data = Z;
		19'b0001111110110111010: color_data = Z;
		19'b0001111110110111011: color_data = Z;
		19'b0001111110110111100: color_data = Z;
		19'b0001111110110111101: color_data = Z;
		19'b0001111110110111110: color_data = Z;
		19'b0001111110110111111: color_data = Z;
		19'b0001111110111000000: color_data = Z;
		19'b0001111110111000001: color_data = Z;
		19'b0010000000011010000: color_data = Z;
		19'b0010000000011010001: color_data = Z;
		19'b0010000000011010010: color_data = Z;
		19'b0010000000011010011: color_data = Z;
		19'b0010000000011010100: color_data = Z;
		19'b0010000000011010101: color_data = Z;
		19'b0010000000011010110: color_data = Z;
		19'b0010000000011010111: color_data = Z;
		19'b0010000000011011000: color_data = Z;
		19'b0010000000011011001: color_data = Z;
		19'b0010000000011011010: color_data = Z;
		19'b0010000000011011011: color_data = Z;
		19'b0010000000011011100: color_data = Z;
		19'b0010000000011011101: color_data = Z;
		19'b0010000000011011110: color_data = Z;
		19'b0010000000011011111: color_data = Z;
		19'b0010000000011100000: color_data = Z;
		19'b0010000000011100001: color_data = Z;
		19'b0010000000011100010: color_data = Z;
		19'b0010000000011100011: color_data = Z;
		19'b0010000000011100100: color_data = Z;
		19'b0010000000011100101: color_data = Z;
		19'b0010000000011100110: color_data = Z;
		19'b0010000000011100111: color_data = Z;
		19'b0010000000011101000: color_data = Z;
		19'b0010000000011101001: color_data = Z;
		19'b0010000000011101010: color_data = Z;
		19'b0010000000011101011: color_data = Z;
		19'b0010000000011101100: color_data = Z;
		19'b0010000000011101101: color_data = Z;
		19'b0010000000011101110: color_data = Z;
		19'b0010000000011101111: color_data = Z;
		19'b0010000000011110000: color_data = Z;
		19'b0010000000011110001: color_data = Z;
		19'b0010000000011110010: color_data = Z;
		19'b0010000000011110011: color_data = Z;
		19'b0010000000011110100: color_data = Z;
		19'b0010000000011110101: color_data = Z;
		19'b0010000000011110110: color_data = Z;
		19'b0010000000011110111: color_data = Z;
		19'b0010000000011111000: color_data = Z;
		19'b0010000000011111001: color_data = Z;
		19'b0010000000011111010: color_data = Z;
		19'b0010000000011111011: color_data = Z;
		19'b0010000000011111100: color_data = Z;
		19'b0010000000011111101: color_data = Z;
		19'b0010000000011111110: color_data = Z;
		19'b0010000000011111111: color_data = Z;
		19'b0010000000100000000: color_data = Z;
		19'b0010000000100000001: color_data = Z;
		19'b0010000000100000010: color_data = Z;
		19'b0010000000100000011: color_data = Z;
		19'b0010000000100000100: color_data = Z;
		19'b0010000000100000101: color_data = Z;
		19'b0010000000100000110: color_data = Z;
		19'b0010000000100000111: color_data = Z;
		19'b0010000000100001000: color_data = Z;
		19'b0010000000100001001: color_data = Z;
		19'b0010000000100001010: color_data = Z;
		19'b0010000000100001011: color_data = Z;
		19'b0010000000100001100: color_data = Z;
		19'b0010000000100001101: color_data = Z;
		19'b0010000000100001110: color_data = Z;
		19'b0010000000100001111: color_data = Z;
		19'b0010000000100010000: color_data = Z;
		19'b0010000000100010001: color_data = Z;
		19'b0010000000100010010: color_data = Z;
		19'b0010000000100010011: color_data = Z;
		19'b0010000000100010100: color_data = Z;
		19'b0010000000100010101: color_data = Z;
		19'b0010000000100010110: color_data = Z;
		19'b0010000000100010111: color_data = Z;
		19'b0010000000100011000: color_data = Z;
		19'b0010000000100011001: color_data = Z;
		19'b0010000000100011010: color_data = Z;
		19'b0010000000100011011: color_data = Z;
		19'b0010000000100011100: color_data = Z;
		19'b0010000000100011101: color_data = Z;
		19'b0010000000100011110: color_data = Z;
		19'b0010000000100011111: color_data = Z;
		19'b0010000000100100000: color_data = Z;
		19'b0010000000100100001: color_data = Z;
		19'b0010000000100100010: color_data = Z;
		19'b0010000000100100011: color_data = Z;
		19'b0010000000100100100: color_data = Z;
		19'b0010000000100100101: color_data = Z;
		19'b0010000000100100110: color_data = Z;
		19'b0010000000100100111: color_data = Z;
		19'b0010000000100101000: color_data = Z;
		19'b0010000000100101001: color_data = Z;
		19'b0010000000100101010: color_data = Z;
		19'b0010000000100101011: color_data = Z;
		19'b0010000000100101100: color_data = Z;
		19'b0010000000100101101: color_data = Z;
		19'b0010000000100101110: color_data = Z;
		19'b0010000000100101111: color_data = Z;
		19'b0010000000100110000: color_data = Z;
		19'b0010000000100110001: color_data = Z;
		19'b0010000000100110010: color_data = Z;
		19'b0010000000100110011: color_data = Z;
		19'b0010000000100110100: color_data = Z;
		19'b0010000000100110101: color_data = Z;
		19'b0010000000100110110: color_data = Z;
		19'b0010000000100110111: color_data = Z;
		19'b0010000000100111000: color_data = Z;
		19'b0010000000100111001: color_data = Z;
		19'b0010000000100111010: color_data = Z;
		19'b0010000000100111011: color_data = Z;
		19'b0010000000100111100: color_data = Z;
		19'b0010000000100111101: color_data = Z;
		19'b0010000000100111110: color_data = Z;
		19'b0010000000100111111: color_data = Z;
		19'b0010000000101000000: color_data = Z;
		19'b0010000000101000001: color_data = Z;
		19'b0010000000101000010: color_data = Z;
		19'b0010000000101000011: color_data = Z;
		19'b0010000000101000100: color_data = Z;
		19'b0010000000101000101: color_data = Z;
		19'b0010000000101000110: color_data = Z;
		19'b0010000000101000111: color_data = Z;
		19'b0010000000101001000: color_data = Z;
		19'b0010000000101001001: color_data = Z;
		19'b0010000000101001010: color_data = Z;
		19'b0010000000101001011: color_data = Z;
		19'b0010000000101001100: color_data = Z;
		19'b0010000000101001101: color_data = Z;
		19'b0010000000101001110: color_data = Z;
		19'b0010000000101001111: color_data = Z;
		19'b0010000000101010000: color_data = Z;
		19'b0010000000101010001: color_data = Z;
		19'b0010000000101010010: color_data = Z;
		19'b0010000000101010011: color_data = Z;
		19'b0010000000101010100: color_data = Z;
		19'b0010000000101010101: color_data = Z;
		19'b0010000000101010110: color_data = Z;
		19'b0010000000101010111: color_data = Z;
		19'b0010000000101011000: color_data = Z;
		19'b0010000000101011001: color_data = Z;
		19'b0010000000101011010: color_data = Z;
		19'b0010000000101011011: color_data = Z;
		19'b0010000000101011100: color_data = Z;
		19'b0010000000101011101: color_data = Z;
		19'b0010000000101011110: color_data = Z;
		19'b0010000000101011111: color_data = Z;
		19'b0010000000101100000: color_data = Z;
		19'b0010000000101100001: color_data = Z;
		19'b0010000000101100010: color_data = Z;
		19'b0010000000101100011: color_data = Z;
		19'b0010000000101100100: color_data = Z;
		19'b0010000000101100101: color_data = Z;
		19'b0010000000101100110: color_data = Z;
		19'b0010000000101100111: color_data = Z;
		19'b0010000000101101000: color_data = Z;
		19'b0010000000101101001: color_data = Z;
		19'b0010000000101101010: color_data = Z;
		19'b0010000000101101011: color_data = Z;
		19'b0010000000101101100: color_data = Z;
		19'b0010000000101101101: color_data = Z;
		19'b0010000000101101110: color_data = Z;
		19'b0010000000101101111: color_data = Z;
		19'b0010000000101110000: color_data = Z;
		19'b0010000000101110001: color_data = Z;
		19'b0010000000101110010: color_data = Z;
		19'b0010000000101110011: color_data = Z;
		19'b0010000000101110100: color_data = Z;
		19'b0010000000101110101: color_data = Z;
		19'b0010000000101110110: color_data = Z;
		19'b0010000000101110111: color_data = Z;
		19'b0010000000101111000: color_data = Z;
		19'b0010000000101111001: color_data = Z;
		19'b0010000000101111010: color_data = Z;
		19'b0010000000101111011: color_data = Z;
		19'b0010000000101111100: color_data = Z;
		19'b0010000000101111101: color_data = Z;
		19'b0010000000101111110: color_data = Z;
		19'b0010000000101111111: color_data = Z;
		19'b0010000000110000000: color_data = Z;
		19'b0010000000110000001: color_data = Z;
		19'b0010000000110000010: color_data = Z;
		19'b0010000000110000011: color_data = Z;
		19'b0010000000110000100: color_data = Z;
		19'b0010000000110000101: color_data = Z;
		19'b0010000000110000110: color_data = Z;
		19'b0010000000110000111: color_data = Z;
		19'b0010000000110001000: color_data = Z;
		19'b0010000000110001001: color_data = Z;
		19'b0010000000110001010: color_data = Z;
		19'b0010000000110001011: color_data = Z;
		19'b0010000000110001100: color_data = Z;
		19'b0010000000110001101: color_data = Z;
		19'b0010000000110001110: color_data = Z;
		19'b0010000000110001111: color_data = Z;
		19'b0010000000110010000: color_data = Z;
		19'b0010000000110010001: color_data = Z;
		19'b0010000000110010010: color_data = Z;
		19'b0010000000110010011: color_data = Z;
		19'b0010000000110010100: color_data = Z;
		19'b0010000000110010101: color_data = Z;
		19'b0010000000110010110: color_data = Z;
		19'b0010000000110010111: color_data = Z;
		19'b0010000000110011000: color_data = Z;
		19'b0010000000110011001: color_data = Z;
		19'b0010000000110011010: color_data = Z;
		19'b0010000000110011011: color_data = Z;
		19'b0010000000110011100: color_data = Z;
		19'b0010000000110011101: color_data = Z;
		19'b0010000000110011110: color_data = Z;
		19'b0010000000110011111: color_data = Z;
		19'b0010000000110100000: color_data = Z;
		19'b0010000000110100001: color_data = Z;
		19'b0010000000110100010: color_data = Z;
		19'b0010000000110100011: color_data = Z;
		19'b0010000000110100100: color_data = Z;
		19'b0010000000110100101: color_data = Z;
		19'b0010000000110100110: color_data = Z;
		19'b0010000000110100111: color_data = Z;
		19'b0010000000110101000: color_data = Z;
		19'b0010000000110101100: color_data = Z;
		19'b0010000000110101101: color_data = Z;
		19'b0010000000110101110: color_data = Z;
		19'b0010000000110101111: color_data = Z;
		19'b0010000000110110000: color_data = Z;
		19'b0010000000110110001: color_data = Z;
		19'b0010000000110110110: color_data = Z;
		19'b0010000000110110111: color_data = Z;
		19'b0010000000110111000: color_data = Z;
		19'b0010000000110111001: color_data = Z;
		19'b0010000000110111010: color_data = Z;
		19'b0010000000110111011: color_data = Z;
		19'b0010000000110111100: color_data = Z;
		19'b0010000000110111101: color_data = Z;
		19'b0010000000110111110: color_data = Z;
		19'b0010000000110111111: color_data = Z;
		19'b0010000000111000000: color_data = Z;
		19'b0010000000111000001: color_data = Z;
		19'b0010000000111000010: color_data = Z;
		19'b0010000010011010000: color_data = Z;
		19'b0010000010011010001: color_data = Z;
		19'b0010000010011010010: color_data = Z;
		19'b0010000010011010011: color_data = Z;
		19'b0010000010011010100: color_data = Z;
		19'b0010000010011010101: color_data = Z;
		19'b0010000010011010110: color_data = Z;
		19'b0010000010011010111: color_data = Z;
		19'b0010000010011011000: color_data = Z;
		19'b0010000010011011001: color_data = Z;
		19'b0010000010011011010: color_data = Z;
		19'b0010000010011011011: color_data = Z;
		19'b0010000010011011100: color_data = Z;
		19'b0010000010011011101: color_data = Z;
		19'b0010000010011011110: color_data = Z;
		19'b0010000010011011111: color_data = Z;
		19'b0010000010011100000: color_data = Z;
		19'b0010000010011100001: color_data = Z;
		19'b0010000010011100010: color_data = Z;
		19'b0010000010011100011: color_data = Z;
		19'b0010000010011100100: color_data = Z;
		19'b0010000010011100101: color_data = Z;
		19'b0010000010011100110: color_data = Z;
		19'b0010000010011100111: color_data = Z;
		19'b0010000010011101000: color_data = Z;
		19'b0010000010011101001: color_data = Z;
		19'b0010000010011101010: color_data = Z;
		19'b0010000010011101011: color_data = Z;
		19'b0010000010011101100: color_data = Z;
		19'b0010000010011101101: color_data = Z;
		19'b0010000010011101110: color_data = Z;
		19'b0010000010011101111: color_data = Z;
		19'b0010000010011110000: color_data = Z;
		19'b0010000010011110001: color_data = Z;
		19'b0010000010011110010: color_data = Z;
		19'b0010000010011110011: color_data = Z;
		19'b0010000010011110100: color_data = Z;
		19'b0010000010011110101: color_data = Z;
		19'b0010000010011110110: color_data = Z;
		19'b0010000010011110111: color_data = Z;
		19'b0010000010011111000: color_data = Z;
		19'b0010000010011111001: color_data = Z;
		19'b0010000010011111010: color_data = Z;
		19'b0010000010011111011: color_data = Z;
		19'b0010000010011111100: color_data = Z;
		19'b0010000010011111101: color_data = Z;
		19'b0010000010011111110: color_data = Z;
		19'b0010000010011111111: color_data = Z;
		19'b0010000010100000000: color_data = Z;
		19'b0010000010100000001: color_data = Z;
		19'b0010000010100000010: color_data = Z;
		19'b0010000010100000011: color_data = Z;
		19'b0010000010100000100: color_data = Z;
		19'b0010000010100000101: color_data = Z;
		19'b0010000010100000110: color_data = Z;
		19'b0010000010100000111: color_data = Z;
		19'b0010000010100001000: color_data = Z;
		19'b0010000010100001001: color_data = Z;
		19'b0010000010100001010: color_data = Z;
		19'b0010000010100001011: color_data = Z;
		19'b0010000010100001100: color_data = Z;
		19'b0010000010100001101: color_data = Z;
		19'b0010000010100001110: color_data = Z;
		19'b0010000010100001111: color_data = Z;
		19'b0010000010100010000: color_data = Z;
		19'b0010000010100010001: color_data = Z;
		19'b0010000010100010010: color_data = Z;
		19'b0010000010100010011: color_data = Z;
		19'b0010000010100010100: color_data = Z;
		19'b0010000010100010101: color_data = Z;
		19'b0010000010100010110: color_data = Z;
		19'b0010000010100010111: color_data = Z;
		19'b0010000010100011000: color_data = Z;
		19'b0010000010100011001: color_data = Z;
		19'b0010000010100011010: color_data = Z;
		19'b0010000010100011011: color_data = Z;
		19'b0010000010100011100: color_data = Z;
		19'b0010000010100011101: color_data = Z;
		19'b0010000010100011110: color_data = Z;
		19'b0010000010100011111: color_data = Z;
		19'b0010000010100100000: color_data = Z;
		19'b0010000010100100001: color_data = Z;
		19'b0010000010100100010: color_data = Z;
		19'b0010000010100100011: color_data = Z;
		19'b0010000010100100100: color_data = Z;
		19'b0010000010100100101: color_data = Z;
		19'b0010000010100100110: color_data = Z;
		19'b0010000010100100111: color_data = Z;
		19'b0010000010100101000: color_data = Z;
		19'b0010000010100101001: color_data = Z;
		19'b0010000010100101010: color_data = Z;
		19'b0010000010100101011: color_data = Z;
		19'b0010000010100101100: color_data = Z;
		19'b0010000010100101101: color_data = Z;
		19'b0010000010100101110: color_data = Z;
		19'b0010000010100101111: color_data = Z;
		19'b0010000010100110000: color_data = Z;
		19'b0010000010100110001: color_data = Z;
		19'b0010000010100110010: color_data = Z;
		19'b0010000010100110011: color_data = Z;
		19'b0010000010100110100: color_data = Z;
		19'b0010000010100110101: color_data = Z;
		19'b0010000010100110110: color_data = Z;
		19'b0010000010100110111: color_data = Z;
		19'b0010000010100111000: color_data = Z;
		19'b0010000010100111001: color_data = Z;
		19'b0010000010100111010: color_data = Z;
		19'b0010000010100111011: color_data = Z;
		19'b0010000010100111100: color_data = Z;
		19'b0010000010100111101: color_data = Z;
		19'b0010000010100111110: color_data = Z;
		19'b0010000010100111111: color_data = Z;
		19'b0010000010101000000: color_data = Z;
		19'b0010000010101000001: color_data = Z;
		19'b0010000010101000010: color_data = Z;
		19'b0010000010101000011: color_data = Z;
		19'b0010000010101000100: color_data = Z;
		19'b0010000010101000101: color_data = Z;
		19'b0010000010101000110: color_data = Z;
		19'b0010000010101000111: color_data = Z;
		19'b0010000010101001000: color_data = Z;
		19'b0010000010101001001: color_data = Z;
		19'b0010000010101001010: color_data = Z;
		19'b0010000010101001011: color_data = Z;
		19'b0010000010101001100: color_data = Z;
		19'b0010000010101001101: color_data = Z;
		19'b0010000010101001110: color_data = Z;
		19'b0010000010101001111: color_data = Z;
		19'b0010000010101010000: color_data = Z;
		19'b0010000010101010001: color_data = Z;
		19'b0010000010101010010: color_data = Z;
		19'b0010000010101010011: color_data = Z;
		19'b0010000010101010100: color_data = Z;
		19'b0010000010101010101: color_data = Z;
		19'b0010000010101010110: color_data = Z;
		19'b0010000010101010111: color_data = Z;
		19'b0010000010101011000: color_data = Z;
		19'b0010000010101011001: color_data = Z;
		19'b0010000010101011010: color_data = Z;
		19'b0010000010101011011: color_data = Z;
		19'b0010000010101011100: color_data = Z;
		19'b0010000010101011101: color_data = Z;
		19'b0010000010101011110: color_data = Z;
		19'b0010000010101011111: color_data = Z;
		19'b0010000010101100000: color_data = Z;
		19'b0010000010101100001: color_data = Z;
		19'b0010000010101100010: color_data = Z;
		19'b0010000010101100011: color_data = Z;
		19'b0010000010101100100: color_data = Z;
		19'b0010000010101100101: color_data = Z;
		19'b0010000010101100110: color_data = Z;
		19'b0010000010101100111: color_data = Z;
		19'b0010000010101101000: color_data = Z;
		19'b0010000010101101001: color_data = Z;
		19'b0010000010101101010: color_data = Z;
		19'b0010000010101101011: color_data = Z;
		19'b0010000010101101100: color_data = Z;
		19'b0010000010101101101: color_data = Z;
		19'b0010000010101101110: color_data = Z;
		19'b0010000010101101111: color_data = Z;
		19'b0010000010101110000: color_data = Z;
		19'b0010000010101110001: color_data = Z;
		19'b0010000010101110010: color_data = Z;
		19'b0010000010101110011: color_data = Z;
		19'b0010000010101110100: color_data = Z;
		19'b0010000010101110101: color_data = Z;
		19'b0010000010101110110: color_data = Z;
		19'b0010000010101110111: color_data = Z;
		19'b0010000010101111000: color_data = Z;
		19'b0010000010101111001: color_data = Z;
		19'b0010000010101111010: color_data = Z;
		19'b0010000010101111011: color_data = Z;
		19'b0010000010101111100: color_data = Z;
		19'b0010000010101111101: color_data = Z;
		19'b0010000010101111110: color_data = Z;
		19'b0010000010101111111: color_data = Z;
		19'b0010000010110000000: color_data = Z;
		19'b0010000010110000001: color_data = Z;
		19'b0010000010110000010: color_data = Z;
		19'b0010000010110000011: color_data = Z;
		19'b0010000010110000100: color_data = Z;
		19'b0010000010110000101: color_data = Z;
		19'b0010000010110000110: color_data = Z;
		19'b0010000010110000111: color_data = Z;
		19'b0010000010110001000: color_data = Z;
		19'b0010000010110001001: color_data = Z;
		19'b0010000010110001010: color_data = Z;
		19'b0010000010110001011: color_data = Z;
		19'b0010000010110001100: color_data = Z;
		19'b0010000010110001101: color_data = Z;
		19'b0010000010110001110: color_data = Z;
		19'b0010000010110001111: color_data = Z;
		19'b0010000010110010000: color_data = Z;
		19'b0010000010110010001: color_data = Z;
		19'b0010000010110010010: color_data = Z;
		19'b0010000010110010011: color_data = Z;
		19'b0010000010110010100: color_data = Z;
		19'b0010000010110010101: color_data = Z;
		19'b0010000010110010110: color_data = Z;
		19'b0010000010110010111: color_data = Z;
		19'b0010000010110011000: color_data = Z;
		19'b0010000010110011001: color_data = Z;
		19'b0010000010110011010: color_data = Z;
		19'b0010000010110011011: color_data = Z;
		19'b0010000010110011100: color_data = Z;
		19'b0010000010110011101: color_data = Z;
		19'b0010000010110011110: color_data = Z;
		19'b0010000010110011111: color_data = Z;
		19'b0010000010110100000: color_data = Z;
		19'b0010000010110100001: color_data = Z;
		19'b0010000010110100010: color_data = Z;
		19'b0010000010110100011: color_data = Z;
		19'b0010000010110100100: color_data = Z;
		19'b0010000010110100101: color_data = Z;
		19'b0010000010110100110: color_data = Z;
		19'b0010000010110100111: color_data = Z;
		19'b0010000010110101000: color_data = Z;
		19'b0010000010110101100: color_data = Z;
		19'b0010000010110101101: color_data = Z;
		19'b0010000010110101110: color_data = Z;
		19'b0010000010110101111: color_data = Z;
		19'b0010000010110110000: color_data = Z;
		19'b0010000010110110001: color_data = Z;
		19'b0010000010110110111: color_data = Z;
		19'b0010000010110111000: color_data = Z;
		19'b0010000010110111001: color_data = Z;
		19'b0010000010110111010: color_data = Z;
		19'b0010000010110111011: color_data = Z;
		19'b0010000010110111100: color_data = Z;
		19'b0010000010110111101: color_data = Z;
		19'b0010000010110111110: color_data = Z;
		19'b0010000010110111111: color_data = Z;
		19'b0010000010111000000: color_data = Z;
		19'b0010000010111000001: color_data = Z;
		19'b0010000010111000010: color_data = Z;
		19'b0010000010111000011: color_data = Z;
		19'b0010000100011001111: color_data = Z;
		19'b0010000100011010000: color_data = Z;
		19'b0010000100011010001: color_data = Z;
		19'b0010000100011010010: color_data = Z;
		19'b0010000100011010011: color_data = Z;
		19'b0010000100011010100: color_data = Z;
		19'b0010000100011010101: color_data = Z;
		19'b0010000100011010110: color_data = Z;
		19'b0010000100011010111: color_data = Z;
		19'b0010000100011011000: color_data = Z;
		19'b0010000100011011001: color_data = Z;
		19'b0010000100011011010: color_data = Z;
		19'b0010000100011011011: color_data = Z;
		19'b0010000100011011100: color_data = Z;
		19'b0010000100011011101: color_data = Z;
		19'b0010000100011011110: color_data = Z;
		19'b0010000100011011111: color_data = Z;
		19'b0010000100011100000: color_data = Z;
		19'b0010000100011100001: color_data = Z;
		19'b0010000100011100010: color_data = Z;
		19'b0010000100011100011: color_data = Z;
		19'b0010000100011100100: color_data = Z;
		19'b0010000100011100101: color_data = Z;
		19'b0010000100011100110: color_data = Z;
		19'b0010000100011100111: color_data = Z;
		19'b0010000100011101000: color_data = Z;
		19'b0010000100011101001: color_data = Z;
		19'b0010000100011101010: color_data = Z;
		19'b0010000100011101011: color_data = Z;
		19'b0010000100011101100: color_data = Z;
		19'b0010000100011101101: color_data = Z;
		19'b0010000100011101110: color_data = Z;
		19'b0010000100011101111: color_data = Z;
		19'b0010000100011110000: color_data = Z;
		19'b0010000100011110001: color_data = Z;
		19'b0010000100011110010: color_data = Z;
		19'b0010000100011110011: color_data = Z;
		19'b0010000100011110100: color_data = Z;
		19'b0010000100011110101: color_data = Z;
		19'b0010000100011110110: color_data = Z;
		19'b0010000100011110111: color_data = Z;
		19'b0010000100011111000: color_data = Z;
		19'b0010000100011111001: color_data = Z;
		19'b0010000100011111010: color_data = Z;
		19'b0010000100011111011: color_data = Z;
		19'b0010000100011111100: color_data = Z;
		19'b0010000100011111101: color_data = Z;
		19'b0010000100011111110: color_data = Z;
		19'b0010000100011111111: color_data = Z;
		19'b0010000100100000000: color_data = Z;
		19'b0010000100100000001: color_data = Z;
		19'b0010000100100000010: color_data = Z;
		19'b0010000100100000011: color_data = Z;
		19'b0010000100100000100: color_data = Z;
		19'b0010000100100000101: color_data = Z;
		19'b0010000100100000110: color_data = Z;
		19'b0010000100100000111: color_data = Z;
		19'b0010000100100001000: color_data = Z;
		19'b0010000100100001001: color_data = Z;
		19'b0010000100100001010: color_data = Z;
		19'b0010000100100001011: color_data = Z;
		19'b0010000100100001100: color_data = Z;
		19'b0010000100100001101: color_data = Z;
		19'b0010000100100001110: color_data = Z;
		19'b0010000100100001111: color_data = Z;
		19'b0010000100100010000: color_data = Z;
		19'b0010000100100010001: color_data = Z;
		19'b0010000100100010010: color_data = Z;
		19'b0010000100100010011: color_data = Z;
		19'b0010000100100010100: color_data = Z;
		19'b0010000100100010101: color_data = Z;
		19'b0010000100100010110: color_data = Z;
		19'b0010000100100010111: color_data = Z;
		19'b0010000100100011000: color_data = Z;
		19'b0010000100100011001: color_data = Z;
		19'b0010000100100011010: color_data = Z;
		19'b0010000100100011011: color_data = Z;
		19'b0010000100100011100: color_data = Z;
		19'b0010000100100011101: color_data = Z;
		19'b0010000100100011110: color_data = Z;
		19'b0010000100100011111: color_data = Z;
		19'b0010000100100100000: color_data = Z;
		19'b0010000100100100001: color_data = Z;
		19'b0010000100100100010: color_data = Z;
		19'b0010000100100100011: color_data = Z;
		19'b0010000100100100100: color_data = Z;
		19'b0010000100100100101: color_data = Z;
		19'b0010000100100100110: color_data = Z;
		19'b0010000100100100111: color_data = Z;
		19'b0010000100100101000: color_data = Z;
		19'b0010000100100101001: color_data = Z;
		19'b0010000100100101010: color_data = Z;
		19'b0010000100100101011: color_data = Z;
		19'b0010000100100101100: color_data = Z;
		19'b0010000100100101101: color_data = Z;
		19'b0010000100100101110: color_data = Z;
		19'b0010000100100101111: color_data = Z;
		19'b0010000100100110000: color_data = Z;
		19'b0010000100100110001: color_data = Z;
		19'b0010000100100110010: color_data = Z;
		19'b0010000100100110011: color_data = Z;
		19'b0010000100100110100: color_data = Z;
		19'b0010000100100110101: color_data = Z;
		19'b0010000100100110110: color_data = Z;
		19'b0010000100100110111: color_data = Z;
		19'b0010000100100111000: color_data = Z;
		19'b0010000100100111001: color_data = Z;
		19'b0010000100100111010: color_data = Z;
		19'b0010000100100111011: color_data = Z;
		19'b0010000100100111100: color_data = Z;
		19'b0010000100100111101: color_data = Z;
		19'b0010000100100111110: color_data = Z;
		19'b0010000100100111111: color_data = Z;
		19'b0010000100101000000: color_data = Z;
		19'b0010000100101000001: color_data = Z;
		19'b0010000100101000010: color_data = Z;
		19'b0010000100101000011: color_data = Z;
		19'b0010000100101000100: color_data = Z;
		19'b0010000100101000101: color_data = Z;
		19'b0010000100101000110: color_data = Z;
		19'b0010000100101000111: color_data = Z;
		19'b0010000100101001000: color_data = Z;
		19'b0010000100101001001: color_data = Z;
		19'b0010000100101001010: color_data = Z;
		19'b0010000100101001011: color_data = Z;
		19'b0010000100101001100: color_data = Z;
		19'b0010000100101001101: color_data = Z;
		19'b0010000100101001110: color_data = Z;
		19'b0010000100101001111: color_data = Z;
		19'b0010000100101010000: color_data = Z;
		19'b0010000100101010001: color_data = Z;
		19'b0010000100101010010: color_data = Z;
		19'b0010000100101010011: color_data = Z;
		19'b0010000100101010100: color_data = Z;
		19'b0010000100101010101: color_data = Z;
		19'b0010000100101010110: color_data = Z;
		19'b0010000100101010111: color_data = Z;
		19'b0010000100101011000: color_data = Z;
		19'b0010000100101011001: color_data = Z;
		19'b0010000100101011010: color_data = Z;
		19'b0010000100101011011: color_data = Z;
		19'b0010000100101011100: color_data = Z;
		19'b0010000100101011101: color_data = Z;
		19'b0010000100101011110: color_data = Z;
		19'b0010000100101011111: color_data = Z;
		19'b0010000100101100000: color_data = Z;
		19'b0010000100101100001: color_data = Z;
		19'b0010000100101100010: color_data = Z;
		19'b0010000100101100011: color_data = Z;
		19'b0010000100101100100: color_data = Z;
		19'b0010000100101100101: color_data = Z;
		19'b0010000100101100110: color_data = Z;
		19'b0010000100101100111: color_data = Z;
		19'b0010000100101101000: color_data = Z;
		19'b0010000100101101001: color_data = Z;
		19'b0010000100101101010: color_data = Z;
		19'b0010000100101101011: color_data = Z;
		19'b0010000100101101100: color_data = Z;
		19'b0010000100101101101: color_data = Z;
		19'b0010000100101101110: color_data = Z;
		19'b0010000100101101111: color_data = Z;
		19'b0010000100101110000: color_data = Z;
		19'b0010000100101110001: color_data = Z;
		19'b0010000100101110010: color_data = Z;
		19'b0010000100101110011: color_data = Z;
		19'b0010000100101110100: color_data = Z;
		19'b0010000100101110101: color_data = Z;
		19'b0010000100101110110: color_data = Z;
		19'b0010000100101110111: color_data = Z;
		19'b0010000100101111000: color_data = Z;
		19'b0010000100101111001: color_data = Z;
		19'b0010000100101111010: color_data = Z;
		19'b0010000100101111011: color_data = Z;
		19'b0010000100101111100: color_data = Z;
		19'b0010000100101111101: color_data = Z;
		19'b0010000100101111110: color_data = Z;
		19'b0010000100101111111: color_data = Z;
		19'b0010000100110000000: color_data = Z;
		19'b0010000100110000001: color_data = Z;
		19'b0010000100110000010: color_data = Z;
		19'b0010000100110000011: color_data = Z;
		19'b0010000100110000100: color_data = Z;
		19'b0010000100110000101: color_data = Z;
		19'b0010000100110000110: color_data = Z;
		19'b0010000100110000111: color_data = Z;
		19'b0010000100110001000: color_data = Z;
		19'b0010000100110001001: color_data = Z;
		19'b0010000100110001010: color_data = Z;
		19'b0010000100110001011: color_data = Z;
		19'b0010000100110001100: color_data = Z;
		19'b0010000100110001101: color_data = Z;
		19'b0010000100110001110: color_data = Z;
		19'b0010000100110001111: color_data = Z;
		19'b0010000100110010000: color_data = Z;
		19'b0010000100110010001: color_data = Z;
		19'b0010000100110010010: color_data = Z;
		19'b0010000100110010011: color_data = Z;
		19'b0010000100110010100: color_data = Z;
		19'b0010000100110010101: color_data = Z;
		19'b0010000100110010110: color_data = Z;
		19'b0010000100110010111: color_data = Z;
		19'b0010000100110011000: color_data = Z;
		19'b0010000100110011001: color_data = Z;
		19'b0010000100110011010: color_data = Z;
		19'b0010000100110011011: color_data = Z;
		19'b0010000100110011100: color_data = Z;
		19'b0010000100110011101: color_data = Z;
		19'b0010000100110011110: color_data = Z;
		19'b0010000100110011111: color_data = Z;
		19'b0010000100110100000: color_data = Z;
		19'b0010000100110100001: color_data = Z;
		19'b0010000100110100010: color_data = Z;
		19'b0010000100110100011: color_data = Z;
		19'b0010000100110100100: color_data = Z;
		19'b0010000100110100101: color_data = Z;
		19'b0010000100110100110: color_data = Z;
		19'b0010000100110100111: color_data = Z;
		19'b0010000100110101000: color_data = Z;
		19'b0010000100110101001: color_data = Z;
		19'b0010000100110101101: color_data = Z;
		19'b0010000100110101110: color_data = Z;
		19'b0010000100110101111: color_data = Z;
		19'b0010000100110110000: color_data = Z;
		19'b0010000100110110001: color_data = Z;
		19'b0010000100110110010: color_data = Z;
		19'b0010000100110110111: color_data = Z;
		19'b0010000100110111000: color_data = Z;
		19'b0010000100110111001: color_data = Z;
		19'b0010000100110111010: color_data = Z;
		19'b0010000100110111011: color_data = Z;
		19'b0010000100110111100: color_data = Z;
		19'b0010000100110111101: color_data = Z;
		19'b0010000100110111110: color_data = Z;
		19'b0010000100110111111: color_data = Z;
		19'b0010000100111000000: color_data = Z;
		19'b0010000100111000001: color_data = Z;
		19'b0010000100111000010: color_data = Z;
		19'b0010000100111000011: color_data = Z;
		19'b0010000110011001110: color_data = Z;
		19'b0010000110011001111: color_data = Z;
		19'b0010000110011010000: color_data = Z;
		19'b0010000110011010001: color_data = Z;
		19'b0010000110011010010: color_data = Z;
		19'b0010000110011010011: color_data = Z;
		19'b0010000110011010100: color_data = Z;
		19'b0010000110011010101: color_data = Z;
		19'b0010000110011010110: color_data = Z;
		19'b0010000110011010111: color_data = Z;
		19'b0010000110011011000: color_data = Z;
		19'b0010000110011011001: color_data = Z;
		19'b0010000110011011010: color_data = Z;
		19'b0010000110011011011: color_data = Z;
		19'b0010000110011011100: color_data = Z;
		19'b0010000110011011101: color_data = Z;
		19'b0010000110011011110: color_data = Z;
		19'b0010000110011011111: color_data = Z;
		19'b0010000110011100000: color_data = Z;
		19'b0010000110011100001: color_data = Z;
		19'b0010000110011100010: color_data = Z;
		19'b0010000110011100011: color_data = Z;
		19'b0010000110011100100: color_data = Z;
		19'b0010000110011100101: color_data = Z;
		19'b0010000110011100110: color_data = Z;
		19'b0010000110011100111: color_data = Z;
		19'b0010000110011101000: color_data = Z;
		19'b0010000110011101001: color_data = Z;
		19'b0010000110011101010: color_data = Z;
		19'b0010000110011101011: color_data = Z;
		19'b0010000110011101100: color_data = Z;
		19'b0010000110011101101: color_data = Z;
		19'b0010000110011101110: color_data = Z;
		19'b0010000110011101111: color_data = Z;
		19'b0010000110011110000: color_data = Z;
		19'b0010000110011110001: color_data = Z;
		19'b0010000110011110010: color_data = Z;
		19'b0010000110011110011: color_data = Z;
		19'b0010000110011110100: color_data = Z;
		19'b0010000110011110101: color_data = Z;
		19'b0010000110011110110: color_data = Z;
		19'b0010000110011110111: color_data = Z;
		19'b0010000110011111000: color_data = Z;
		19'b0010000110011111001: color_data = Z;
		19'b0010000110011111010: color_data = Z;
		19'b0010000110011111011: color_data = Z;
		19'b0010000110011111100: color_data = Z;
		19'b0010000110011111101: color_data = Z;
		19'b0010000110011111110: color_data = Z;
		19'b0010000110011111111: color_data = Z;
		19'b0010000110100000000: color_data = Z;
		19'b0010000110100000001: color_data = Z;
		19'b0010000110100000010: color_data = Z;
		19'b0010000110100000011: color_data = Z;
		19'b0010000110100000100: color_data = Z;
		19'b0010000110100000101: color_data = Z;
		19'b0010000110100000110: color_data = Z;
		19'b0010000110100000111: color_data = Z;
		19'b0010000110100001000: color_data = Z;
		19'b0010000110100001001: color_data = Z;
		19'b0010000110100001010: color_data = Z;
		19'b0010000110100001011: color_data = Z;
		19'b0010000110100001100: color_data = Z;
		19'b0010000110100001101: color_data = Z;
		19'b0010000110100001110: color_data = Z;
		19'b0010000110100001111: color_data = Z;
		19'b0010000110100010000: color_data = Z;
		19'b0010000110100010001: color_data = Z;
		19'b0010000110100010010: color_data = Z;
		19'b0010000110100010011: color_data = Z;
		19'b0010000110100010100: color_data = Z;
		19'b0010000110100010101: color_data = Z;
		19'b0010000110100010110: color_data = Z;
		19'b0010000110100010111: color_data = Z;
		19'b0010000110100011000: color_data = Z;
		19'b0010000110100011001: color_data = Z;
		19'b0010000110100011010: color_data = Z;
		19'b0010000110100011011: color_data = Z;
		19'b0010000110100011100: color_data = Z;
		19'b0010000110100011101: color_data = Z;
		19'b0010000110100011110: color_data = Z;
		19'b0010000110100011111: color_data = Z;
		19'b0010000110100100000: color_data = Z;
		19'b0010000110100100001: color_data = Z;
		19'b0010000110100100010: color_data = Z;
		19'b0010000110100100011: color_data = Z;
		19'b0010000110100100100: color_data = Z;
		19'b0010000110100100101: color_data = Z;
		19'b0010000110100100110: color_data = Z;
		19'b0010000110100100111: color_data = Z;
		19'b0010000110100101000: color_data = Z;
		19'b0010000110100101001: color_data = Z;
		19'b0010000110100101010: color_data = Z;
		19'b0010000110100101011: color_data = Z;
		19'b0010000110100101100: color_data = Z;
		19'b0010000110100101101: color_data = Z;
		19'b0010000110100101110: color_data = Z;
		19'b0010000110100101111: color_data = Z;
		19'b0010000110100110000: color_data = Z;
		19'b0010000110100110001: color_data = Z;
		19'b0010000110100110010: color_data = Z;
		19'b0010000110100110011: color_data = Z;
		19'b0010000110100110100: color_data = Z;
		19'b0010000110100110101: color_data = Z;
		19'b0010000110100110110: color_data = Z;
		19'b0010000110100110111: color_data = Z;
		19'b0010000110100111000: color_data = Z;
		19'b0010000110100111001: color_data = Z;
		19'b0010000110100111010: color_data = Z;
		19'b0010000110100111011: color_data = Z;
		19'b0010000110100111100: color_data = Z;
		19'b0010000110100111101: color_data = Z;
		19'b0010000110100111110: color_data = Z;
		19'b0010000110100111111: color_data = Z;
		19'b0010000110101000000: color_data = Z;
		19'b0010000110101000001: color_data = Z;
		19'b0010000110101000010: color_data = Z;
		19'b0010000110101000011: color_data = Z;
		19'b0010000110101000100: color_data = Z;
		19'b0010000110101000101: color_data = Z;
		19'b0010000110101000110: color_data = Z;
		19'b0010000110101000111: color_data = Z;
		19'b0010000110101001000: color_data = Z;
		19'b0010000110101001001: color_data = Z;
		19'b0010000110101001010: color_data = Z;
		19'b0010000110101001011: color_data = Z;
		19'b0010000110101001100: color_data = Z;
		19'b0010000110101001101: color_data = Z;
		19'b0010000110101001110: color_data = Z;
		19'b0010000110101001111: color_data = Z;
		19'b0010000110101010000: color_data = Z;
		19'b0010000110101010001: color_data = Z;
		19'b0010000110101010010: color_data = Z;
		19'b0010000110101010011: color_data = Z;
		19'b0010000110101010100: color_data = Z;
		19'b0010000110101010101: color_data = Z;
		19'b0010000110101010110: color_data = Z;
		19'b0010000110101010111: color_data = Z;
		19'b0010000110101011000: color_data = Z;
		19'b0010000110101011001: color_data = Z;
		19'b0010000110101011010: color_data = Z;
		19'b0010000110101011011: color_data = Z;
		19'b0010000110101011100: color_data = Z;
		19'b0010000110101011101: color_data = Z;
		19'b0010000110101011110: color_data = Z;
		19'b0010000110101011111: color_data = Z;
		19'b0010000110101100000: color_data = Z;
		19'b0010000110101100001: color_data = Z;
		19'b0010000110101100010: color_data = Z;
		19'b0010000110101100011: color_data = Z;
		19'b0010000110101100100: color_data = Z;
		19'b0010000110101100101: color_data = Z;
		19'b0010000110101100110: color_data = Z;
		19'b0010000110101100111: color_data = Z;
		19'b0010000110101101000: color_data = Z;
		19'b0010000110101101001: color_data = Z;
		19'b0010000110101101010: color_data = Z;
		19'b0010000110101101011: color_data = Z;
		19'b0010000110101101100: color_data = Z;
		19'b0010000110101101101: color_data = Z;
		19'b0010000110101101110: color_data = Z;
		19'b0010000110101101111: color_data = Z;
		19'b0010000110101110000: color_data = Z;
		19'b0010000110101110001: color_data = Z;
		19'b0010000110101110010: color_data = Z;
		19'b0010000110101110011: color_data = Z;
		19'b0010000110101110100: color_data = Z;
		19'b0010000110101110101: color_data = Z;
		19'b0010000110101110110: color_data = Z;
		19'b0010000110101110111: color_data = Z;
		19'b0010000110101111000: color_data = Z;
		19'b0010000110101111001: color_data = Z;
		19'b0010000110101111010: color_data = Z;
		19'b0010000110101111011: color_data = Z;
		19'b0010000110101111100: color_data = Z;
		19'b0010000110101111101: color_data = Z;
		19'b0010000110101111110: color_data = Z;
		19'b0010000110101111111: color_data = Z;
		19'b0010000110110000000: color_data = Z;
		19'b0010000110110000001: color_data = Z;
		19'b0010000110110000010: color_data = Z;
		19'b0010000110110000011: color_data = Z;
		19'b0010000110110000100: color_data = Z;
		19'b0010000110110000101: color_data = Z;
		19'b0010000110110000110: color_data = Z;
		19'b0010000110110000111: color_data = Z;
		19'b0010000110110001000: color_data = Z;
		19'b0010000110110001001: color_data = Z;
		19'b0010000110110001010: color_data = Z;
		19'b0010000110110001011: color_data = Z;
		19'b0010000110110001100: color_data = Z;
		19'b0010000110110001101: color_data = Z;
		19'b0010000110110001110: color_data = Z;
		19'b0010000110110001111: color_data = Z;
		19'b0010000110110010000: color_data = Z;
		19'b0010000110110010001: color_data = Z;
		19'b0010000110110010010: color_data = Z;
		19'b0010000110110010011: color_data = Z;
		19'b0010000110110010100: color_data = Z;
		19'b0010000110110010101: color_data = Z;
		19'b0010000110110010110: color_data = Z;
		19'b0010000110110010111: color_data = Z;
		19'b0010000110110011000: color_data = Z;
		19'b0010000110110011001: color_data = Z;
		19'b0010000110110011010: color_data = Z;
		19'b0010000110110011011: color_data = Z;
		19'b0010000110110011100: color_data = Z;
		19'b0010000110110011101: color_data = Z;
		19'b0010000110110011110: color_data = Z;
		19'b0010000110110011111: color_data = Z;
		19'b0010000110110100000: color_data = Z;
		19'b0010000110110100001: color_data = Z;
		19'b0010000110110100010: color_data = Z;
		19'b0010000110110100011: color_data = Z;
		19'b0010000110110100100: color_data = Z;
		19'b0010000110110100101: color_data = Z;
		19'b0010000110110100110: color_data = Z;
		19'b0010000110110100111: color_data = Z;
		19'b0010000110110101000: color_data = Z;
		19'b0010000110110101001: color_data = Z;
		19'b0010000110110101101: color_data = Z;
		19'b0010000110110101110: color_data = Z;
		19'b0010000110110101111: color_data = Z;
		19'b0010000110110110000: color_data = Z;
		19'b0010000110110110001: color_data = Z;
		19'b0010000110110110010: color_data = Z;
		19'b0010000110110111000: color_data = Z;
		19'b0010000110110111001: color_data = Z;
		19'b0010000110110111010: color_data = Z;
		19'b0010000110110111011: color_data = Z;
		19'b0010000110110111100: color_data = Z;
		19'b0010000110110111101: color_data = Z;
		19'b0010000110110111110: color_data = Z;
		19'b0010000110110111111: color_data = Z;
		19'b0010000110111000000: color_data = Z;
		19'b0010000110111000001: color_data = Z;
		19'b0010000110111000010: color_data = Z;
		19'b0010000110111000011: color_data = Z;
		19'b0010001000011001110: color_data = Z;
		19'b0010001000011001111: color_data = Z;
		19'b0010001000011010000: color_data = Z;
		19'b0010001000011010001: color_data = Z;
		19'b0010001000011010010: color_data = Z;
		19'b0010001000011010011: color_data = Z;
		19'b0010001000011010100: color_data = Z;
		19'b0010001000011010101: color_data = Z;
		19'b0010001000011010110: color_data = Z;
		19'b0010001000011010111: color_data = Z;
		19'b0010001000011011000: color_data = Z;
		19'b0010001000011011001: color_data = Z;
		19'b0010001000011011010: color_data = Z;
		19'b0010001000011011011: color_data = Z;
		19'b0010001000011011100: color_data = Z;
		19'b0010001000011011101: color_data = Z;
		19'b0010001000011011110: color_data = Z;
		19'b0010001000011011111: color_data = Z;
		19'b0010001000011100000: color_data = Z;
		19'b0010001000011100001: color_data = Z;
		19'b0010001000011100010: color_data = Z;
		19'b0010001000011100011: color_data = Z;
		19'b0010001000011100100: color_data = Z;
		19'b0010001000011100101: color_data = Z;
		19'b0010001000011100110: color_data = Z;
		19'b0010001000011100111: color_data = Z;
		19'b0010001000011101000: color_data = Z;
		19'b0010001000011101001: color_data = Z;
		19'b0010001000011101010: color_data = Z;
		19'b0010001000011101011: color_data = Z;
		19'b0010001000011101100: color_data = Z;
		19'b0010001000011101101: color_data = Z;
		19'b0010001000011101110: color_data = Z;
		19'b0010001000011101111: color_data = Z;
		19'b0010001000011110000: color_data = Z;
		19'b0010001000011110001: color_data = Z;
		19'b0010001000011110010: color_data = Z;
		19'b0010001000011110011: color_data = Z;
		19'b0010001000011110100: color_data = Z;
		19'b0010001000011110101: color_data = Z;
		19'b0010001000011110110: color_data = Z;
		19'b0010001000011110111: color_data = Z;
		19'b0010001000011111000: color_data = Z;
		19'b0010001000011111001: color_data = Z;
		19'b0010001000011111010: color_data = Z;
		19'b0010001000011111011: color_data = Z;
		19'b0010001000011111100: color_data = Z;
		19'b0010001000011111101: color_data = Z;
		19'b0010001000011111110: color_data = Z;
		19'b0010001000011111111: color_data = Z;
		19'b0010001000100000000: color_data = Z;
		19'b0010001000100000001: color_data = Z;
		19'b0010001000100000010: color_data = Z;
		19'b0010001000100000011: color_data = Z;
		19'b0010001000100000100: color_data = Z;
		19'b0010001000100000101: color_data = Z;
		19'b0010001000100000110: color_data = Z;
		19'b0010001000100000111: color_data = Z;
		19'b0010001000100001000: color_data = Z;
		19'b0010001000100001001: color_data = Z;
		19'b0010001000100001010: color_data = Z;
		19'b0010001000100001011: color_data = Z;
		19'b0010001000100001100: color_data = Z;
		19'b0010001000100001101: color_data = Z;
		19'b0010001000100001110: color_data = Z;
		19'b0010001000100001111: color_data = Z;
		19'b0010001000100010000: color_data = Z;
		19'b0010001000100010001: color_data = Z;
		19'b0010001000100010010: color_data = Z;
		19'b0010001000100010011: color_data = Z;
		19'b0010001000100010100: color_data = Z;
		19'b0010001000100010101: color_data = Z;
		19'b0010001000100010110: color_data = Z;
		19'b0010001000100010111: color_data = Z;
		19'b0010001000100011000: color_data = Z;
		19'b0010001000100011001: color_data = Z;
		19'b0010001000100011010: color_data = Z;
		19'b0010001000100011011: color_data = Z;
		19'b0010001000100011100: color_data = Z;
		19'b0010001000100011101: color_data = Z;
		19'b0010001000100011110: color_data = Z;
		19'b0010001000100011111: color_data = Z;
		19'b0010001000100100000: color_data = Z;
		19'b0010001000100100001: color_data = Z;
		19'b0010001000100100010: color_data = Z;
		19'b0010001000100100011: color_data = Z;
		19'b0010001000100100100: color_data = Z;
		19'b0010001000100100101: color_data = Z;
		19'b0010001000100100110: color_data = Z;
		19'b0010001000100100111: color_data = Z;
		19'b0010001000100101000: color_data = Z;
		19'b0010001000100101001: color_data = Z;
		19'b0010001000100101010: color_data = Z;
		19'b0010001000100101011: color_data = Z;
		19'b0010001000100101100: color_data = Z;
		19'b0010001000100101101: color_data = Z;
		19'b0010001000100101110: color_data = Z;
		19'b0010001000100101111: color_data = Z;
		19'b0010001000100110000: color_data = Z;
		19'b0010001000100110001: color_data = Z;
		19'b0010001000100110010: color_data = Z;
		19'b0010001000100110011: color_data = Z;
		19'b0010001000100110100: color_data = Z;
		19'b0010001000100110101: color_data = Z;
		19'b0010001000100110110: color_data = Z;
		19'b0010001000100110111: color_data = Z;
		19'b0010001000100111000: color_data = Z;
		19'b0010001000100111001: color_data = Z;
		19'b0010001000100111010: color_data = Z;
		19'b0010001000100111011: color_data = Z;
		19'b0010001000100111100: color_data = Z;
		19'b0010001000100111101: color_data = Z;
		19'b0010001000100111110: color_data = Z;
		19'b0010001000100111111: color_data = Z;
		19'b0010001000101000000: color_data = Z;
		19'b0010001000101000001: color_data = Z;
		19'b0010001000101000010: color_data = Z;
		19'b0010001000101000011: color_data = Z;
		19'b0010001000101000100: color_data = Z;
		19'b0010001000101000101: color_data = Z;
		19'b0010001000101000110: color_data = Z;
		19'b0010001000101000111: color_data = Z;
		19'b0010001000101001000: color_data = Z;
		19'b0010001000101001001: color_data = Z;
		19'b0010001000101001010: color_data = Z;
		19'b0010001000101001011: color_data = Z;
		19'b0010001000101001100: color_data = Z;
		19'b0010001000101001101: color_data = Z;
		19'b0010001000101001110: color_data = Z;
		19'b0010001000101001111: color_data = Z;
		19'b0010001000101010000: color_data = Z;
		19'b0010001000101010001: color_data = Z;
		19'b0010001000101010010: color_data = Z;
		19'b0010001000101010011: color_data = Z;
		19'b0010001000101010100: color_data = Z;
		19'b0010001000101010101: color_data = Z;
		19'b0010001000101010110: color_data = Z;
		19'b0010001000101010111: color_data = Z;
		19'b0010001000101011000: color_data = Z;
		19'b0010001000101011001: color_data = Z;
		19'b0010001000101011010: color_data = Z;
		19'b0010001000101011011: color_data = Z;
		19'b0010001000101011100: color_data = Z;
		19'b0010001000101011101: color_data = Z;
		19'b0010001000101011110: color_data = Z;
		19'b0010001000101011111: color_data = Z;
		19'b0010001000101100000: color_data = Z;
		19'b0010001000101100001: color_data = Z;
		19'b0010001000101100010: color_data = Z;
		19'b0010001000101100011: color_data = Z;
		19'b0010001000101100100: color_data = Z;
		19'b0010001000101100101: color_data = Z;
		19'b0010001000101100110: color_data = Z;
		19'b0010001000101100111: color_data = Z;
		19'b0010001000101101000: color_data = Z;
		19'b0010001000101101001: color_data = Z;
		19'b0010001000101101010: color_data = Z;
		19'b0010001000101101011: color_data = Z;
		19'b0010001000101101100: color_data = Z;
		19'b0010001000101101101: color_data = Z;
		19'b0010001000101101110: color_data = Z;
		19'b0010001000101101111: color_data = Z;
		19'b0010001000101110000: color_data = Z;
		19'b0010001000101110001: color_data = Z;
		19'b0010001000101110010: color_data = Z;
		19'b0010001000101110011: color_data = Z;
		19'b0010001000101110100: color_data = Z;
		19'b0010001000101110101: color_data = Z;
		19'b0010001000101110110: color_data = Z;
		19'b0010001000101110111: color_data = Z;
		19'b0010001000101111000: color_data = Z;
		19'b0010001000101111001: color_data = Z;
		19'b0010001000101111010: color_data = Z;
		19'b0010001000101111011: color_data = Z;
		19'b0010001000101111100: color_data = Z;
		19'b0010001000101111101: color_data = Z;
		19'b0010001000101111110: color_data = Z;
		19'b0010001000101111111: color_data = Z;
		19'b0010001000110000000: color_data = Z;
		19'b0010001000110000001: color_data = Z;
		19'b0010001000110000010: color_data = Z;
		19'b0010001000110000011: color_data = Z;
		19'b0010001000110000100: color_data = Z;
		19'b0010001000110000101: color_data = Z;
		19'b0010001000110000110: color_data = Z;
		19'b0010001000110000111: color_data = Z;
		19'b0010001000110001000: color_data = Z;
		19'b0010001000110001001: color_data = Z;
		19'b0010001000110001010: color_data = Z;
		19'b0010001000110001011: color_data = Z;
		19'b0010001000110001100: color_data = Z;
		19'b0010001000110001101: color_data = Z;
		19'b0010001000110001110: color_data = Z;
		19'b0010001000110001111: color_data = Z;
		19'b0010001000110010000: color_data = Z;
		19'b0010001000110010001: color_data = Z;
		19'b0010001000110010010: color_data = Z;
		19'b0010001000110010011: color_data = Z;
		19'b0010001000110010100: color_data = Z;
		19'b0010001000110010101: color_data = Z;
		19'b0010001000110010110: color_data = Z;
		19'b0010001000110010111: color_data = Z;
		19'b0010001000110011000: color_data = Z;
		19'b0010001000110011001: color_data = Z;
		19'b0010001000110011010: color_data = Z;
		19'b0010001000110011011: color_data = Z;
		19'b0010001000110011100: color_data = Z;
		19'b0010001000110011101: color_data = Z;
		19'b0010001000110011110: color_data = Z;
		19'b0010001000110011111: color_data = Z;
		19'b0010001000110100000: color_data = Z;
		19'b0010001000110100001: color_data = Z;
		19'b0010001000110100010: color_data = Z;
		19'b0010001000110100011: color_data = Z;
		19'b0010001000110100100: color_data = Z;
		19'b0010001000110100101: color_data = Z;
		19'b0010001000110100110: color_data = Z;
		19'b0010001000110100111: color_data = Z;
		19'b0010001000110101000: color_data = Z;
		19'b0010001000110101001: color_data = Z;
		19'b0010001000110101110: color_data = Z;
		19'b0010001000110101111: color_data = Z;
		19'b0010001000110110000: color_data = Z;
		19'b0010001000110110001: color_data = Z;
		19'b0010001000110110010: color_data = Z;
		19'b0010001000110110011: color_data = Z;
		19'b0010001000110111000: color_data = Z;
		19'b0010001000110111001: color_data = Z;
		19'b0010001000110111010: color_data = Z;
		19'b0010001000110111011: color_data = Z;
		19'b0010001000110111100: color_data = Z;
		19'b0010001000110111101: color_data = Z;
		19'b0010001000110111110: color_data = Z;
		19'b0010001000110111111: color_data = Z;
		19'b0010001000111000000: color_data = Z;
		19'b0010001000111000001: color_data = Z;
		19'b0010001000111000010: color_data = Z;
		19'b0010001000111000011: color_data = Z;
		19'b0010001000111000100: color_data = Z;
		19'b0010001010011001101: color_data = Z;
		19'b0010001010011001110: color_data = Z;
		19'b0010001010011001111: color_data = Z;
		19'b0010001010011010000: color_data = Z;
		19'b0010001010011010001: color_data = Z;
		19'b0010001010011010010: color_data = Z;
		19'b0010001010011010011: color_data = Z;
		19'b0010001010011010100: color_data = Z;
		19'b0010001010011010101: color_data = Z;
		19'b0010001010011010110: color_data = Z;
		19'b0010001010011010111: color_data = Z;
		19'b0010001010011011000: color_data = Z;
		19'b0010001010011011001: color_data = Z;
		19'b0010001010011011010: color_data = Z;
		19'b0010001010011011011: color_data = Z;
		19'b0010001010011011100: color_data = Z;
		19'b0010001010011011101: color_data = Z;
		19'b0010001010011011110: color_data = Z;
		19'b0010001010011011111: color_data = Z;
		19'b0010001010011100000: color_data = Z;
		19'b0010001010011100001: color_data = Z;
		19'b0010001010011100010: color_data = Z;
		19'b0010001010011100011: color_data = Z;
		19'b0010001010011100100: color_data = Z;
		19'b0010001010011100101: color_data = Z;
		19'b0010001010011100110: color_data = Z;
		19'b0010001010011100111: color_data = Z;
		19'b0010001010011101000: color_data = Z;
		19'b0010001010011101001: color_data = Z;
		19'b0010001010011101010: color_data = Z;
		19'b0010001010011101011: color_data = Z;
		19'b0010001010011101100: color_data = Z;
		19'b0010001010011101101: color_data = Z;
		19'b0010001010011101110: color_data = Z;
		19'b0010001010011101111: color_data = Z;
		19'b0010001010011110000: color_data = Z;
		19'b0010001010011110001: color_data = Z;
		19'b0010001010011110010: color_data = Z;
		19'b0010001010011110011: color_data = Z;
		19'b0010001010011110100: color_data = Z;
		19'b0010001010011110101: color_data = Z;
		19'b0010001010011110110: color_data = Z;
		19'b0010001010011110111: color_data = Z;
		19'b0010001010011111000: color_data = Z;
		19'b0010001010011111001: color_data = Z;
		19'b0010001010011111010: color_data = Z;
		19'b0010001010011111011: color_data = Z;
		19'b0010001010011111100: color_data = Z;
		19'b0010001010011111101: color_data = Z;
		19'b0010001010011111110: color_data = Z;
		19'b0010001010011111111: color_data = Z;
		19'b0010001010100000000: color_data = Z;
		19'b0010001010100000001: color_data = Z;
		19'b0010001010100000010: color_data = Z;
		19'b0010001010100000011: color_data = Z;
		19'b0010001010100000100: color_data = Z;
		19'b0010001010100000101: color_data = Z;
		19'b0010001010100000110: color_data = Z;
		19'b0010001010100000111: color_data = Z;
		19'b0010001010100001000: color_data = Z;
		19'b0010001010100001001: color_data = Z;
		19'b0010001010100001010: color_data = Z;
		19'b0010001010100001011: color_data = Z;
		19'b0010001010100001100: color_data = Z;
		19'b0010001010100001101: color_data = Z;
		19'b0010001010100001110: color_data = Z;
		19'b0010001010100001111: color_data = Z;
		19'b0010001010100010000: color_data = Z;
		19'b0010001010100010001: color_data = Z;
		19'b0010001010100010010: color_data = Z;
		19'b0010001010100010011: color_data = Z;
		19'b0010001010100010100: color_data = Z;
		19'b0010001010100010101: color_data = Z;
		19'b0010001010100010110: color_data = Z;
		19'b0010001010100010111: color_data = Z;
		19'b0010001010100011000: color_data = Z;
		19'b0010001010100011001: color_data = Z;
		19'b0010001010100011010: color_data = Z;
		19'b0010001010100011011: color_data = Z;
		19'b0010001010100011100: color_data = Z;
		19'b0010001010100011101: color_data = Z;
		19'b0010001010100011110: color_data = Z;
		19'b0010001010100011111: color_data = Z;
		19'b0010001010100100000: color_data = Z;
		19'b0010001010100100001: color_data = Z;
		19'b0010001010100100010: color_data = Z;
		19'b0010001010100100011: color_data = Z;
		19'b0010001010100100100: color_data = Z;
		19'b0010001010100100101: color_data = Z;
		19'b0010001010100100110: color_data = Z;
		19'b0010001010100100111: color_data = Z;
		19'b0010001010100101000: color_data = Z;
		19'b0010001010100101001: color_data = Z;
		19'b0010001010100101010: color_data = Z;
		19'b0010001010100101011: color_data = Z;
		19'b0010001010100101100: color_data = Z;
		19'b0010001010100101101: color_data = Z;
		19'b0010001010100101110: color_data = Z;
		19'b0010001010100101111: color_data = Z;
		19'b0010001010100110000: color_data = Z;
		19'b0010001010100110001: color_data = Z;
		19'b0010001010100110010: color_data = Z;
		19'b0010001010100110011: color_data = Z;
		19'b0010001010100110100: color_data = Z;
		19'b0010001010100110101: color_data = Z;
		19'b0010001010100110110: color_data = Z;
		19'b0010001010100110111: color_data = Z;
		19'b0010001010100111000: color_data = Z;
		19'b0010001010100111001: color_data = Z;
		19'b0010001010100111010: color_data = Z;
		19'b0010001010100111011: color_data = Z;
		19'b0010001010100111100: color_data = Z;
		19'b0010001010100111101: color_data = Z;
		19'b0010001010100111110: color_data = Z;
		19'b0010001010100111111: color_data = Z;
		19'b0010001010101000000: color_data = Z;
		19'b0010001010101000001: color_data = Z;
		19'b0010001010101000010: color_data = Z;
		19'b0010001010101000011: color_data = Z;
		19'b0010001010101000100: color_data = Z;
		19'b0010001010101000101: color_data = Z;
		19'b0010001010101000110: color_data = Z;
		19'b0010001010101000111: color_data = Z;
		19'b0010001010101001000: color_data = Z;
		19'b0010001010101001001: color_data = Z;
		19'b0010001010101001010: color_data = Z;
		19'b0010001010101001011: color_data = Z;
		19'b0010001010101001100: color_data = Z;
		19'b0010001010101001101: color_data = Z;
		19'b0010001010101001110: color_data = Z;
		19'b0010001010101001111: color_data = Z;
		19'b0010001010101010000: color_data = Z;
		19'b0010001010101010001: color_data = Z;
		19'b0010001010101010010: color_data = Z;
		19'b0010001010101010011: color_data = Z;
		19'b0010001010101010100: color_data = Z;
		19'b0010001010101010101: color_data = Z;
		19'b0010001010101010110: color_data = Z;
		19'b0010001010101010111: color_data = Z;
		19'b0010001010101011000: color_data = Z;
		19'b0010001010101011001: color_data = Z;
		19'b0010001010101011010: color_data = Z;
		19'b0010001010101011011: color_data = Z;
		19'b0010001010101011100: color_data = Z;
		19'b0010001010101011101: color_data = Z;
		19'b0010001010101011110: color_data = Z;
		19'b0010001010101011111: color_data = Z;
		19'b0010001010101100000: color_data = Z;
		19'b0010001010101100001: color_data = Z;
		19'b0010001010101100010: color_data = Z;
		19'b0010001010101100011: color_data = Z;
		19'b0010001010101100100: color_data = Z;
		19'b0010001010101100101: color_data = Z;
		19'b0010001010101100110: color_data = Z;
		19'b0010001010101100111: color_data = Z;
		19'b0010001010101101000: color_data = Z;
		19'b0010001010101101001: color_data = Z;
		19'b0010001010101101010: color_data = Z;
		19'b0010001010101101011: color_data = Z;
		19'b0010001010101101100: color_data = Z;
		19'b0010001010101101101: color_data = Z;
		19'b0010001010101101110: color_data = Z;
		19'b0010001010101101111: color_data = Z;
		19'b0010001010101110000: color_data = Z;
		19'b0010001010101110001: color_data = Z;
		19'b0010001010101110010: color_data = Z;
		19'b0010001010101110011: color_data = Z;
		19'b0010001010101110100: color_data = Z;
		19'b0010001010101110101: color_data = Z;
		19'b0010001010101110110: color_data = Z;
		19'b0010001010101110111: color_data = Z;
		19'b0010001010101111000: color_data = Z;
		19'b0010001010101111001: color_data = Z;
		19'b0010001010101111010: color_data = Z;
		19'b0010001010101111011: color_data = Z;
		19'b0010001010101111100: color_data = Z;
		19'b0010001010101111101: color_data = Z;
		19'b0010001010101111110: color_data = Z;
		19'b0010001010101111111: color_data = Z;
		19'b0010001010110000000: color_data = Z;
		19'b0010001010110000001: color_data = Z;
		19'b0010001010110000010: color_data = Z;
		19'b0010001010110000011: color_data = Z;
		19'b0010001010110000100: color_data = Z;
		19'b0010001010110000101: color_data = Z;
		19'b0010001010110000110: color_data = Z;
		19'b0010001010110000111: color_data = Z;
		19'b0010001010110001000: color_data = Z;
		19'b0010001010110001001: color_data = Z;
		19'b0010001010110001010: color_data = Z;
		19'b0010001010110001011: color_data = Z;
		19'b0010001010110001100: color_data = Z;
		19'b0010001010110001101: color_data = Z;
		19'b0010001010110001110: color_data = Z;
		19'b0010001010110001111: color_data = Z;
		19'b0010001010110010000: color_data = Z;
		19'b0010001010110010001: color_data = Z;
		19'b0010001010110010010: color_data = Z;
		19'b0010001010110010011: color_data = Z;
		19'b0010001010110010100: color_data = Z;
		19'b0010001010110010101: color_data = Z;
		19'b0010001010110010110: color_data = Z;
		19'b0010001010110010111: color_data = Z;
		19'b0010001010110011000: color_data = Z;
		19'b0010001010110011001: color_data = Z;
		19'b0010001010110011010: color_data = Z;
		19'b0010001010110011011: color_data = Z;
		19'b0010001010110011100: color_data = Z;
		19'b0010001010110011101: color_data = Z;
		19'b0010001010110011110: color_data = Z;
		19'b0010001010110011111: color_data = Z;
		19'b0010001010110100000: color_data = Z;
		19'b0010001010110100001: color_data = Z;
		19'b0010001010110100010: color_data = Z;
		19'b0010001010110100011: color_data = Z;
		19'b0010001010110100100: color_data = Z;
		19'b0010001010110100101: color_data = Z;
		19'b0010001010110100110: color_data = Z;
		19'b0010001010110100111: color_data = Z;
		19'b0010001010110101000: color_data = Z;
		19'b0010001010110101001: color_data = Z;
		19'b0010001010110101010: color_data = Z;
		19'b0010001010110101111: color_data = Z;
		19'b0010001010110110000: color_data = Z;
		19'b0010001010110110001: color_data = Z;
		19'b0010001010110110010: color_data = Z;
		19'b0010001010110110011: color_data = Z;
		19'b0010001010110111000: color_data = Z;
		19'b0010001010110111001: color_data = Z;
		19'b0010001010110111010: color_data = Z;
		19'b0010001010110111011: color_data = Z;
		19'b0010001010110111100: color_data = Z;
		19'b0010001010110111101: color_data = Z;
		19'b0010001010110111110: color_data = Z;
		19'b0010001010110111111: color_data = Z;
		19'b0010001010111000000: color_data = Z;
		19'b0010001010111000001: color_data = Z;
		19'b0010001010111000010: color_data = Z;
		19'b0010001010111000011: color_data = Z;
		19'b0010001010111000100: color_data = Z;
		19'b0010001010111000101: color_data = Z;
		19'b0010001100011001101: color_data = Z;
		19'b0010001100011001110: color_data = Z;
		19'b0010001100011001111: color_data = Z;
		19'b0010001100011010000: color_data = Z;
		19'b0010001100011010001: color_data = Z;
		19'b0010001100011010010: color_data = Z;
		19'b0010001100011010011: color_data = Z;
		19'b0010001100011010100: color_data = Z;
		19'b0010001100011010101: color_data = Z;
		19'b0010001100011010110: color_data = Z;
		19'b0010001100011010111: color_data = Z;
		19'b0010001100011011000: color_data = Z;
		19'b0010001100011011001: color_data = Z;
		19'b0010001100011011010: color_data = Z;
		19'b0010001100011011011: color_data = Z;
		19'b0010001100011011100: color_data = Z;
		19'b0010001100011011101: color_data = Z;
		19'b0010001100011011110: color_data = Z;
		19'b0010001100011011111: color_data = Z;
		19'b0010001100011100000: color_data = Z;
		19'b0010001100011100001: color_data = Z;
		19'b0010001100011100010: color_data = Z;
		19'b0010001100011100011: color_data = Z;
		19'b0010001100011100100: color_data = Z;
		19'b0010001100011100101: color_data = Z;
		19'b0010001100011100110: color_data = Z;
		19'b0010001100011100111: color_data = Z;
		19'b0010001100011101000: color_data = Z;
		19'b0010001100011101001: color_data = Z;
		19'b0010001100011101010: color_data = Z;
		19'b0010001100011101011: color_data = Z;
		19'b0010001100011101100: color_data = Z;
		19'b0010001100011101101: color_data = Z;
		19'b0010001100011101110: color_data = Z;
		19'b0010001100011101111: color_data = Z;
		19'b0010001100011110000: color_data = Z;
		19'b0010001100011110001: color_data = Z;
		19'b0010001100011110010: color_data = Z;
		19'b0010001100011110011: color_data = Z;
		19'b0010001100011110100: color_data = Z;
		19'b0010001100011110101: color_data = Z;
		19'b0010001100011110110: color_data = Z;
		19'b0010001100011110111: color_data = Z;
		19'b0010001100011111000: color_data = Z;
		19'b0010001100011111001: color_data = Z;
		19'b0010001100011111010: color_data = Z;
		19'b0010001100011111011: color_data = Z;
		19'b0010001100011111100: color_data = Z;
		19'b0010001100011111101: color_data = Z;
		19'b0010001100011111110: color_data = Z;
		19'b0010001100011111111: color_data = Z;
		19'b0010001100100000000: color_data = Z;
		19'b0010001100100000001: color_data = Z;
		19'b0010001100100000010: color_data = Z;
		19'b0010001100100000011: color_data = Z;
		19'b0010001100100000100: color_data = Z;
		19'b0010001100100000101: color_data = Z;
		19'b0010001100100000110: color_data = Z;
		19'b0010001100100000111: color_data = Z;
		19'b0010001100100001000: color_data = Z;
		19'b0010001100100001001: color_data = Z;
		19'b0010001100100001010: color_data = Z;
		19'b0010001100100001011: color_data = Z;
		19'b0010001100100001100: color_data = Z;
		19'b0010001100100001101: color_data = Z;
		19'b0010001100100001110: color_data = Z;
		19'b0010001100100001111: color_data = Z;
		19'b0010001100100010000: color_data = Z;
		19'b0010001100100010001: color_data = Z;
		19'b0010001100100010010: color_data = Z;
		19'b0010001100100010011: color_data = Z;
		19'b0010001100100010100: color_data = Z;
		19'b0010001100100010101: color_data = Z;
		19'b0010001100100010110: color_data = Z;
		19'b0010001100100010111: color_data = Z;
		19'b0010001100100011000: color_data = Z;
		19'b0010001100100011001: color_data = Z;
		19'b0010001100100011010: color_data = Z;
		19'b0010001100100011011: color_data = Z;
		19'b0010001100100011100: color_data = Z;
		19'b0010001100100011101: color_data = Z;
		19'b0010001100100011110: color_data = Z;
		19'b0010001100100011111: color_data = Z;
		19'b0010001100100100000: color_data = Z;
		19'b0010001100100100001: color_data = Z;
		19'b0010001100100100010: color_data = Z;
		19'b0010001100100100011: color_data = Z;
		19'b0010001100100100100: color_data = Z;
		19'b0010001100100100101: color_data = Z;
		19'b0010001100100100110: color_data = Z;
		19'b0010001100100100111: color_data = Z;
		19'b0010001100100101000: color_data = Z;
		19'b0010001100100101001: color_data = Z;
		19'b0010001100100101010: color_data = Z;
		19'b0010001100100101011: color_data = Z;
		19'b0010001100100101100: color_data = Z;
		19'b0010001100100101101: color_data = Z;
		19'b0010001100100101110: color_data = Z;
		19'b0010001100100101111: color_data = Z;
		19'b0010001100100110000: color_data = Z;
		19'b0010001100100110001: color_data = Z;
		19'b0010001100100110010: color_data = Z;
		19'b0010001100100110011: color_data = Z;
		19'b0010001100100110100: color_data = Z;
		19'b0010001100100110101: color_data = Z;
		19'b0010001100100110110: color_data = Z;
		19'b0010001100100110111: color_data = Z;
		19'b0010001100100111000: color_data = Z;
		19'b0010001100100111001: color_data = Z;
		19'b0010001100100111010: color_data = Z;
		19'b0010001100100111011: color_data = Z;
		19'b0010001100100111100: color_data = Z;
		19'b0010001100100111101: color_data = Z;
		19'b0010001100100111110: color_data = Z;
		19'b0010001100100111111: color_data = Z;
		19'b0010001100101000000: color_data = Z;
		19'b0010001100101000001: color_data = Z;
		19'b0010001100101000010: color_data = Z;
		19'b0010001100101000011: color_data = Z;
		19'b0010001100101000100: color_data = Z;
		19'b0010001100101000101: color_data = Z;
		19'b0010001100101000110: color_data = Z;
		19'b0010001100101000111: color_data = Z;
		19'b0010001100101001000: color_data = Z;
		19'b0010001100101001001: color_data = Z;
		19'b0010001100101001010: color_data = Z;
		19'b0010001100101001011: color_data = Z;
		19'b0010001100101001100: color_data = Z;
		19'b0010001100101001101: color_data = Z;
		19'b0010001100101001110: color_data = Z;
		19'b0010001100101001111: color_data = Z;
		19'b0010001100101010000: color_data = Z;
		19'b0010001100101010001: color_data = Z;
		19'b0010001100101010010: color_data = Z;
		19'b0010001100101010011: color_data = Z;
		19'b0010001100101010100: color_data = Z;
		19'b0010001100101010101: color_data = Z;
		19'b0010001100101010110: color_data = Z;
		19'b0010001100101010111: color_data = Z;
		19'b0010001100101011000: color_data = Z;
		19'b0010001100101011001: color_data = Z;
		19'b0010001100101011010: color_data = Z;
		19'b0010001100101011011: color_data = Z;
		19'b0010001100101011100: color_data = Z;
		19'b0010001100101011101: color_data = Z;
		19'b0010001100101011110: color_data = Z;
		19'b0010001100101011111: color_data = Z;
		19'b0010001100101100000: color_data = Z;
		19'b0010001100101100001: color_data = Z;
		19'b0010001100101100010: color_data = Z;
		19'b0010001100101100011: color_data = Z;
		19'b0010001100101100100: color_data = Z;
		19'b0010001100101100101: color_data = Z;
		19'b0010001100101100110: color_data = Z;
		19'b0010001100101100111: color_data = Z;
		19'b0010001100101101000: color_data = Z;
		19'b0010001100101101001: color_data = Z;
		19'b0010001100101101010: color_data = Z;
		19'b0010001100101101011: color_data = Z;
		19'b0010001100101101100: color_data = Z;
		19'b0010001100101101101: color_data = Z;
		19'b0010001100101101110: color_data = Z;
		19'b0010001100101101111: color_data = Z;
		19'b0010001100101110000: color_data = Z;
		19'b0010001100101110001: color_data = Z;
		19'b0010001100101110010: color_data = Z;
		19'b0010001100101110011: color_data = Z;
		19'b0010001100101110100: color_data = Z;
		19'b0010001100101110101: color_data = Z;
		19'b0010001100101110110: color_data = Z;
		19'b0010001100101110111: color_data = Z;
		19'b0010001100101111000: color_data = Z;
		19'b0010001100101111001: color_data = Z;
		19'b0010001100101111010: color_data = Z;
		19'b0010001100101111011: color_data = Z;
		19'b0010001100101111100: color_data = Z;
		19'b0010001100101111101: color_data = Z;
		19'b0010001100101111110: color_data = Z;
		19'b0010001100101111111: color_data = Z;
		19'b0010001100110000000: color_data = Z;
		19'b0010001100110000001: color_data = Z;
		19'b0010001100110000010: color_data = Z;
		19'b0010001100110000011: color_data = Z;
		19'b0010001100110000100: color_data = Z;
		19'b0010001100110000101: color_data = Z;
		19'b0010001100110000110: color_data = Z;
		19'b0010001100110000111: color_data = Z;
		19'b0010001100110001000: color_data = Z;
		19'b0010001100110001001: color_data = Z;
		19'b0010001100110001010: color_data = Z;
		19'b0010001100110001011: color_data = Z;
		19'b0010001100110001100: color_data = Z;
		19'b0010001100110001101: color_data = Z;
		19'b0010001100110001110: color_data = Z;
		19'b0010001100110001111: color_data = Z;
		19'b0010001100110010000: color_data = Z;
		19'b0010001100110010001: color_data = Z;
		19'b0010001100110010010: color_data = Z;
		19'b0010001100110010011: color_data = Z;
		19'b0010001100110010100: color_data = Z;
		19'b0010001100110010101: color_data = Z;
		19'b0010001100110010110: color_data = Z;
		19'b0010001100110010111: color_data = Z;
		19'b0010001100110011000: color_data = Z;
		19'b0010001100110011001: color_data = Z;
		19'b0010001100110011010: color_data = Z;
		19'b0010001100110011011: color_data = Z;
		19'b0010001100110011100: color_data = Z;
		19'b0010001100110011101: color_data = Z;
		19'b0010001100110011110: color_data = Z;
		19'b0010001100110011111: color_data = Z;
		19'b0010001100110100000: color_data = Z;
		19'b0010001100110100001: color_data = Z;
		19'b0010001100110100010: color_data = Z;
		19'b0010001100110100011: color_data = Z;
		19'b0010001100110100100: color_data = Z;
		19'b0010001100110100101: color_data = Z;
		19'b0010001100110100110: color_data = Z;
		19'b0010001100110100111: color_data = Z;
		19'b0010001100110101000: color_data = Z;
		19'b0010001100110101001: color_data = Z;
		19'b0010001100110101010: color_data = Z;
		19'b0010001100110101111: color_data = Z;
		19'b0010001100110110000: color_data = Z;
		19'b0010001100110110001: color_data = Z;
		19'b0010001100110110010: color_data = Z;
		19'b0010001100110110011: color_data = Z;
		19'b0010001100110111001: color_data = Z;
		19'b0010001100110111010: color_data = Z;
		19'b0010001100110111011: color_data = Z;
		19'b0010001100110111100: color_data = Z;
		19'b0010001100110111101: color_data = Z;
		19'b0010001100110111110: color_data = Z;
		19'b0010001100110111111: color_data = Z;
		19'b0010001100111000000: color_data = Z;
		19'b0010001100111000001: color_data = Z;
		19'b0010001100111000010: color_data = Z;
		19'b0010001100111000011: color_data = Z;
		19'b0010001100111000100: color_data = Z;
		19'b0010001100111000101: color_data = Z;
		19'b0010001100111000110: color_data = Z;
		19'b0010001110011001100: color_data = Z;
		19'b0010001110011001101: color_data = Z;
		19'b0010001110011001110: color_data = Z;
		19'b0010001110011001111: color_data = Z;
		19'b0010001110011010000: color_data = Z;
		19'b0010001110011010001: color_data = Z;
		19'b0010001110011010010: color_data = Z;
		19'b0010001110011010011: color_data = Z;
		19'b0010001110011010100: color_data = Z;
		19'b0010001110011010101: color_data = Z;
		19'b0010001110011010110: color_data = Z;
		19'b0010001110011010111: color_data = Z;
		19'b0010001110011011000: color_data = Z;
		19'b0010001110011011001: color_data = Z;
		19'b0010001110011011010: color_data = Z;
		19'b0010001110011011011: color_data = Z;
		19'b0010001110011011100: color_data = Z;
		19'b0010001110011011101: color_data = Z;
		19'b0010001110011011110: color_data = Z;
		19'b0010001110011011111: color_data = Z;
		19'b0010001110011100000: color_data = Z;
		19'b0010001110011100001: color_data = Z;
		19'b0010001110011100010: color_data = Z;
		19'b0010001110011100011: color_data = Z;
		19'b0010001110011100100: color_data = Z;
		19'b0010001110011100101: color_data = Z;
		19'b0010001110011100110: color_data = Z;
		19'b0010001110011100111: color_data = Z;
		19'b0010001110011101000: color_data = Z;
		19'b0010001110011101001: color_data = Z;
		19'b0010001110011101010: color_data = Z;
		19'b0010001110011101011: color_data = Z;
		19'b0010001110011101100: color_data = Z;
		19'b0010001110011101101: color_data = Z;
		19'b0010001110011101110: color_data = Z;
		19'b0010001110011101111: color_data = Z;
		19'b0010001110011110000: color_data = Z;
		19'b0010001110011110001: color_data = Z;
		19'b0010001110011110010: color_data = Z;
		19'b0010001110011110011: color_data = Z;
		19'b0010001110011110100: color_data = Z;
		19'b0010001110011110101: color_data = Z;
		19'b0010001110011110110: color_data = Z;
		19'b0010001110011110111: color_data = Z;
		19'b0010001110011111000: color_data = Z;
		19'b0010001110011111001: color_data = Z;
		19'b0010001110011111010: color_data = Z;
		19'b0010001110011111011: color_data = Z;
		19'b0010001110011111100: color_data = Z;
		19'b0010001110011111101: color_data = Z;
		19'b0010001110011111110: color_data = Z;
		19'b0010001110011111111: color_data = Z;
		19'b0010001110100000000: color_data = Z;
		19'b0010001110100000001: color_data = Z;
		19'b0010001110100000010: color_data = Z;
		19'b0010001110100000011: color_data = Z;
		19'b0010001110100000100: color_data = Z;
		19'b0010001110100000101: color_data = Z;
		19'b0010001110100000110: color_data = Z;
		19'b0010001110100000111: color_data = Z;
		19'b0010001110100001000: color_data = Z;
		19'b0010001110100001001: color_data = Z;
		19'b0010001110100001010: color_data = Z;
		19'b0010001110100001011: color_data = Z;
		19'b0010001110100001100: color_data = Z;
		19'b0010001110100001101: color_data = Z;
		19'b0010001110100001110: color_data = Z;
		19'b0010001110100001111: color_data = Z;
		19'b0010001110100010000: color_data = Z;
		19'b0010001110100010001: color_data = Z;
		19'b0010001110100010010: color_data = Z;
		19'b0010001110100010011: color_data = Z;
		19'b0010001110100010100: color_data = Z;
		19'b0010001110100010101: color_data = Z;
		19'b0010001110100010110: color_data = Z;
		19'b0010001110100010111: color_data = Z;
		19'b0010001110100011000: color_data = Z;
		19'b0010001110100011001: color_data = Z;
		19'b0010001110100011010: color_data = Z;
		19'b0010001110100011011: color_data = Z;
		19'b0010001110100011100: color_data = Z;
		19'b0010001110100011101: color_data = Z;
		19'b0010001110100011110: color_data = Z;
		19'b0010001110100011111: color_data = Z;
		19'b0010001110100100000: color_data = Z;
		19'b0010001110100100001: color_data = Z;
		19'b0010001110100100010: color_data = Z;
		19'b0010001110100100011: color_data = Z;
		19'b0010001110100100100: color_data = Z;
		19'b0010001110100100101: color_data = Z;
		19'b0010001110100100110: color_data = Z;
		19'b0010001110100100111: color_data = Z;
		19'b0010001110100101000: color_data = Z;
		19'b0010001110100101001: color_data = Z;
		19'b0010001110100101010: color_data = Z;
		19'b0010001110100101011: color_data = Z;
		19'b0010001110100101100: color_data = Z;
		19'b0010001110100101101: color_data = Z;
		19'b0010001110100101110: color_data = Z;
		19'b0010001110100101111: color_data = Z;
		19'b0010001110100110000: color_data = Z;
		19'b0010001110100110001: color_data = Z;
		19'b0010001110100110010: color_data = Z;
		19'b0010001110100110011: color_data = Z;
		19'b0010001110100110100: color_data = Z;
		19'b0010001110100110101: color_data = Z;
		19'b0010001110100110110: color_data = Z;
		19'b0010001110100110111: color_data = Z;
		19'b0010001110100111000: color_data = Z;
		19'b0010001110100111001: color_data = Z;
		19'b0010001110100111010: color_data = Z;
		19'b0010001110100111011: color_data = Z;
		19'b0010001110100111100: color_data = Z;
		19'b0010001110100111101: color_data = Z;
		19'b0010001110100111110: color_data = Z;
		19'b0010001110100111111: color_data = Z;
		19'b0010001110101000000: color_data = Z;
		19'b0010001110101000001: color_data = Z;
		19'b0010001110101000010: color_data = Z;
		19'b0010001110101000011: color_data = Z;
		19'b0010001110101000100: color_data = Z;
		19'b0010001110101000101: color_data = Z;
		19'b0010001110101000110: color_data = Z;
		19'b0010001110101000111: color_data = Z;
		19'b0010001110101001000: color_data = Z;
		19'b0010001110101001001: color_data = Z;
		19'b0010001110101001010: color_data = Z;
		19'b0010001110101001011: color_data = Z;
		19'b0010001110101001100: color_data = Z;
		19'b0010001110101001101: color_data = Z;
		19'b0010001110101001110: color_data = Z;
		19'b0010001110101001111: color_data = Z;
		19'b0010001110101010000: color_data = Z;
		19'b0010001110101010001: color_data = Z;
		19'b0010001110101010010: color_data = Z;
		19'b0010001110101010011: color_data = Z;
		19'b0010001110101010100: color_data = Z;
		19'b0010001110101010101: color_data = Z;
		19'b0010001110101010110: color_data = Z;
		19'b0010001110101010111: color_data = Z;
		19'b0010001110101011000: color_data = Z;
		19'b0010001110101011001: color_data = Z;
		19'b0010001110101011010: color_data = Z;
		19'b0010001110101011011: color_data = Z;
		19'b0010001110101011100: color_data = Z;
		19'b0010001110101011101: color_data = Z;
		19'b0010001110101011110: color_data = Z;
		19'b0010001110101011111: color_data = Z;
		19'b0010001110101100000: color_data = Z;
		19'b0010001110101100001: color_data = Z;
		19'b0010001110101100010: color_data = Z;
		19'b0010001110101100011: color_data = Z;
		19'b0010001110101100100: color_data = Z;
		19'b0010001110101100101: color_data = Z;
		19'b0010001110101100110: color_data = Z;
		19'b0010001110101100111: color_data = Z;
		19'b0010001110101101000: color_data = Z;
		19'b0010001110101101001: color_data = Z;
		19'b0010001110101101010: color_data = Z;
		19'b0010001110101101011: color_data = Z;
		19'b0010001110101101100: color_data = Z;
		19'b0010001110101101101: color_data = Z;
		19'b0010001110101101110: color_data = Z;
		19'b0010001110101101111: color_data = Z;
		19'b0010001110101110000: color_data = Z;
		19'b0010001110101110001: color_data = Z;
		19'b0010001110101110010: color_data = Z;
		19'b0010001110101110011: color_data = Z;
		19'b0010001110101110100: color_data = Z;
		19'b0010001110101110101: color_data = Z;
		19'b0010001110101110110: color_data = Z;
		19'b0010001110101110111: color_data = Z;
		19'b0010001110101111000: color_data = Z;
		19'b0010001110101111001: color_data = Z;
		19'b0010001110101111010: color_data = Z;
		19'b0010001110101111011: color_data = Z;
		19'b0010001110101111100: color_data = Z;
		19'b0010001110101111101: color_data = Z;
		19'b0010001110101111110: color_data = Z;
		19'b0010001110101111111: color_data = Z;
		19'b0010001110110000000: color_data = Z;
		19'b0010001110110000001: color_data = Z;
		19'b0010001110110000010: color_data = Z;
		19'b0010001110110000011: color_data = Z;
		19'b0010001110110000100: color_data = Z;
		19'b0010001110110000101: color_data = Z;
		19'b0010001110110000110: color_data = Z;
		19'b0010001110110000111: color_data = Z;
		19'b0010001110110001000: color_data = Z;
		19'b0010001110110001001: color_data = Z;
		19'b0010001110110001010: color_data = Z;
		19'b0010001110110001011: color_data = Z;
		19'b0010001110110001100: color_data = Z;
		19'b0010001110110001101: color_data = Z;
		19'b0010001110110001110: color_data = Z;
		19'b0010001110110001111: color_data = Z;
		19'b0010001110110010000: color_data = Z;
		19'b0010001110110010001: color_data = Z;
		19'b0010001110110010010: color_data = Z;
		19'b0010001110110010011: color_data = Z;
		19'b0010001110110010100: color_data = Z;
		19'b0010001110110010101: color_data = Z;
		19'b0010001110110010110: color_data = Z;
		19'b0010001110110010111: color_data = Z;
		19'b0010001110110011000: color_data = Z;
		19'b0010001110110011001: color_data = Z;
		19'b0010001110110011010: color_data = Z;
		19'b0010001110110011011: color_data = Z;
		19'b0010001110110011100: color_data = Z;
		19'b0010001110110011101: color_data = Z;
		19'b0010001110110011110: color_data = Z;
		19'b0010001110110011111: color_data = Z;
		19'b0010001110110100000: color_data = Z;
		19'b0010001110110100001: color_data = Z;
		19'b0010001110110100010: color_data = Z;
		19'b0010001110110100011: color_data = Z;
		19'b0010001110110100100: color_data = Z;
		19'b0010001110110100101: color_data = Z;
		19'b0010001110110100110: color_data = Z;
		19'b0010001110110100111: color_data = Z;
		19'b0010001110110101000: color_data = Z;
		19'b0010001110110101001: color_data = Z;
		19'b0010001110110101010: color_data = Z;
		19'b0010001110110101011: color_data = Z;
		19'b0010001110110110000: color_data = Z;
		19'b0010001110110110001: color_data = Z;
		19'b0010001110110110010: color_data = Z;
		19'b0010001110110110011: color_data = Z;
		19'b0010001110110111001: color_data = Z;
		19'b0010001110110111010: color_data = Z;
		19'b0010001110110111011: color_data = Z;
		19'b0010001110110111100: color_data = Z;
		19'b0010001110110111101: color_data = Z;
		19'b0010001110110111110: color_data = Z;
		19'b0010001110110111111: color_data = Z;
		19'b0010001110111000000: color_data = Z;
		19'b0010001110111000001: color_data = Z;
		19'b0010001110111000010: color_data = Z;
		19'b0010001110111000011: color_data = Z;
		19'b0010001110111000100: color_data = Z;
		19'b0010001110111000101: color_data = Z;
		19'b0010001110111000110: color_data = Z;
		19'b0010001110111000111: color_data = Z;
		19'b0010010000011001011: color_data = Z;
		19'b0010010000011001100: color_data = Z;
		19'b0010010000011001101: color_data = Z;
		19'b0010010000011001110: color_data = Z;
		19'b0010010000011001111: color_data = Z;
		19'b0010010000011010000: color_data = Z;
		19'b0010010000011010001: color_data = Z;
		19'b0010010000011010010: color_data = Z;
		19'b0010010000011010011: color_data = Z;
		19'b0010010000011010100: color_data = Z;
		19'b0010010000011010101: color_data = Z;
		19'b0010010000011010110: color_data = Z;
		19'b0010010000011010111: color_data = Z;
		19'b0010010000011011000: color_data = Z;
		19'b0010010000011011001: color_data = Z;
		19'b0010010000011011010: color_data = Z;
		19'b0010010000011011011: color_data = Z;
		19'b0010010000011011100: color_data = Z;
		19'b0010010000011011101: color_data = Z;
		19'b0010010000011011110: color_data = Z;
		19'b0010010000011011111: color_data = Z;
		19'b0010010000011100000: color_data = Z;
		19'b0010010000011100001: color_data = Z;
		19'b0010010000011100010: color_data = Z;
		19'b0010010000011100011: color_data = Z;
		19'b0010010000011100100: color_data = Z;
		19'b0010010000011100101: color_data = Z;
		19'b0010010000011100110: color_data = Z;
		19'b0010010000011100111: color_data = Z;
		19'b0010010000011101000: color_data = Z;
		19'b0010010000011101001: color_data = Z;
		19'b0010010000011101010: color_data = Z;
		19'b0010010000011101011: color_data = Z;
		19'b0010010000011101100: color_data = Z;
		19'b0010010000011101101: color_data = Z;
		19'b0010010000011101110: color_data = Z;
		19'b0010010000011101111: color_data = Z;
		19'b0010010000011110000: color_data = Z;
		19'b0010010000011110001: color_data = Z;
		19'b0010010000011110010: color_data = Z;
		19'b0010010000011110011: color_data = Z;
		19'b0010010000011110100: color_data = Z;
		19'b0010010000011110101: color_data = Z;
		19'b0010010000011110110: color_data = Z;
		19'b0010010000011110111: color_data = Z;
		19'b0010010000011111000: color_data = Z;
		19'b0010010000011111001: color_data = Z;
		19'b0010010000011111010: color_data = Z;
		19'b0010010000011111011: color_data = Z;
		19'b0010010000011111100: color_data = Z;
		19'b0010010000011111101: color_data = Z;
		19'b0010010000011111110: color_data = Z;
		19'b0010010000011111111: color_data = Z;
		19'b0010010000100000000: color_data = Z;
		19'b0010010000100000001: color_data = Z;
		19'b0010010000100000010: color_data = Z;
		19'b0010010000100000011: color_data = Z;
		19'b0010010000100000100: color_data = Z;
		19'b0010010000100000101: color_data = Z;
		19'b0010010000100000110: color_data = Z;
		19'b0010010000100000111: color_data = Z;
		19'b0010010000100001000: color_data = Z;
		19'b0010010000100001001: color_data = Z;
		19'b0010010000100001010: color_data = Z;
		19'b0010010000100001011: color_data = Z;
		19'b0010010000100001100: color_data = Z;
		19'b0010010000100001101: color_data = Z;
		19'b0010010000100001110: color_data = Z;
		19'b0010010000100001111: color_data = Z;
		19'b0010010000100010000: color_data = Z;
		19'b0010010000100010001: color_data = Z;
		19'b0010010000100010010: color_data = Z;
		19'b0010010000100010011: color_data = Z;
		19'b0010010000100010100: color_data = Z;
		19'b0010010000100010101: color_data = Z;
		19'b0010010000100010110: color_data = Z;
		19'b0010010000100010111: color_data = Z;
		19'b0010010000100011000: color_data = Z;
		19'b0010010000100011001: color_data = Z;
		19'b0010010000100011010: color_data = Z;
		19'b0010010000100011011: color_data = Z;
		19'b0010010000100011100: color_data = Z;
		19'b0010010000100011101: color_data = Z;
		19'b0010010000100011110: color_data = Z;
		19'b0010010000100011111: color_data = Z;
		19'b0010010000100100000: color_data = Z;
		19'b0010010000100100001: color_data = Z;
		19'b0010010000100100010: color_data = Z;
		19'b0010010000100100011: color_data = Z;
		19'b0010010000100100100: color_data = Z;
		19'b0010010000100100101: color_data = Z;
		19'b0010010000100100110: color_data = Z;
		19'b0010010000100100111: color_data = Z;
		19'b0010010000100101000: color_data = Z;
		19'b0010010000100101001: color_data = Z;
		19'b0010010000100101010: color_data = Z;
		19'b0010010000100101011: color_data = Z;
		19'b0010010000100101100: color_data = Z;
		19'b0010010000100101101: color_data = Z;
		19'b0010010000100101110: color_data = Z;
		19'b0010010000100101111: color_data = Z;
		19'b0010010000100110000: color_data = Z;
		19'b0010010000100110001: color_data = Z;
		19'b0010010000100110010: color_data = Z;
		19'b0010010000100110011: color_data = Z;
		19'b0010010000100110100: color_data = Z;
		19'b0010010000100110101: color_data = Z;
		19'b0010010000100110110: color_data = Z;
		19'b0010010000100110111: color_data = Z;
		19'b0010010000100111000: color_data = Z;
		19'b0010010000100111001: color_data = Z;
		19'b0010010000100111010: color_data = Z;
		19'b0010010000100111011: color_data = Z;
		19'b0010010000100111100: color_data = Z;
		19'b0010010000100111101: color_data = Z;
		19'b0010010000100111110: color_data = Z;
		19'b0010010000100111111: color_data = Z;
		19'b0010010000101000000: color_data = Z;
		19'b0010010000101000001: color_data = Z;
		19'b0010010000101000010: color_data = Z;
		19'b0010010000101000011: color_data = Z;
		19'b0010010000101000100: color_data = Z;
		19'b0010010000101000101: color_data = Z;
		19'b0010010000101000110: color_data = Z;
		19'b0010010000101000111: color_data = Z;
		19'b0010010000101001000: color_data = Z;
		19'b0010010000101001001: color_data = Z;
		19'b0010010000101001010: color_data = Z;
		19'b0010010000101001011: color_data = Z;
		19'b0010010000101001100: color_data = Z;
		19'b0010010000101001101: color_data = Z;
		19'b0010010000101001110: color_data = Z;
		19'b0010010000101001111: color_data = Z;
		19'b0010010000101010000: color_data = Z;
		19'b0010010000101010001: color_data = Z;
		19'b0010010000101010010: color_data = Z;
		19'b0010010000101010011: color_data = Z;
		19'b0010010000101010100: color_data = Z;
		19'b0010010000101010101: color_data = Z;
		19'b0010010000101010110: color_data = Z;
		19'b0010010000101010111: color_data = Z;
		19'b0010010000101011000: color_data = Z;
		19'b0010010000101011001: color_data = Z;
		19'b0010010000101011010: color_data = Z;
		19'b0010010000101011011: color_data = Z;
		19'b0010010000101011100: color_data = Z;
		19'b0010010000101011101: color_data = Z;
		19'b0010010000101011110: color_data = Z;
		19'b0010010000101011111: color_data = Z;
		19'b0010010000101100000: color_data = Z;
		19'b0010010000101100001: color_data = Z;
		19'b0010010000101100010: color_data = Z;
		19'b0010010000101100011: color_data = Z;
		19'b0010010000101100100: color_data = Z;
		19'b0010010000101100101: color_data = Z;
		19'b0010010000101100110: color_data = Z;
		19'b0010010000101100111: color_data = Z;
		19'b0010010000101101000: color_data = Z;
		19'b0010010000101101001: color_data = Z;
		19'b0010010000101101010: color_data = Z;
		19'b0010010000101101011: color_data = Z;
		19'b0010010000101101100: color_data = Z;
		19'b0010010000101101101: color_data = Z;
		19'b0010010000101101110: color_data = Z;
		19'b0010010000101101111: color_data = Z;
		19'b0010010000101110000: color_data = Z;
		19'b0010010000101110001: color_data = Z;
		19'b0010010000101110010: color_data = Z;
		19'b0010010000101110011: color_data = Z;
		19'b0010010000101110100: color_data = Z;
		19'b0010010000101110101: color_data = Z;
		19'b0010010000101110110: color_data = Z;
		19'b0010010000101110111: color_data = Z;
		19'b0010010000101111000: color_data = Z;
		19'b0010010000101111001: color_data = Z;
		19'b0010010000101111010: color_data = Z;
		19'b0010010000101111011: color_data = Z;
		19'b0010010000101111100: color_data = Z;
		19'b0010010000101111101: color_data = Z;
		19'b0010010000101111110: color_data = Z;
		19'b0010010000101111111: color_data = Z;
		19'b0010010000110000000: color_data = Z;
		19'b0010010000110000001: color_data = Z;
		19'b0010010000110000010: color_data = Z;
		19'b0010010000110000011: color_data = Z;
		19'b0010010000110000100: color_data = Z;
		19'b0010010000110000101: color_data = Z;
		19'b0010010000110000110: color_data = Z;
		19'b0010010000110000111: color_data = Z;
		19'b0010010000110001000: color_data = Z;
		19'b0010010000110001001: color_data = Z;
		19'b0010010000110001010: color_data = Z;
		19'b0010010000110001011: color_data = Z;
		19'b0010010000110001100: color_data = Z;
		19'b0010010000110001101: color_data = Z;
		19'b0010010000110001110: color_data = Z;
		19'b0010010000110001111: color_data = Z;
		19'b0010010000110010000: color_data = Z;
		19'b0010010000110010001: color_data = Z;
		19'b0010010000110010010: color_data = Z;
		19'b0010010000110010011: color_data = Z;
		19'b0010010000110010100: color_data = Z;
		19'b0010010000110010101: color_data = Z;
		19'b0010010000110010110: color_data = Z;
		19'b0010010000110010111: color_data = Z;
		19'b0010010000110011000: color_data = Z;
		19'b0010010000110011001: color_data = Z;
		19'b0010010000110011010: color_data = Z;
		19'b0010010000110011011: color_data = Z;
		19'b0010010000110011100: color_data = Z;
		19'b0010010000110011101: color_data = Z;
		19'b0010010000110011110: color_data = Z;
		19'b0010010000110011111: color_data = Z;
		19'b0010010000110100000: color_data = Z;
		19'b0010010000110100001: color_data = Z;
		19'b0010010000110100010: color_data = Z;
		19'b0010010000110100011: color_data = Z;
		19'b0010010000110100100: color_data = Z;
		19'b0010010000110100101: color_data = Z;
		19'b0010010000110100110: color_data = Z;
		19'b0010010000110100111: color_data = Z;
		19'b0010010000110101000: color_data = Z;
		19'b0010010000110101001: color_data = Z;
		19'b0010010000110101010: color_data = Z;
		19'b0010010000110101011: color_data = Z;
		19'b0010010000110110000: color_data = Z;
		19'b0010010000110110001: color_data = Z;
		19'b0010010000110110010: color_data = Z;
		19'b0010010000110110011: color_data = Z;
		19'b0010010000110110100: color_data = Z;
		19'b0010010000110111010: color_data = Z;
		19'b0010010000110111011: color_data = Z;
		19'b0010010000110111100: color_data = Z;
		19'b0010010000110111101: color_data = Z;
		19'b0010010000110111110: color_data = Z;
		19'b0010010000110111111: color_data = Z;
		19'b0010010000111000000: color_data = Z;
		19'b0010010000111000001: color_data = Z;
		19'b0010010000111000010: color_data = Z;
		19'b0010010000111000011: color_data = Z;
		19'b0010010000111000100: color_data = Z;
		19'b0010010000111000101: color_data = Z;
		19'b0010010000111000110: color_data = Z;
		19'b0010010000111000111: color_data = Z;
		19'b0010010000111001000: color_data = Z;
		19'b0010010010011001011: color_data = Z;
		19'b0010010010011001100: color_data = Z;
		19'b0010010010011001101: color_data = Z;
		19'b0010010010011001110: color_data = Z;
		19'b0010010010011001111: color_data = Z;
		19'b0010010010011010000: color_data = Z;
		19'b0010010010011010001: color_data = Z;
		19'b0010010010011010010: color_data = Z;
		19'b0010010010011010011: color_data = Z;
		19'b0010010010011010100: color_data = Z;
		19'b0010010010011010101: color_data = Z;
		19'b0010010010011010110: color_data = Z;
		19'b0010010010011010111: color_data = Z;
		19'b0010010010011011000: color_data = Z;
		19'b0010010010011011001: color_data = Z;
		19'b0010010010011011010: color_data = Z;
		19'b0010010010011011011: color_data = Z;
		19'b0010010010011011100: color_data = Z;
		19'b0010010010011011101: color_data = Z;
		19'b0010010010011011110: color_data = Z;
		19'b0010010010011011111: color_data = Z;
		19'b0010010010011100000: color_data = Z;
		19'b0010010010011100001: color_data = Z;
		19'b0010010010011100010: color_data = Z;
		19'b0010010010011100011: color_data = Z;
		19'b0010010010011100100: color_data = Z;
		19'b0010010010011100101: color_data = Z;
		19'b0010010010011100110: color_data = Z;
		19'b0010010010011100111: color_data = Z;
		19'b0010010010011101000: color_data = Z;
		19'b0010010010011101001: color_data = Z;
		19'b0010010010011101010: color_data = Z;
		19'b0010010010011101011: color_data = Z;
		19'b0010010010011101100: color_data = Z;
		19'b0010010010011101101: color_data = Z;
		19'b0010010010011101110: color_data = Z;
		19'b0010010010011101111: color_data = Z;
		19'b0010010010011110000: color_data = Z;
		19'b0010010010011110001: color_data = Z;
		19'b0010010010011110010: color_data = Z;
		19'b0010010010011110011: color_data = Z;
		19'b0010010010011110100: color_data = Z;
		19'b0010010010011110101: color_data = Z;
		19'b0010010010011110110: color_data = Z;
		19'b0010010010011110111: color_data = Z;
		19'b0010010010011111000: color_data = Z;
		19'b0010010010011111001: color_data = Z;
		19'b0010010010011111010: color_data = Z;
		19'b0010010010011111011: color_data = Z;
		19'b0010010010011111100: color_data = Z;
		19'b0010010010011111101: color_data = Z;
		19'b0010010010011111110: color_data = Z;
		19'b0010010010011111111: color_data = Z;
		19'b0010010010100000000: color_data = Z;
		19'b0010010010100000001: color_data = Z;
		19'b0010010010100000010: color_data = Z;
		19'b0010010010100000011: color_data = Z;
		19'b0010010010100000100: color_data = Z;
		19'b0010010010100000101: color_data = Z;
		19'b0010010010100000110: color_data = Z;
		19'b0010010010100000111: color_data = Z;
		19'b0010010010100001000: color_data = Z;
		19'b0010010010100001001: color_data = Z;
		19'b0010010010100001010: color_data = Z;
		19'b0010010010100001011: color_data = Z;
		19'b0010010010100001100: color_data = Z;
		19'b0010010010100001101: color_data = Z;
		19'b0010010010100001110: color_data = Z;
		19'b0010010010100001111: color_data = Z;
		19'b0010010010100010000: color_data = Z;
		19'b0010010010100010001: color_data = Z;
		19'b0010010010100010010: color_data = Z;
		19'b0010010010100010011: color_data = Z;
		19'b0010010010100010100: color_data = Z;
		19'b0010010010100010101: color_data = Z;
		19'b0010010010100010110: color_data = Z;
		19'b0010010010100010111: color_data = Z;
		19'b0010010010100011000: color_data = Z;
		19'b0010010010100011001: color_data = Z;
		19'b0010010010100011010: color_data = Z;
		19'b0010010010100011011: color_data = Z;
		19'b0010010010100011100: color_data = Z;
		19'b0010010010100011101: color_data = Z;
		19'b0010010010100011110: color_data = Z;
		19'b0010010010100011111: color_data = Z;
		19'b0010010010100100000: color_data = Z;
		19'b0010010010100100001: color_data = Z;
		19'b0010010010100100010: color_data = Z;
		19'b0010010010100100011: color_data = Z;
		19'b0010010010100100100: color_data = Z;
		19'b0010010010100100101: color_data = Z;
		19'b0010010010100100110: color_data = Z;
		19'b0010010010100100111: color_data = Z;
		19'b0010010010100101000: color_data = Z;
		19'b0010010010100101001: color_data = Z;
		19'b0010010010100101010: color_data = Z;
		19'b0010010010100101011: color_data = Z;
		19'b0010010010100101100: color_data = Z;
		19'b0010010010100101101: color_data = Z;
		19'b0010010010100101110: color_data = Z;
		19'b0010010010100101111: color_data = Z;
		19'b0010010010100110000: color_data = Z;
		19'b0010010010100110001: color_data = Z;
		19'b0010010010100110010: color_data = Z;
		19'b0010010010100110011: color_data = Z;
		19'b0010010010100110100: color_data = Z;
		19'b0010010010100110101: color_data = Z;
		19'b0010010010100110110: color_data = Z;
		19'b0010010010100110111: color_data = Z;
		19'b0010010010100111000: color_data = Z;
		19'b0010010010100111001: color_data = Z;
		19'b0010010010100111010: color_data = Z;
		19'b0010010010100111011: color_data = Z;
		19'b0010010010100111100: color_data = Z;
		19'b0010010010100111101: color_data = Z;
		19'b0010010010100111110: color_data = Z;
		19'b0010010010100111111: color_data = Z;
		19'b0010010010101000000: color_data = Z;
		19'b0010010010101000001: color_data = Z;
		19'b0010010010101000010: color_data = Z;
		19'b0010010010101000011: color_data = Z;
		19'b0010010010101000100: color_data = Z;
		19'b0010010010101000101: color_data = Z;
		19'b0010010010101000110: color_data = Z;
		19'b0010010010101000111: color_data = Z;
		19'b0010010010101001000: color_data = Z;
		19'b0010010010101001001: color_data = Z;
		19'b0010010010101001010: color_data = Z;
		19'b0010010010101001011: color_data = Z;
		19'b0010010010101001100: color_data = Z;
		19'b0010010010101001101: color_data = Z;
		19'b0010010010101001110: color_data = Z;
		19'b0010010010101001111: color_data = Z;
		19'b0010010010101010000: color_data = Z;
		19'b0010010010101010001: color_data = Z;
		19'b0010010010101010010: color_data = Z;
		19'b0010010010101010011: color_data = Z;
		19'b0010010010101010100: color_data = Z;
		19'b0010010010101010101: color_data = Z;
		19'b0010010010101010110: color_data = Z;
		19'b0010010010101010111: color_data = Z;
		19'b0010010010101011000: color_data = Z;
		19'b0010010010101011001: color_data = Z;
		19'b0010010010101011010: color_data = Z;
		19'b0010010010101011011: color_data = Z;
		19'b0010010010101011100: color_data = Z;
		19'b0010010010101011101: color_data = Z;
		19'b0010010010101011110: color_data = Z;
		19'b0010010010101011111: color_data = Z;
		19'b0010010010101100000: color_data = Z;
		19'b0010010010101100001: color_data = Z;
		19'b0010010010101100010: color_data = Z;
		19'b0010010010101100011: color_data = Z;
		19'b0010010010101100100: color_data = Z;
		19'b0010010010101100101: color_data = Z;
		19'b0010010010101100110: color_data = Z;
		19'b0010010010101100111: color_data = Z;
		19'b0010010010101101000: color_data = Z;
		19'b0010010010101101001: color_data = Z;
		19'b0010010010101101010: color_data = Z;
		19'b0010010010101101011: color_data = Z;
		19'b0010010010101101100: color_data = Z;
		19'b0010010010101101101: color_data = Z;
		19'b0010010010101101110: color_data = Z;
		19'b0010010010101101111: color_data = Z;
		19'b0010010010101110000: color_data = Z;
		19'b0010010010101110001: color_data = Z;
		19'b0010010010101110010: color_data = Z;
		19'b0010010010101110011: color_data = Z;
		19'b0010010010101110100: color_data = Z;
		19'b0010010010101110101: color_data = Z;
		19'b0010010010101110110: color_data = Z;
		19'b0010010010101110111: color_data = Z;
		19'b0010010010101111000: color_data = Z;
		19'b0010010010101111001: color_data = Z;
		19'b0010010010101111010: color_data = Z;
		19'b0010010010101111011: color_data = Z;
		19'b0010010010101111100: color_data = Z;
		19'b0010010010101111101: color_data = Z;
		19'b0010010010101111110: color_data = Z;
		19'b0010010010101111111: color_data = Z;
		19'b0010010010110000000: color_data = Z;
		19'b0010010010110000001: color_data = Z;
		19'b0010010010110000010: color_data = Z;
		19'b0010010010110000011: color_data = Z;
		19'b0010010010110000100: color_data = Z;
		19'b0010010010110000101: color_data = Z;
		19'b0010010010110000110: color_data = Z;
		19'b0010010010110000111: color_data = Z;
		19'b0010010010110001000: color_data = Z;
		19'b0010010010110001001: color_data = Z;
		19'b0010010010110001010: color_data = Z;
		19'b0010010010110001011: color_data = Z;
		19'b0010010010110001100: color_data = Z;
		19'b0010010010110001101: color_data = Z;
		19'b0010010010110001110: color_data = Z;
		19'b0010010010110001111: color_data = Z;
		19'b0010010010110010000: color_data = Z;
		19'b0010010010110010001: color_data = Z;
		19'b0010010010110010010: color_data = Z;
		19'b0010010010110010011: color_data = Z;
		19'b0010010010110010100: color_data = Z;
		19'b0010010010110010101: color_data = Z;
		19'b0010010010110010110: color_data = Z;
		19'b0010010010110010111: color_data = Z;
		19'b0010010010110011000: color_data = Z;
		19'b0010010010110011001: color_data = Z;
		19'b0010010010110011010: color_data = Z;
		19'b0010010010110011011: color_data = Z;
		19'b0010010010110011100: color_data = Z;
		19'b0010010010110011101: color_data = Z;
		19'b0010010010110011110: color_data = Z;
		19'b0010010010110011111: color_data = Z;
		19'b0010010010110100000: color_data = Z;
		19'b0010010010110100001: color_data = Z;
		19'b0010010010110100010: color_data = Z;
		19'b0010010010110100011: color_data = Z;
		19'b0010010010110100100: color_data = Z;
		19'b0010010010110100101: color_data = Z;
		19'b0010010010110100110: color_data = Z;
		19'b0010010010110100111: color_data = Z;
		19'b0010010010110101000: color_data = Z;
		19'b0010010010110101001: color_data = Z;
		19'b0010010010110101010: color_data = Z;
		19'b0010010010110101011: color_data = Z;
		19'b0010010010110110001: color_data = Z;
		19'b0010010010110110010: color_data = Z;
		19'b0010010010110110011: color_data = Z;
		19'b0010010010110110100: color_data = Z;
		19'b0010010010110110101: color_data = Z;
		19'b0010010010110111010: color_data = Z;
		19'b0010010010110111011: color_data = Z;
		19'b0010010010110111100: color_data = Z;
		19'b0010010010110111101: color_data = Z;
		19'b0010010010110111110: color_data = Z;
		19'b0010010010110111111: color_data = Z;
		19'b0010010010111000000: color_data = Z;
		19'b0010010010111000001: color_data = Z;
		19'b0010010010111000010: color_data = Z;
		19'b0010010010111000011: color_data = Z;
		19'b0010010010111000100: color_data = Z;
		19'b0010010010111000101: color_data = Z;
		19'b0010010010111000110: color_data = Z;
		19'b0010010010111000111: color_data = Z;
		19'b0010010100011001010: color_data = Z;
		19'b0010010100011001011: color_data = Z;
		19'b0010010100011001100: color_data = Z;
		19'b0010010100011001101: color_data = Z;
		19'b0010010100011001110: color_data = Z;
		19'b0010010100011001111: color_data = Z;
		19'b0010010100011010000: color_data = Z;
		19'b0010010100011010001: color_data = Z;
		19'b0010010100011010010: color_data = Z;
		19'b0010010100011010011: color_data = Z;
		19'b0010010100011010100: color_data = Z;
		19'b0010010100011010101: color_data = Z;
		19'b0010010100011010110: color_data = Z;
		19'b0010010100011010111: color_data = Z;
		19'b0010010100011011000: color_data = Z;
		19'b0010010100011011001: color_data = Z;
		19'b0010010100011011010: color_data = Z;
		19'b0010010100011011011: color_data = Z;
		19'b0010010100011011100: color_data = Z;
		19'b0010010100011011101: color_data = Z;
		19'b0010010100011011110: color_data = Z;
		19'b0010010100011011111: color_data = Z;
		19'b0010010100011100000: color_data = Z;
		19'b0010010100011100001: color_data = Z;
		19'b0010010100011100010: color_data = Z;
		19'b0010010100011100011: color_data = Z;
		19'b0010010100011100100: color_data = Z;
		19'b0010010100011100101: color_data = Z;
		19'b0010010100011100110: color_data = Z;
		19'b0010010100011100111: color_data = Z;
		19'b0010010100011101000: color_data = Z;
		19'b0010010100011101001: color_data = Z;
		19'b0010010100011101010: color_data = Z;
		19'b0010010100011101011: color_data = Z;
		19'b0010010100011101100: color_data = Z;
		19'b0010010100011101101: color_data = Z;
		19'b0010010100011101110: color_data = Z;
		19'b0010010100011101111: color_data = Z;
		19'b0010010100011110000: color_data = Z;
		19'b0010010100011110001: color_data = Z;
		19'b0010010100011110010: color_data = Z;
		19'b0010010100011110011: color_data = Z;
		19'b0010010100011110100: color_data = Z;
		19'b0010010100011110101: color_data = Z;
		19'b0010010100011110110: color_data = Z;
		19'b0010010100011110111: color_data = Z;
		19'b0010010100011111000: color_data = Z;
		19'b0010010100011111001: color_data = Z;
		19'b0010010100011111010: color_data = Z;
		19'b0010010100011111011: color_data = Z;
		19'b0010010100011111100: color_data = Z;
		19'b0010010100011111101: color_data = Z;
		19'b0010010100011111110: color_data = Z;
		19'b0010010100011111111: color_data = Z;
		19'b0010010100100000000: color_data = Z;
		19'b0010010100100000001: color_data = Z;
		19'b0010010100100000010: color_data = Z;
		19'b0010010100100000011: color_data = Z;
		19'b0010010100100000100: color_data = Z;
		19'b0010010100100000101: color_data = Z;
		19'b0010010100100000110: color_data = Z;
		19'b0010010100100000111: color_data = Z;
		19'b0010010100100001000: color_data = Z;
		19'b0010010100100001001: color_data = Z;
		19'b0010010100100001010: color_data = Z;
		19'b0010010100100001011: color_data = Z;
		19'b0010010100100001100: color_data = Z;
		19'b0010010100100001101: color_data = Z;
		19'b0010010100100001110: color_data = Z;
		19'b0010010100100001111: color_data = Z;
		19'b0010010100100010000: color_data = Z;
		19'b0010010100100010001: color_data = Z;
		19'b0010010100100010010: color_data = Z;
		19'b0010010100100010011: color_data = Z;
		19'b0010010100100010100: color_data = Z;
		19'b0010010100100010101: color_data = Z;
		19'b0010010100100010110: color_data = Z;
		19'b0010010100100010111: color_data = Z;
		19'b0010010100100011000: color_data = Z;
		19'b0010010100100011001: color_data = Z;
		19'b0010010100100011010: color_data = Z;
		19'b0010010100100011011: color_data = Z;
		19'b0010010100100011100: color_data = Z;
		19'b0010010100100011101: color_data = Z;
		19'b0010010100100011110: color_data = Z;
		19'b0010010100100011111: color_data = Z;
		19'b0010010100100100000: color_data = Z;
		19'b0010010100100100001: color_data = Z;
		19'b0010010100100100010: color_data = Z;
		19'b0010010100100100011: color_data = Z;
		19'b0010010100100100100: color_data = Z;
		19'b0010010100100100101: color_data = Z;
		19'b0010010100100100110: color_data = Z;
		19'b0010010100100100111: color_data = Z;
		19'b0010010100100101000: color_data = Z;
		19'b0010010100100101001: color_data = Z;
		19'b0010010100100101010: color_data = Z;
		19'b0010010100100101011: color_data = Z;
		19'b0010010100100101100: color_data = Z;
		19'b0010010100100101101: color_data = Z;
		19'b0010010100100101110: color_data = Z;
		19'b0010010100100101111: color_data = Z;
		19'b0010010100100110000: color_data = Z;
		19'b0010010100100110001: color_data = Z;
		19'b0010010100100110010: color_data = Z;
		19'b0010010100100110011: color_data = Z;
		19'b0010010100100110100: color_data = Z;
		19'b0010010100100110101: color_data = Z;
		19'b0010010100100110110: color_data = Z;
		19'b0010010100100110111: color_data = Z;
		19'b0010010100100111000: color_data = Z;
		19'b0010010100100111001: color_data = Z;
		19'b0010010100100111010: color_data = Z;
		19'b0010010100100111011: color_data = Z;
		19'b0010010100100111100: color_data = Z;
		19'b0010010100100111101: color_data = Z;
		19'b0010010100100111110: color_data = Z;
		19'b0010010100100111111: color_data = Z;
		19'b0010010100101000000: color_data = Z;
		19'b0010010100101000001: color_data = Z;
		19'b0010010100101000010: color_data = Z;
		19'b0010010100101000011: color_data = Z;
		19'b0010010100101000100: color_data = Z;
		19'b0010010100101000101: color_data = Z;
		19'b0010010100101000110: color_data = Z;
		19'b0010010100101000111: color_data = Z;
		19'b0010010100101001000: color_data = Z;
		19'b0010010100101001001: color_data = Z;
		19'b0010010100101001010: color_data = Z;
		19'b0010010100101001011: color_data = Z;
		19'b0010010100101001100: color_data = Z;
		19'b0010010100101001101: color_data = Z;
		19'b0010010100101001110: color_data = Z;
		19'b0010010100101001111: color_data = Z;
		19'b0010010100101010000: color_data = Z;
		19'b0010010100101010001: color_data = Z;
		19'b0010010100101010010: color_data = Z;
		19'b0010010100101010011: color_data = Z;
		19'b0010010100101010100: color_data = Z;
		19'b0010010100101010101: color_data = Z;
		19'b0010010100101010110: color_data = Z;
		19'b0010010100101010111: color_data = Z;
		19'b0010010100101011000: color_data = Z;
		19'b0010010100101011001: color_data = Z;
		19'b0010010100101011010: color_data = Z;
		19'b0010010100101011011: color_data = Z;
		19'b0010010100101011100: color_data = Z;
		19'b0010010100101011101: color_data = Z;
		19'b0010010100101011110: color_data = Z;
		19'b0010010100101011111: color_data = Z;
		19'b0010010100101100000: color_data = Z;
		19'b0010010100101100001: color_data = Z;
		19'b0010010100101100010: color_data = Z;
		19'b0010010100101100011: color_data = Z;
		19'b0010010100101100100: color_data = Z;
		19'b0010010100101100101: color_data = Z;
		19'b0010010100101100110: color_data = Z;
		19'b0010010100101100111: color_data = Z;
		19'b0010010100101101000: color_data = Z;
		19'b0010010100101101001: color_data = Z;
		19'b0010010100101101010: color_data = Z;
		19'b0010010100101101011: color_data = Z;
		19'b0010010100101101100: color_data = Z;
		19'b0010010100101101101: color_data = Z;
		19'b0010010100101101110: color_data = Z;
		19'b0010010100101101111: color_data = Z;
		19'b0010010100101110000: color_data = Z;
		19'b0010010100101110001: color_data = Z;
		19'b0010010100101110010: color_data = Z;
		19'b0010010100101110011: color_data = Z;
		19'b0010010100101110100: color_data = Z;
		19'b0010010100101110101: color_data = Z;
		19'b0010010100101110110: color_data = Z;
		19'b0010010100101110111: color_data = Z;
		19'b0010010100101111000: color_data = Z;
		19'b0010010100101111001: color_data = Z;
		19'b0010010100101111010: color_data = Z;
		19'b0010010100101111011: color_data = Z;
		19'b0010010100101111100: color_data = Z;
		19'b0010010100101111101: color_data = Z;
		19'b0010010100101111110: color_data = Z;
		19'b0010010100101111111: color_data = Z;
		19'b0010010100110000000: color_data = Z;
		19'b0010010100110000001: color_data = Z;
		19'b0010010100110000010: color_data = Z;
		19'b0010010100110000011: color_data = Z;
		19'b0010010100110000100: color_data = Z;
		19'b0010010100110000101: color_data = Z;
		19'b0010010100110000110: color_data = Z;
		19'b0010010100110000111: color_data = Z;
		19'b0010010100110001000: color_data = Z;
		19'b0010010100110001001: color_data = Z;
		19'b0010010100110001010: color_data = Z;
		19'b0010010100110001011: color_data = Z;
		19'b0010010100110001100: color_data = Z;
		19'b0010010100110001101: color_data = Z;
		19'b0010010100110001110: color_data = Z;
		19'b0010010100110001111: color_data = Z;
		19'b0010010100110010000: color_data = Z;
		19'b0010010100110010001: color_data = Z;
		19'b0010010100110010010: color_data = Z;
		19'b0010010100110010011: color_data = Z;
		19'b0010010100110010100: color_data = Z;
		19'b0010010100110010101: color_data = Z;
		19'b0010010100110010110: color_data = Z;
		19'b0010010100110010111: color_data = Z;
		19'b0010010100110011000: color_data = Z;
		19'b0010010100110011001: color_data = Z;
		19'b0010010100110011010: color_data = Z;
		19'b0010010100110011011: color_data = Z;
		19'b0010010100110011100: color_data = Z;
		19'b0010010100110011101: color_data = Z;
		19'b0010010100110011110: color_data = Z;
		19'b0010010100110011111: color_data = Z;
		19'b0010010100110100000: color_data = Z;
		19'b0010010100110100001: color_data = Z;
		19'b0010010100110100010: color_data = Z;
		19'b0010010100110100011: color_data = Z;
		19'b0010010100110100100: color_data = Z;
		19'b0010010100110100101: color_data = Z;
		19'b0010010100110100110: color_data = Z;
		19'b0010010100110100111: color_data = Z;
		19'b0010010100110101000: color_data = Z;
		19'b0010010100110101001: color_data = Z;
		19'b0010010100110101010: color_data = Z;
		19'b0010010100110101011: color_data = Z;
		19'b0010010100110101100: color_data = Z;
		19'b0010010100110110001: color_data = Z;
		19'b0010010100110110010: color_data = Z;
		19'b0010010100110110100: color_data = Z;
		19'b0010010100110110101: color_data = Z;
		19'b0010010100110110110: color_data = Z;
		19'b0010010100110111011: color_data = Z;
		19'b0010010100110111100: color_data = Z;
		19'b0010010100110111101: color_data = Z;
		19'b0010010100110111110: color_data = Z;
		19'b0010010100110111111: color_data = Z;
		19'b0010010100111000000: color_data = Z;
		19'b0010010100111000001: color_data = Z;
		19'b0010010100111000010: color_data = Z;
		19'b0010010100111000011: color_data = Z;
		19'b0010010100111000100: color_data = Z;
		19'b0010010100111000101: color_data = Z;
		19'b0010010100111000110: color_data = Z;
		19'b0010010100111000111: color_data = Z;
		19'b0010010100111001000: color_data = Z;
		19'b0010010110011001010: color_data = Z;
		19'b0010010110011001011: color_data = Z;
		19'b0010010110011001100: color_data = Z;
		19'b0010010110011001101: color_data = Z;
		19'b0010010110011001110: color_data = Z;
		19'b0010010110011001111: color_data = Z;
		19'b0010010110011010000: color_data = Z;
		19'b0010010110011010001: color_data = Z;
		19'b0010010110011010010: color_data = Z;
		19'b0010010110011010011: color_data = Z;
		19'b0010010110011010100: color_data = Z;
		19'b0010010110011010101: color_data = Z;
		19'b0010010110011010110: color_data = Z;
		19'b0010010110011010111: color_data = Z;
		19'b0010010110011011000: color_data = Z;
		19'b0010010110011011001: color_data = Z;
		19'b0010010110011011010: color_data = Z;
		19'b0010010110011011011: color_data = Z;
		19'b0010010110011011100: color_data = Z;
		19'b0010010110011011101: color_data = Z;
		19'b0010010110011011110: color_data = Z;
		19'b0010010110011011111: color_data = Z;
		19'b0010010110011100000: color_data = Z;
		19'b0010010110011100001: color_data = Z;
		19'b0010010110011100010: color_data = Z;
		19'b0010010110011100011: color_data = Z;
		19'b0010010110011100100: color_data = Z;
		19'b0010010110011100101: color_data = Z;
		19'b0010010110011100110: color_data = Z;
		19'b0010010110011100111: color_data = Z;
		19'b0010010110011101000: color_data = Z;
		19'b0010010110011101001: color_data = Z;
		19'b0010010110011101010: color_data = Z;
		19'b0010010110011101011: color_data = Z;
		19'b0010010110011101100: color_data = Z;
		19'b0010010110011101101: color_data = Z;
		19'b0010010110011101110: color_data = Z;
		19'b0010010110011101111: color_data = Z;
		19'b0010010110011110000: color_data = Z;
		19'b0010010110011110001: color_data = Z;
		19'b0010010110011110010: color_data = Z;
		19'b0010010110011110011: color_data = Z;
		19'b0010010110011110100: color_data = Z;
		19'b0010010110011110101: color_data = Z;
		19'b0010010110011110110: color_data = Z;
		19'b0010010110011110111: color_data = Z;
		19'b0010010110011111000: color_data = Z;
		19'b0010010110011111001: color_data = Z;
		19'b0010010110011111010: color_data = Z;
		19'b0010010110011111011: color_data = Z;
		19'b0010010110011111100: color_data = Z;
		19'b0010010110011111101: color_data = Z;
		19'b0010010110011111110: color_data = Z;
		19'b0010010110011111111: color_data = Z;
		19'b0010010110100000000: color_data = Z;
		19'b0010010110100000001: color_data = Z;
		19'b0010010110100000010: color_data = Z;
		19'b0010010110100000011: color_data = Z;
		19'b0010010110100000100: color_data = Z;
		19'b0010010110100000101: color_data = Z;
		19'b0010010110100000110: color_data = Z;
		19'b0010010110100000111: color_data = Z;
		19'b0010010110100001000: color_data = Z;
		19'b0010010110100001001: color_data = Z;
		19'b0010010110100001010: color_data = Z;
		19'b0010010110100001011: color_data = Z;
		19'b0010010110100001100: color_data = Z;
		19'b0010010110100001101: color_data = Z;
		19'b0010010110100001110: color_data = Z;
		19'b0010010110100001111: color_data = Z;
		19'b0010010110100010000: color_data = Z;
		19'b0010010110100010001: color_data = Z;
		19'b0010010110100010010: color_data = Z;
		19'b0010010110100010011: color_data = Z;
		19'b0010010110100010100: color_data = Z;
		19'b0010010110100010101: color_data = Z;
		19'b0010010110100010110: color_data = Z;
		19'b0010010110100010111: color_data = Z;
		19'b0010010110100011000: color_data = Z;
		19'b0010010110100011001: color_data = Z;
		19'b0010010110100011010: color_data = Z;
		19'b0010010110100011011: color_data = Z;
		19'b0010010110100011100: color_data = Z;
		19'b0010010110100011101: color_data = Z;
		19'b0010010110100011110: color_data = Z;
		19'b0010010110100011111: color_data = Z;
		19'b0010010110100100000: color_data = Z;
		19'b0010010110100100001: color_data = Z;
		19'b0010010110100100010: color_data = Z;
		19'b0010010110100100011: color_data = Z;
		19'b0010010110100100100: color_data = Z;
		19'b0010010110100100101: color_data = Z;
		19'b0010010110100100110: color_data = Z;
		19'b0010010110100100111: color_data = Z;
		19'b0010010110100101000: color_data = Z;
		19'b0010010110100101001: color_data = Z;
		19'b0010010110100101010: color_data = Z;
		19'b0010010110100101011: color_data = Z;
		19'b0010010110100101100: color_data = Z;
		19'b0010010110100101101: color_data = Z;
		19'b0010010110100101110: color_data = Z;
		19'b0010010110100101111: color_data = Z;
		19'b0010010110100110000: color_data = Z;
		19'b0010010110100110001: color_data = Z;
		19'b0010010110100110010: color_data = Z;
		19'b0010010110100110011: color_data = Z;
		19'b0010010110100110100: color_data = Z;
		19'b0010010110100110101: color_data = Z;
		19'b0010010110100110110: color_data = Z;
		19'b0010010110100110111: color_data = Z;
		19'b0010010110100111000: color_data = Z;
		19'b0010010110100111001: color_data = Z;
		19'b0010010110100111010: color_data = Z;
		19'b0010010110100111011: color_data = Z;
		19'b0010010110100111100: color_data = Z;
		19'b0010010110100111101: color_data = Z;
		19'b0010010110100111110: color_data = Z;
		19'b0010010110100111111: color_data = Z;
		19'b0010010110101000000: color_data = Z;
		19'b0010010110101000001: color_data = Z;
		19'b0010010110101000010: color_data = Z;
		19'b0010010110101000011: color_data = Z;
		19'b0010010110101000100: color_data = Z;
		19'b0010010110101000101: color_data = Z;
		19'b0010010110101000110: color_data = Z;
		19'b0010010110101000111: color_data = Z;
		19'b0010010110101001000: color_data = Z;
		19'b0010010110101001001: color_data = Z;
		19'b0010010110101001010: color_data = Z;
		19'b0010010110101001011: color_data = Z;
		19'b0010010110101001100: color_data = Z;
		19'b0010010110101001101: color_data = Z;
		19'b0010010110101001110: color_data = Z;
		19'b0010010110101001111: color_data = Z;
		19'b0010010110101010000: color_data = Z;
		19'b0010010110101010001: color_data = Z;
		19'b0010010110101010010: color_data = Z;
		19'b0010010110101010011: color_data = Z;
		19'b0010010110101010100: color_data = Z;
		19'b0010010110101010101: color_data = Z;
		19'b0010010110101010110: color_data = Z;
		19'b0010010110101010111: color_data = Z;
		19'b0010010110101011000: color_data = Z;
		19'b0010010110101011001: color_data = Z;
		19'b0010010110101011010: color_data = Z;
		19'b0010010110101011011: color_data = Z;
		19'b0010010110101011100: color_data = Z;
		19'b0010010110101011101: color_data = Z;
		19'b0010010110101011110: color_data = Z;
		19'b0010010110101011111: color_data = Z;
		19'b0010010110101100000: color_data = Z;
		19'b0010010110101100001: color_data = Z;
		19'b0010010110101100010: color_data = Z;
		19'b0010010110101100011: color_data = Z;
		19'b0010010110101100100: color_data = Z;
		19'b0010010110101100101: color_data = Z;
		19'b0010010110101100110: color_data = Z;
		19'b0010010110101100111: color_data = Z;
		19'b0010010110101101000: color_data = Z;
		19'b0010010110101101001: color_data = Z;
		19'b0010010110101101010: color_data = Z;
		19'b0010010110101101011: color_data = Z;
		19'b0010010110101101100: color_data = Z;
		19'b0010010110101101101: color_data = Z;
		19'b0010010110101101110: color_data = Z;
		19'b0010010110101101111: color_data = Z;
		19'b0010010110101110000: color_data = Z;
		19'b0010010110101110001: color_data = Z;
		19'b0010010110101110010: color_data = Z;
		19'b0010010110101110011: color_data = Z;
		19'b0010010110101110100: color_data = Z;
		19'b0010010110101110101: color_data = Z;
		19'b0010010110101110110: color_data = Z;
		19'b0010010110101110111: color_data = Z;
		19'b0010010110101111000: color_data = Z;
		19'b0010010110101111001: color_data = Z;
		19'b0010010110101111010: color_data = Z;
		19'b0010010110101111011: color_data = Z;
		19'b0010010110101111100: color_data = Z;
		19'b0010010110101111101: color_data = Z;
		19'b0010010110101111110: color_data = Z;
		19'b0010010110101111111: color_data = Z;
		19'b0010010110110000000: color_data = Z;
		19'b0010010110110000001: color_data = Z;
		19'b0010010110110000010: color_data = Z;
		19'b0010010110110000011: color_data = Z;
		19'b0010010110110000100: color_data = Z;
		19'b0010010110110000101: color_data = Z;
		19'b0010010110110000110: color_data = Z;
		19'b0010010110110000111: color_data = Z;
		19'b0010010110110001000: color_data = Z;
		19'b0010010110110001001: color_data = Z;
		19'b0010010110110001010: color_data = Z;
		19'b0010010110110001011: color_data = Z;
		19'b0010010110110001100: color_data = Z;
		19'b0010010110110001101: color_data = Z;
		19'b0010010110110001110: color_data = Z;
		19'b0010010110110001111: color_data = Z;
		19'b0010010110110010000: color_data = Z;
		19'b0010010110110010001: color_data = Z;
		19'b0010010110110010010: color_data = Z;
		19'b0010010110110010011: color_data = Z;
		19'b0010010110110010100: color_data = Z;
		19'b0010010110110010101: color_data = Z;
		19'b0010010110110010110: color_data = Z;
		19'b0010010110110010111: color_data = Z;
		19'b0010010110110011000: color_data = Z;
		19'b0010010110110011001: color_data = Z;
		19'b0010010110110011010: color_data = Z;
		19'b0010010110110011011: color_data = Z;
		19'b0010010110110011100: color_data = Z;
		19'b0010010110110011101: color_data = Z;
		19'b0010010110110011110: color_data = Z;
		19'b0010010110110011111: color_data = Z;
		19'b0010010110110100000: color_data = Z;
		19'b0010010110110100001: color_data = Z;
		19'b0010010110110100010: color_data = Z;
		19'b0010010110110100011: color_data = Z;
		19'b0010010110110100100: color_data = Z;
		19'b0010010110110100101: color_data = Z;
		19'b0010010110110100110: color_data = Z;
		19'b0010010110110100111: color_data = Z;
		19'b0010010110110101000: color_data = Z;
		19'b0010010110110101001: color_data = Z;
		19'b0010010110110101010: color_data = Z;
		19'b0010010110110101011: color_data = Z;
		19'b0010010110110101100: color_data = Z;
		19'b0010010110110110001: color_data = Z;
		19'b0010010110110110010: color_data = Z;
		19'b0010010110110110100: color_data = Z;
		19'b0010010110110110101: color_data = Z;
		19'b0010010110110110110: color_data = Z;
		19'b0010010110110110111: color_data = Z;
		19'b0010010110110111011: color_data = Z;
		19'b0010010110110111100: color_data = Z;
		19'b0010010110110111101: color_data = Z;
		19'b0010010110110111110: color_data = Z;
		19'b0010010110110111111: color_data = Z;
		19'b0010010110111000000: color_data = Z;
		19'b0010010110111000001: color_data = Z;
		19'b0010010110111000010: color_data = Z;
		19'b0010010110111000011: color_data = Z;
		19'b0010010110111000100: color_data = Z;
		19'b0010010110111000101: color_data = Z;
		19'b0010010110111000110: color_data = Z;
		19'b0010010110111000111: color_data = Z;
		19'b0010010110111001000: color_data = Z;
		19'b0010011000011001001: color_data = Z;
		19'b0010011000011001010: color_data = Z;
		19'b0010011000011001011: color_data = Z;
		19'b0010011000011001100: color_data = Z;
		19'b0010011000011001101: color_data = Z;
		19'b0010011000011001110: color_data = Z;
		19'b0010011000011001111: color_data = Z;
		19'b0010011000011010000: color_data = Z;
		19'b0010011000011010001: color_data = Z;
		19'b0010011000011010010: color_data = Z;
		19'b0010011000011010011: color_data = Z;
		19'b0010011000011010100: color_data = Z;
		19'b0010011000011010101: color_data = Z;
		19'b0010011000011010110: color_data = Z;
		19'b0010011000011010111: color_data = Z;
		19'b0010011000011011000: color_data = Z;
		19'b0010011000011011001: color_data = Z;
		19'b0010011000011011010: color_data = Z;
		19'b0010011000011011011: color_data = Z;
		19'b0010011000011011100: color_data = Z;
		19'b0010011000011011101: color_data = Z;
		19'b0010011000011011110: color_data = Z;
		19'b0010011000011011111: color_data = Z;
		19'b0010011000011100000: color_data = Z;
		19'b0010011000011100001: color_data = Z;
		19'b0010011000011100010: color_data = Z;
		19'b0010011000011100011: color_data = Z;
		19'b0010011000011100100: color_data = Z;
		19'b0010011000011100101: color_data = Z;
		19'b0010011000011100110: color_data = Z;
		19'b0010011000011100111: color_data = Z;
		19'b0010011000011101000: color_data = Z;
		19'b0010011000011101001: color_data = Z;
		19'b0010011000011101010: color_data = Z;
		19'b0010011000011101011: color_data = Z;
		19'b0010011000011101100: color_data = Z;
		19'b0010011000011101101: color_data = Z;
		19'b0010011000011101110: color_data = Z;
		19'b0010011000011101111: color_data = Z;
		19'b0010011000011110000: color_data = Z;
		19'b0010011000011110001: color_data = Z;
		19'b0010011000011110010: color_data = Z;
		19'b0010011000011110011: color_data = Z;
		19'b0010011000011110100: color_data = Z;
		19'b0010011000011110101: color_data = Z;
		19'b0010011000011110110: color_data = Z;
		19'b0010011000011110111: color_data = Z;
		19'b0010011000011111000: color_data = Z;
		19'b0010011000011111001: color_data = Z;
		19'b0010011000011111010: color_data = Z;
		19'b0010011000011111011: color_data = Z;
		19'b0010011000011111100: color_data = Z;
		19'b0010011000011111101: color_data = Z;
		19'b0010011000011111110: color_data = Z;
		19'b0010011000011111111: color_data = Z;
		19'b0010011000100000000: color_data = Z;
		19'b0010011000100000001: color_data = Z;
		19'b0010011000100000010: color_data = Z;
		19'b0010011000100000011: color_data = Z;
		19'b0010011000100000100: color_data = Z;
		19'b0010011000100000101: color_data = Z;
		19'b0010011000100000110: color_data = Z;
		19'b0010011000100000111: color_data = Z;
		19'b0010011000100001000: color_data = Z;
		19'b0010011000100001001: color_data = Z;
		19'b0010011000100001010: color_data = Z;
		19'b0010011000100001011: color_data = Z;
		19'b0010011000100001100: color_data = Z;
		19'b0010011000100001101: color_data = Z;
		19'b0010011000100001110: color_data = Z;
		19'b0010011000100001111: color_data = Z;
		19'b0010011000100010000: color_data = Z;
		19'b0010011000100010001: color_data = Z;
		19'b0010011000100010010: color_data = Z;
		19'b0010011000100010011: color_data = Z;
		19'b0010011000100010100: color_data = Z;
		19'b0010011000100010101: color_data = Z;
		19'b0010011000100010110: color_data = Z;
		19'b0010011000100010111: color_data = Z;
		19'b0010011000100011000: color_data = Z;
		19'b0010011000100011001: color_data = Z;
		19'b0010011000100011010: color_data = Z;
		19'b0010011000100011011: color_data = Z;
		19'b0010011000100011100: color_data = Z;
		19'b0010011000100011101: color_data = Z;
		19'b0010011000100011110: color_data = Z;
		19'b0010011000100011111: color_data = Z;
		19'b0010011000100100000: color_data = Z;
		19'b0010011000100100001: color_data = Z;
		19'b0010011000100100010: color_data = Z;
		19'b0010011000100100011: color_data = Z;
		19'b0010011000100100100: color_data = Z;
		19'b0010011000100100101: color_data = Z;
		19'b0010011000100100110: color_data = Z;
		19'b0010011000100100111: color_data = Z;
		19'b0010011000100101000: color_data = Z;
		19'b0010011000100101001: color_data = Z;
		19'b0010011000100101010: color_data = Z;
		19'b0010011000100101011: color_data = Z;
		19'b0010011000100101100: color_data = Z;
		19'b0010011000100101101: color_data = Z;
		19'b0010011000100101110: color_data = Z;
		19'b0010011000100101111: color_data = Z;
		19'b0010011000100110000: color_data = Z;
		19'b0010011000100110001: color_data = Z;
		19'b0010011000100110010: color_data = Z;
		19'b0010011000100110011: color_data = Z;
		19'b0010011000100110100: color_data = Z;
		19'b0010011000100110101: color_data = Z;
		19'b0010011000100110110: color_data = Z;
		19'b0010011000100110111: color_data = Z;
		19'b0010011000100111000: color_data = Z;
		19'b0010011000100111001: color_data = Z;
		19'b0010011000100111010: color_data = Z;
		19'b0010011000100111011: color_data = Z;
		19'b0010011000100111100: color_data = Z;
		19'b0010011000100111101: color_data = Z;
		19'b0010011000100111110: color_data = Z;
		19'b0010011000100111111: color_data = Z;
		19'b0010011000101000000: color_data = Z;
		19'b0010011000101000001: color_data = Z;
		19'b0010011000101000010: color_data = Z;
		19'b0010011000101000011: color_data = Z;
		19'b0010011000101000100: color_data = Z;
		19'b0010011000101000101: color_data = Z;
		19'b0010011000101000110: color_data = Z;
		19'b0010011000101000111: color_data = Z;
		19'b0010011000101001000: color_data = Z;
		19'b0010011000101001001: color_data = Z;
		19'b0010011000101001010: color_data = Z;
		19'b0010011000101001011: color_data = Z;
		19'b0010011000101001100: color_data = Z;
		19'b0010011000101001101: color_data = Z;
		19'b0010011000101001110: color_data = Z;
		19'b0010011000101001111: color_data = Z;
		19'b0010011000101010000: color_data = Z;
		19'b0010011000101010001: color_data = Z;
		19'b0010011000101010010: color_data = Z;
		19'b0010011000101010011: color_data = Z;
		19'b0010011000101010100: color_data = Z;
		19'b0010011000101010101: color_data = Z;
		19'b0010011000101010110: color_data = Z;
		19'b0010011000101010111: color_data = Z;
		19'b0010011000101011000: color_data = Z;
		19'b0010011000101011001: color_data = Z;
		19'b0010011000101011010: color_data = Z;
		19'b0010011000101011011: color_data = Z;
		19'b0010011000101011100: color_data = Z;
		19'b0010011000101011101: color_data = Z;
		19'b0010011000101011110: color_data = Z;
		19'b0010011000101011111: color_data = Z;
		19'b0010011000101100000: color_data = Z;
		19'b0010011000101100001: color_data = Z;
		19'b0010011000101100010: color_data = Z;
		19'b0010011000101100011: color_data = Z;
		19'b0010011000101100100: color_data = Z;
		19'b0010011000101100101: color_data = Z;
		19'b0010011000101100110: color_data = Z;
		19'b0010011000101100111: color_data = Z;
		19'b0010011000101101000: color_data = Z;
		19'b0010011000101101001: color_data = Z;
		19'b0010011000101101010: color_data = Z;
		19'b0010011000101101011: color_data = Z;
		19'b0010011000101101100: color_data = Z;
		19'b0010011000101101101: color_data = Z;
		19'b0010011000101101110: color_data = Z;
		19'b0010011000101101111: color_data = Z;
		19'b0010011000101110000: color_data = Z;
		19'b0010011000101110001: color_data = Z;
		19'b0010011000101110010: color_data = Z;
		19'b0010011000101110011: color_data = Z;
		19'b0010011000101110100: color_data = Z;
		19'b0010011000101110101: color_data = Z;
		19'b0010011000101110110: color_data = Z;
		19'b0010011000101110111: color_data = Z;
		19'b0010011000101111000: color_data = Z;
		19'b0010011000101111001: color_data = Z;
		19'b0010011000101111010: color_data = Z;
		19'b0010011000101111011: color_data = Z;
		19'b0010011000101111100: color_data = Z;
		19'b0010011000101111101: color_data = Z;
		19'b0010011000101111110: color_data = Z;
		19'b0010011000101111111: color_data = Z;
		19'b0010011000110000000: color_data = Z;
		19'b0010011000110000001: color_data = Z;
		19'b0010011000110000010: color_data = Z;
		19'b0010011000110000011: color_data = Z;
		19'b0010011000110000100: color_data = Z;
		19'b0010011000110000101: color_data = Z;
		19'b0010011000110000110: color_data = Z;
		19'b0010011000110000111: color_data = Z;
		19'b0010011000110001000: color_data = Z;
		19'b0010011000110001001: color_data = Z;
		19'b0010011000110001010: color_data = Z;
		19'b0010011000110001011: color_data = Z;
		19'b0010011000110001100: color_data = Z;
		19'b0010011000110001101: color_data = Z;
		19'b0010011000110001110: color_data = Z;
		19'b0010011000110001111: color_data = Z;
		19'b0010011000110010000: color_data = Z;
		19'b0010011000110010001: color_data = Z;
		19'b0010011000110010010: color_data = Z;
		19'b0010011000110010011: color_data = Z;
		19'b0010011000110010100: color_data = Z;
		19'b0010011000110010101: color_data = Z;
		19'b0010011000110010110: color_data = Z;
		19'b0010011000110010111: color_data = Z;
		19'b0010011000110011000: color_data = Z;
		19'b0010011000110011001: color_data = Z;
		19'b0010011000110011010: color_data = Z;
		19'b0010011000110011011: color_data = Z;
		19'b0010011000110011100: color_data = Z;
		19'b0010011000110011101: color_data = Z;
		19'b0010011000110011110: color_data = Z;
		19'b0010011000110011111: color_data = Z;
		19'b0010011000110100000: color_data = Z;
		19'b0010011000110100001: color_data = Z;
		19'b0010011000110100010: color_data = Z;
		19'b0010011000110100011: color_data = Z;
		19'b0010011000110100100: color_data = Z;
		19'b0010011000110100101: color_data = Z;
		19'b0010011000110100110: color_data = Z;
		19'b0010011000110100111: color_data = Z;
		19'b0010011000110101000: color_data = Z;
		19'b0010011000110101001: color_data = Z;
		19'b0010011000110101010: color_data = Z;
		19'b0010011000110101011: color_data = Z;
		19'b0010011000110101100: color_data = Z;
		19'b0010011000110101101: color_data = Z;
		19'b0010011000110110010: color_data = Z;
		19'b0010011000110110011: color_data = Z;
		19'b0010011000110110101: color_data = Z;
		19'b0010011000110110110: color_data = Z;
		19'b0010011000110110111: color_data = Z;
		19'b0010011000110111000: color_data = Z;
		19'b0010011000110111011: color_data = Z;
		19'b0010011000110111100: color_data = Z;
		19'b0010011000110111101: color_data = Z;
		19'b0010011000110111110: color_data = Z;
		19'b0010011000110111111: color_data = Z;
		19'b0010011000111000000: color_data = Z;
		19'b0010011000111000001: color_data = Z;
		19'b0010011000111000010: color_data = Z;
		19'b0010011000111000011: color_data = Z;
		19'b0010011000111000100: color_data = Z;
		19'b0010011000111000101: color_data = Z;
		19'b0010011000111000110: color_data = Z;
		19'b0010011000111000111: color_data = Z;
		19'b0010011000111001000: color_data = Z;
		19'b0010011000111001001: color_data = Z;
		19'b0010011010011001001: color_data = Z;
		19'b0010011010011001010: color_data = Z;
		19'b0010011010011001011: color_data = Z;
		19'b0010011010011001100: color_data = Z;
		19'b0010011010011001101: color_data = Z;
		19'b0010011010011001110: color_data = Z;
		19'b0010011010011001111: color_data = Z;
		19'b0010011010011010000: color_data = Z;
		19'b0010011010011010001: color_data = Z;
		19'b0010011010011010010: color_data = Z;
		19'b0010011010011010011: color_data = Z;
		19'b0010011010011010100: color_data = Z;
		19'b0010011010011010101: color_data = Z;
		19'b0010011010011010110: color_data = Z;
		19'b0010011010011010111: color_data = Z;
		19'b0010011010011011000: color_data = Z;
		19'b0010011010011011001: color_data = Z;
		19'b0010011010011011010: color_data = Z;
		19'b0010011010011011011: color_data = Z;
		19'b0010011010011011100: color_data = Z;
		19'b0010011010011011101: color_data = Z;
		19'b0010011010011011110: color_data = Z;
		19'b0010011010011011111: color_data = Z;
		19'b0010011010011100000: color_data = Z;
		19'b0010011010011100001: color_data = Z;
		19'b0010011010011100010: color_data = Z;
		19'b0010011010011100011: color_data = Z;
		19'b0010011010011100100: color_data = Z;
		19'b0010011010011100101: color_data = Z;
		19'b0010011010011100110: color_data = Z;
		19'b0010011010011100111: color_data = Z;
		19'b0010011010011101000: color_data = Z;
		19'b0010011010011101001: color_data = Z;
		19'b0010011010011101010: color_data = Z;
		19'b0010011010011101011: color_data = Z;
		19'b0010011010011101100: color_data = Z;
		19'b0010011010011101101: color_data = Z;
		19'b0010011010011101110: color_data = Z;
		19'b0010011010011101111: color_data = Z;
		19'b0010011010011110000: color_data = Z;
		19'b0010011010011110001: color_data = Z;
		19'b0010011010011110010: color_data = Z;
		19'b0010011010011110011: color_data = Z;
		19'b0010011010011110100: color_data = Z;
		19'b0010011010011110101: color_data = Z;
		19'b0010011010011110110: color_data = Z;
		19'b0010011010011110111: color_data = Z;
		19'b0010011010011111000: color_data = Z;
		19'b0010011010011111001: color_data = Z;
		19'b0010011010011111010: color_data = Z;
		19'b0010011010011111011: color_data = Z;
		19'b0010011010011111100: color_data = Z;
		19'b0010011010011111101: color_data = Z;
		19'b0010011010011111110: color_data = Z;
		19'b0010011010011111111: color_data = Z;
		19'b0010011010100000000: color_data = Z;
		19'b0010011010100000001: color_data = Z;
		19'b0010011010100000010: color_data = Z;
		19'b0010011010100000011: color_data = Z;
		19'b0010011010100000100: color_data = Z;
		19'b0010011010100000101: color_data = Z;
		19'b0010011010100000110: color_data = Z;
		19'b0010011010100000111: color_data = Z;
		19'b0010011010100001000: color_data = Z;
		19'b0010011010100001001: color_data = Z;
		19'b0010011010100001010: color_data = Z;
		19'b0010011010100001011: color_data = Z;
		19'b0010011010100001100: color_data = Z;
		19'b0010011010100001101: color_data = Z;
		19'b0010011010100001110: color_data = Z;
		19'b0010011010100001111: color_data = Z;
		19'b0010011010100010000: color_data = Z;
		19'b0010011010100010001: color_data = Z;
		19'b0010011010100010010: color_data = Z;
		19'b0010011010100010011: color_data = Z;
		19'b0010011010100010100: color_data = Z;
		19'b0010011010100010101: color_data = Z;
		19'b0010011010100010110: color_data = Z;
		19'b0010011010100010111: color_data = Z;
		19'b0010011010100011000: color_data = Z;
		19'b0010011010100011001: color_data = Z;
		19'b0010011010100011010: color_data = Z;
		19'b0010011010100011011: color_data = Z;
		19'b0010011010100011100: color_data = Z;
		19'b0010011010100011101: color_data = Z;
		19'b0010011010100011110: color_data = Z;
		19'b0010011010100011111: color_data = Z;
		19'b0010011010100100000: color_data = Z;
		19'b0010011010100100001: color_data = Z;
		19'b0010011010100100010: color_data = Z;
		19'b0010011010100100011: color_data = Z;
		19'b0010011010100100100: color_data = Z;
		19'b0010011010100100101: color_data = Z;
		19'b0010011010100100110: color_data = Z;
		19'b0010011010100100111: color_data = Z;
		19'b0010011010100101000: color_data = Z;
		19'b0010011010100101001: color_data = Z;
		19'b0010011010100101010: color_data = Z;
		19'b0010011010100101011: color_data = Z;
		19'b0010011010100101100: color_data = Z;
		19'b0010011010100101101: color_data = Z;
		19'b0010011010100101110: color_data = Z;
		19'b0010011010100101111: color_data = Z;
		19'b0010011010100110000: color_data = Z;
		19'b0010011010100110001: color_data = Z;
		19'b0010011010100110010: color_data = Z;
		19'b0010011010100110011: color_data = Z;
		19'b0010011010100110100: color_data = Z;
		19'b0010011010100110101: color_data = Z;
		19'b0010011010100110110: color_data = Z;
		19'b0010011010100110111: color_data = Z;
		19'b0010011010100111000: color_data = Z;
		19'b0010011010100111001: color_data = Z;
		19'b0010011010100111010: color_data = Z;
		19'b0010011010100111011: color_data = Z;
		19'b0010011010100111100: color_data = Z;
		19'b0010011010100111101: color_data = Z;
		19'b0010011010100111110: color_data = Z;
		19'b0010011010100111111: color_data = Z;
		19'b0010011010101000000: color_data = Z;
		19'b0010011010101000001: color_data = Z;
		19'b0010011010101000010: color_data = Z;
		19'b0010011010101000011: color_data = Z;
		19'b0010011010101000100: color_data = Z;
		19'b0010011010101000101: color_data = Z;
		19'b0010011010101000110: color_data = Z;
		19'b0010011010101000111: color_data = Z;
		19'b0010011010101001000: color_data = Z;
		19'b0010011010101001001: color_data = Z;
		19'b0010011010101001010: color_data = Z;
		19'b0010011010101001011: color_data = Z;
		19'b0010011010101001100: color_data = Z;
		19'b0010011010101001101: color_data = Z;
		19'b0010011010101001110: color_data = Z;
		19'b0010011010101001111: color_data = Z;
		19'b0010011010101010000: color_data = Z;
		19'b0010011010101010001: color_data = Z;
		19'b0010011010101010010: color_data = Z;
		19'b0010011010101010011: color_data = Z;
		19'b0010011010101010100: color_data = Z;
		19'b0010011010101010101: color_data = Z;
		19'b0010011010101010110: color_data = Z;
		19'b0010011010101010111: color_data = Z;
		19'b0010011010101011000: color_data = Z;
		19'b0010011010101011001: color_data = Z;
		19'b0010011010101011010: color_data = Z;
		19'b0010011010101011011: color_data = Z;
		19'b0010011010101011100: color_data = Z;
		19'b0010011010101011101: color_data = Z;
		19'b0010011010101011110: color_data = Z;
		19'b0010011010101011111: color_data = Z;
		19'b0010011010101100000: color_data = Z;
		19'b0010011010101100001: color_data = Z;
		19'b0010011010101100010: color_data = Z;
		19'b0010011010101100011: color_data = Z;
		19'b0010011010101100100: color_data = Z;
		19'b0010011010101100101: color_data = Z;
		19'b0010011010101100110: color_data = Z;
		19'b0010011010101100111: color_data = Z;
		19'b0010011010101101000: color_data = Z;
		19'b0010011010101101001: color_data = Z;
		19'b0010011010101101010: color_data = Z;
		19'b0010011010101101011: color_data = Z;
		19'b0010011010101101100: color_data = Z;
		19'b0010011010101101101: color_data = Z;
		19'b0010011010101101110: color_data = Z;
		19'b0010011010101101111: color_data = Z;
		19'b0010011010101110000: color_data = Z;
		19'b0010011010101110001: color_data = Z;
		19'b0010011010101110010: color_data = Z;
		19'b0010011010101110011: color_data = Z;
		19'b0010011010101110100: color_data = Z;
		19'b0010011010101110101: color_data = Z;
		19'b0010011010101110110: color_data = Z;
		19'b0010011010101110111: color_data = Z;
		19'b0010011010101111000: color_data = Z;
		19'b0010011010101111001: color_data = Z;
		19'b0010011010101111010: color_data = Z;
		19'b0010011010101111011: color_data = Z;
		19'b0010011010101111100: color_data = Z;
		19'b0010011010101111101: color_data = Z;
		19'b0010011010101111110: color_data = Z;
		19'b0010011010101111111: color_data = Z;
		19'b0010011010110000000: color_data = Z;
		19'b0010011010110000001: color_data = Z;
		19'b0010011010110000010: color_data = Z;
		19'b0010011010110000011: color_data = Z;
		19'b0010011010110000100: color_data = Z;
		19'b0010011010110000101: color_data = Z;
		19'b0010011010110000110: color_data = Z;
		19'b0010011010110000111: color_data = Z;
		19'b0010011010110001000: color_data = Z;
		19'b0010011010110001001: color_data = Z;
		19'b0010011010110001010: color_data = Z;
		19'b0010011010110001011: color_data = Z;
		19'b0010011010110001100: color_data = Z;
		19'b0010011010110001101: color_data = Z;
		19'b0010011010110001110: color_data = Z;
		19'b0010011010110001111: color_data = Z;
		19'b0010011010110010000: color_data = Z;
		19'b0010011010110010001: color_data = Z;
		19'b0010011010110010010: color_data = Z;
		19'b0010011010110010011: color_data = Z;
		19'b0010011010110010100: color_data = Z;
		19'b0010011010110010101: color_data = Z;
		19'b0010011010110010110: color_data = Z;
		19'b0010011010110010111: color_data = Z;
		19'b0010011010110011000: color_data = Z;
		19'b0010011010110011001: color_data = Z;
		19'b0010011010110011010: color_data = Z;
		19'b0010011010110011011: color_data = Z;
		19'b0010011010110011100: color_data = Z;
		19'b0010011010110011101: color_data = Z;
		19'b0010011010110011110: color_data = Z;
		19'b0010011010110011111: color_data = Z;
		19'b0010011010110100000: color_data = Z;
		19'b0010011010110100001: color_data = Z;
		19'b0010011010110100010: color_data = Z;
		19'b0010011010110100011: color_data = Z;
		19'b0010011010110100100: color_data = Z;
		19'b0010011010110100101: color_data = Z;
		19'b0010011010110100110: color_data = Z;
		19'b0010011010110100111: color_data = Z;
		19'b0010011010110101000: color_data = Z;
		19'b0010011010110101001: color_data = Z;
		19'b0010011010110101010: color_data = Z;
		19'b0010011010110101011: color_data = Z;
		19'b0010011010110101100: color_data = Z;
		19'b0010011010110101101: color_data = Z;
		19'b0010011010110110011: color_data = Z;
		19'b0010011010110110100: color_data = Z;
		19'b0010011010110110101: color_data = Z;
		19'b0010011010110110110: color_data = Z;
		19'b0010011010110110111: color_data = Z;
		19'b0010011010110111000: color_data = Z;
		19'b0010011010110111100: color_data = Z;
		19'b0010011010110111101: color_data = Z;
		19'b0010011010110111110: color_data = Z;
		19'b0010011010110111111: color_data = Z;
		19'b0010011010111000000: color_data = Z;
		19'b0010011010111000001: color_data = Z;
		19'b0010011010111000010: color_data = Z;
		19'b0010011010111000011: color_data = Z;
		19'b0010011010111000100: color_data = Z;
		19'b0010011010111000101: color_data = Z;
		19'b0010011010111000110: color_data = Z;
		19'b0010011010111000111: color_data = Z;
		19'b0010011010111001000: color_data = Z;
		19'b0010011010111001001: color_data = Z;
		19'b0010011100011001010: color_data = Z;
		19'b0010011100011001011: color_data = Z;
		19'b0010011100011001100: color_data = Z;
		19'b0010011100011001101: color_data = Z;
		19'b0010011100011001110: color_data = Z;
		19'b0010011100011001111: color_data = Z;
		19'b0010011100011010000: color_data = Z;
		19'b0010011100011010001: color_data = Z;
		19'b0010011100011010010: color_data = Z;
		19'b0010011100011010011: color_data = Z;
		19'b0010011100011010100: color_data = Z;
		19'b0010011100011010101: color_data = Z;
		19'b0010011100011010110: color_data = Z;
		19'b0010011100011010111: color_data = Z;
		19'b0010011100011011000: color_data = Z;
		19'b0010011100011011001: color_data = Z;
		19'b0010011100011011010: color_data = Z;
		19'b0010011100011011011: color_data = Z;
		19'b0010011100011011100: color_data = Z;
		19'b0010011100011011101: color_data = Z;
		19'b0010011100011011110: color_data = Z;
		19'b0010011100011011111: color_data = Z;
		19'b0010011100011100000: color_data = Z;
		19'b0010011100011100001: color_data = Z;
		19'b0010011100011100010: color_data = Z;
		19'b0010011100011100011: color_data = Z;
		19'b0010011100011100100: color_data = Z;
		19'b0010011100011100101: color_data = Z;
		19'b0010011100011100110: color_data = Z;
		19'b0010011100011100111: color_data = Z;
		19'b0010011100011101000: color_data = Z;
		19'b0010011100011101001: color_data = Z;
		19'b0010011100011101010: color_data = Z;
		19'b0010011100011101011: color_data = Z;
		19'b0010011100011101100: color_data = Z;
		19'b0010011100011101101: color_data = Z;
		19'b0010011100011101110: color_data = Z;
		19'b0010011100011101111: color_data = Z;
		19'b0010011100011110000: color_data = Z;
		19'b0010011100011110001: color_data = Z;
		19'b0010011100011110010: color_data = Z;
		19'b0010011100011110011: color_data = Z;
		19'b0010011100011110100: color_data = Z;
		19'b0010011100011110101: color_data = Z;
		19'b0010011100011110110: color_data = Z;
		19'b0010011100011110111: color_data = Z;
		19'b0010011100011111000: color_data = Z;
		19'b0010011100011111001: color_data = Z;
		19'b0010011100011111010: color_data = Z;
		19'b0010011100011111011: color_data = Z;
		19'b0010011100011111100: color_data = Z;
		19'b0010011100011111101: color_data = Z;
		19'b0010011100011111110: color_data = Z;
		19'b0010011100011111111: color_data = Z;
		19'b0010011100100000000: color_data = Z;
		19'b0010011100100000001: color_data = Z;
		19'b0010011100100000010: color_data = Z;
		19'b0010011100100000011: color_data = Z;
		19'b0010011100100000100: color_data = Z;
		19'b0010011100100000101: color_data = Z;
		19'b0010011100100000110: color_data = Z;
		19'b0010011100100000111: color_data = Z;
		19'b0010011100100001000: color_data = Z;
		19'b0010011100100001001: color_data = Z;
		19'b0010011100100001010: color_data = Z;
		19'b0010011100100001011: color_data = Z;
		19'b0010011100100001100: color_data = Z;
		19'b0010011100100001101: color_data = Z;
		19'b0010011100100001110: color_data = Z;
		19'b0010011100100001111: color_data = Z;
		19'b0010011100100010000: color_data = Z;
		19'b0010011100100010001: color_data = Z;
		19'b0010011100100010010: color_data = Z;
		19'b0010011100100010011: color_data = Z;
		19'b0010011100100010100: color_data = Z;
		19'b0010011100100010101: color_data = Z;
		19'b0010011100100010110: color_data = Z;
		19'b0010011100100010111: color_data = Z;
		19'b0010011100100011000: color_data = Z;
		19'b0010011100100011001: color_data = Z;
		19'b0010011100100011010: color_data = Z;
		19'b0010011100100011011: color_data = Z;
		19'b0010011100100011100: color_data = Z;
		19'b0010011100100011101: color_data = Z;
		19'b0010011100100011110: color_data = Z;
		19'b0010011100100011111: color_data = Z;
		19'b0010011100100100000: color_data = Z;
		19'b0010011100100100001: color_data = Z;
		19'b0010011100100100010: color_data = Z;
		19'b0010011100100100011: color_data = Z;
		19'b0010011100100100100: color_data = Z;
		19'b0010011100100100101: color_data = Z;
		19'b0010011100100100110: color_data = Z;
		19'b0010011100100100111: color_data = Z;
		19'b0010011100100101000: color_data = Z;
		19'b0010011100100101001: color_data = Z;
		19'b0010011100100101010: color_data = Z;
		19'b0010011100100101011: color_data = Z;
		19'b0010011100100101100: color_data = Z;
		19'b0010011100100101101: color_data = Z;
		19'b0010011100100101110: color_data = Z;
		19'b0010011100100101111: color_data = Z;
		19'b0010011100100110000: color_data = Z;
		19'b0010011100100110001: color_data = Z;
		19'b0010011100100110010: color_data = Z;
		19'b0010011100100110011: color_data = Z;
		19'b0010011100100110100: color_data = Z;
		19'b0010011100100110101: color_data = Z;
		19'b0010011100100110110: color_data = Z;
		19'b0010011100100110111: color_data = Z;
		19'b0010011100100111000: color_data = Z;
		19'b0010011100100111001: color_data = Z;
		19'b0010011100100111010: color_data = Z;
		19'b0010011100100111011: color_data = Z;
		19'b0010011100100111100: color_data = Z;
		19'b0010011100100111101: color_data = Z;
		19'b0010011100100111110: color_data = Z;
		19'b0010011100100111111: color_data = Z;
		19'b0010011100101000000: color_data = Z;
		19'b0010011100101000001: color_data = Z;
		19'b0010011100101000010: color_data = Z;
		19'b0010011100101000011: color_data = Z;
		19'b0010011100101000100: color_data = Z;
		19'b0010011100101000101: color_data = Z;
		19'b0010011100101000110: color_data = Z;
		19'b0010011100101000111: color_data = Z;
		19'b0010011100101001000: color_data = Z;
		19'b0010011100101001001: color_data = Z;
		19'b0010011100101001010: color_data = Z;
		19'b0010011100101001011: color_data = Z;
		19'b0010011100101001100: color_data = Z;
		19'b0010011100101001101: color_data = Z;
		19'b0010011100101001110: color_data = Z;
		19'b0010011100101001111: color_data = Z;
		19'b0010011100101010000: color_data = Z;
		19'b0010011100101010001: color_data = Z;
		19'b0010011100101010010: color_data = Z;
		19'b0010011100101010011: color_data = Z;
		19'b0010011100101010100: color_data = Z;
		19'b0010011100101010101: color_data = Z;
		19'b0010011100101010110: color_data = Z;
		19'b0010011100101010111: color_data = Z;
		19'b0010011100101011000: color_data = Z;
		19'b0010011100101011001: color_data = Z;
		19'b0010011100101011010: color_data = Z;
		19'b0010011100101011011: color_data = Z;
		19'b0010011100101011100: color_data = Z;
		19'b0010011100101011101: color_data = Z;
		19'b0010011100101011110: color_data = Z;
		19'b0010011100101011111: color_data = Z;
		19'b0010011100101100000: color_data = Z;
		19'b0010011100101100001: color_data = Z;
		19'b0010011100101100010: color_data = Z;
		19'b0010011100101100011: color_data = Z;
		19'b0010011100101100100: color_data = Z;
		19'b0010011100101100101: color_data = Z;
		19'b0010011100101100110: color_data = Z;
		19'b0010011100101100111: color_data = Z;
		19'b0010011100101101000: color_data = Z;
		19'b0010011100101101001: color_data = Z;
		19'b0010011100101101010: color_data = Z;
		19'b0010011100101101011: color_data = Z;
		19'b0010011100101101100: color_data = Z;
		19'b0010011100101101101: color_data = Z;
		19'b0010011100101101110: color_data = Z;
		19'b0010011100101101111: color_data = Z;
		19'b0010011100101110000: color_data = Z;
		19'b0010011100101110001: color_data = Z;
		19'b0010011100101110010: color_data = Z;
		19'b0010011100101110011: color_data = Z;
		19'b0010011100101110100: color_data = Z;
		19'b0010011100101110101: color_data = Z;
		19'b0010011100101110110: color_data = Z;
		19'b0010011100101110111: color_data = Z;
		19'b0010011100101111000: color_data = Z;
		19'b0010011100101111001: color_data = Z;
		19'b0010011100101111010: color_data = Z;
		19'b0010011100101111011: color_data = Z;
		19'b0010011100101111100: color_data = Z;
		19'b0010011100101111101: color_data = Z;
		19'b0010011100101111110: color_data = Z;
		19'b0010011100101111111: color_data = Z;
		19'b0010011100110000000: color_data = Z;
		19'b0010011100110000001: color_data = Z;
		19'b0010011100110000010: color_data = Z;
		19'b0010011100110000011: color_data = Z;
		19'b0010011100110000100: color_data = Z;
		19'b0010011100110000101: color_data = Z;
		19'b0010011100110000110: color_data = Z;
		19'b0010011100110000111: color_data = Z;
		19'b0010011100110001000: color_data = Z;
		19'b0010011100110001001: color_data = Z;
		19'b0010011100110001010: color_data = Z;
		19'b0010011100110001011: color_data = Z;
		19'b0010011100110001100: color_data = Z;
		19'b0010011100110001101: color_data = Z;
		19'b0010011100110001110: color_data = Z;
		19'b0010011100110001111: color_data = Z;
		19'b0010011100110010000: color_data = Z;
		19'b0010011100110010001: color_data = Z;
		19'b0010011100110010010: color_data = Z;
		19'b0010011100110010011: color_data = Z;
		19'b0010011100110010100: color_data = Z;
		19'b0010011100110010101: color_data = Z;
		19'b0010011100110010110: color_data = Z;
		19'b0010011100110010111: color_data = Z;
		19'b0010011100110011000: color_data = Z;
		19'b0010011100110011001: color_data = Z;
		19'b0010011100110011010: color_data = Z;
		19'b0010011100110011011: color_data = Z;
		19'b0010011100110011100: color_data = Z;
		19'b0010011100110011101: color_data = Z;
		19'b0010011100110011110: color_data = Z;
		19'b0010011100110011111: color_data = Z;
		19'b0010011100110100000: color_data = Z;
		19'b0010011100110100001: color_data = Z;
		19'b0010011100110100010: color_data = Z;
		19'b0010011100110100011: color_data = Z;
		19'b0010011100110100100: color_data = Z;
		19'b0010011100110100101: color_data = Z;
		19'b0010011100110100110: color_data = Z;
		19'b0010011100110100111: color_data = Z;
		19'b0010011100110101000: color_data = Z;
		19'b0010011100110101001: color_data = Z;
		19'b0010011100110101010: color_data = Z;
		19'b0010011100110101011: color_data = Z;
		19'b0010011100110101100: color_data = Z;
		19'b0010011100110101101: color_data = Z;
		19'b0010011100110101110: color_data = Z;
		19'b0010011100110110011: color_data = Z;
		19'b0010011100110110100: color_data = Z;
		19'b0010011100110110101: color_data = Z;
		19'b0010011100110110110: color_data = Z;
		19'b0010011100110110111: color_data = Z;
		19'b0010011100110111000: color_data = Z;
		19'b0010011100110111001: color_data = Z;
		19'b0010011100110111101: color_data = Z;
		19'b0010011100110111110: color_data = Z;
		19'b0010011100110111111: color_data = Z;
		19'b0010011100111000000: color_data = Z;
		19'b0010011100111000001: color_data = Z;
		19'b0010011100111000010: color_data = Z;
		19'b0010011100111000011: color_data = Z;
		19'b0010011100111000100: color_data = Z;
		19'b0010011100111000101: color_data = Z;
		19'b0010011100111000110: color_data = Z;
		19'b0010011100111000111: color_data = Z;
		19'b0010011100111001000: color_data = Z;
		19'b0010011100111001001: color_data = Z;
		19'b0010011100111001010: color_data = Z;
		19'b0010011110011001011: color_data = Z;
		19'b0010011110011001100: color_data = Z;
		19'b0010011110011001101: color_data = Z;
		19'b0010011110011001110: color_data = Z;
		19'b0010011110011001111: color_data = Z;
		19'b0010011110011010000: color_data = Z;
		19'b0010011110011010001: color_data = Z;
		19'b0010011110011010010: color_data = Z;
		19'b0010011110011010011: color_data = Z;
		19'b0010011110011010100: color_data = Z;
		19'b0010011110011010101: color_data = Z;
		19'b0010011110011010110: color_data = Z;
		19'b0010011110011010111: color_data = Z;
		19'b0010011110011011000: color_data = Z;
		19'b0010011110011011001: color_data = Z;
		19'b0010011110011011010: color_data = Z;
		19'b0010011110011011011: color_data = Z;
		19'b0010011110011011100: color_data = Z;
		19'b0010011110011011101: color_data = Z;
		19'b0010011110011011110: color_data = Z;
		19'b0010011110011011111: color_data = Z;
		19'b0010011110011100000: color_data = Z;
		19'b0010011110011100001: color_data = Z;
		19'b0010011110011100010: color_data = Z;
		19'b0010011110011100011: color_data = Z;
		19'b0010011110011100100: color_data = Z;
		19'b0010011110011100101: color_data = Z;
		19'b0010011110011100110: color_data = Z;
		19'b0010011110011100111: color_data = Z;
		19'b0010011110011101000: color_data = Z;
		19'b0010011110011101001: color_data = Z;
		19'b0010011110011101010: color_data = Z;
		19'b0010011110011101011: color_data = Z;
		19'b0010011110011101100: color_data = Z;
		19'b0010011110011101101: color_data = Z;
		19'b0010011110011101110: color_data = Z;
		19'b0010011110011101111: color_data = Z;
		19'b0010011110011110000: color_data = Z;
		19'b0010011110011110001: color_data = Z;
		19'b0010011110011110010: color_data = Z;
		19'b0010011110011110011: color_data = Z;
		19'b0010011110011110100: color_data = Z;
		19'b0010011110011110101: color_data = Z;
		19'b0010011110011110110: color_data = Z;
		19'b0010011110011110111: color_data = Z;
		19'b0010011110011111000: color_data = Z;
		19'b0010011110011111001: color_data = Z;
		19'b0010011110011111010: color_data = Z;
		19'b0010011110011111011: color_data = Z;
		19'b0010011110011111100: color_data = Z;
		19'b0010011110011111101: color_data = Z;
		19'b0010011110011111110: color_data = Z;
		19'b0010011110011111111: color_data = Z;
		19'b0010011110100000000: color_data = Z;
		19'b0010011110100000001: color_data = Z;
		19'b0010011110100000010: color_data = Z;
		19'b0010011110100000011: color_data = Z;
		19'b0010011110100000100: color_data = Z;
		19'b0010011110100000101: color_data = Z;
		19'b0010011110100000110: color_data = Z;
		19'b0010011110100000111: color_data = Z;
		19'b0010011110100001000: color_data = Z;
		19'b0010011110100001001: color_data = Z;
		19'b0010011110100001010: color_data = Z;
		19'b0010011110100001011: color_data = Z;
		19'b0010011110100001100: color_data = Z;
		19'b0010011110100001101: color_data = Z;
		19'b0010011110100001110: color_data = Z;
		19'b0010011110100001111: color_data = Z;
		19'b0010011110100010000: color_data = Z;
		19'b0010011110100010001: color_data = Z;
		19'b0010011110100010010: color_data = Z;
		19'b0010011110100010011: color_data = Z;
		19'b0010011110100010100: color_data = Z;
		19'b0010011110100010101: color_data = Z;
		19'b0010011110100010110: color_data = Z;
		19'b0010011110100010111: color_data = Z;
		19'b0010011110100011000: color_data = Z;
		19'b0010011110100011001: color_data = Z;
		19'b0010011110100011010: color_data = Z;
		19'b0010011110100011011: color_data = Z;
		19'b0010011110100011100: color_data = Z;
		19'b0010011110100011101: color_data = Z;
		19'b0010011110100011110: color_data = Z;
		19'b0010011110100011111: color_data = Z;
		19'b0010011110100100000: color_data = Z;
		19'b0010011110100100001: color_data = Z;
		19'b0010011110100100010: color_data = Z;
		19'b0010011110100100011: color_data = Z;
		19'b0010011110100100100: color_data = Z;
		19'b0010011110100100101: color_data = Z;
		19'b0010011110100100110: color_data = Z;
		19'b0010011110100100111: color_data = Z;
		19'b0010011110100101000: color_data = Z;
		19'b0010011110100101001: color_data = Z;
		19'b0010011110100101010: color_data = Z;
		19'b0010011110100101011: color_data = Z;
		19'b0010011110100101100: color_data = Z;
		19'b0010011110100101101: color_data = Z;
		19'b0010011110100101110: color_data = Z;
		19'b0010011110100101111: color_data = Z;
		19'b0010011110100110000: color_data = Z;
		19'b0010011110100110001: color_data = Z;
		19'b0010011110100110010: color_data = Z;
		19'b0010011110100110011: color_data = Z;
		19'b0010011110100110100: color_data = Z;
		19'b0010011110100110101: color_data = Z;
		19'b0010011110100110110: color_data = Z;
		19'b0010011110100110111: color_data = Z;
		19'b0010011110100111000: color_data = Z;
		19'b0010011110100111001: color_data = Z;
		19'b0010011110100111010: color_data = Z;
		19'b0010011110100111011: color_data = Z;
		19'b0010011110100111100: color_data = Z;
		19'b0010011110100111101: color_data = Z;
		19'b0010011110100111110: color_data = Z;
		19'b0010011110100111111: color_data = Z;
		19'b0010011110101000000: color_data = Z;
		19'b0010011110101000001: color_data = Z;
		19'b0010011110101000010: color_data = Z;
		19'b0010011110101000011: color_data = Z;
		19'b0010011110101000100: color_data = Z;
		19'b0010011110101000101: color_data = Z;
		19'b0010011110101000110: color_data = Z;
		19'b0010011110101000111: color_data = Z;
		19'b0010011110101001000: color_data = Z;
		19'b0010011110101001001: color_data = Z;
		19'b0010011110101001010: color_data = Z;
		19'b0010011110101001011: color_data = Z;
		19'b0010011110101001100: color_data = Z;
		19'b0010011110101001101: color_data = Z;
		19'b0010011110101001110: color_data = Z;
		19'b0010011110101001111: color_data = Z;
		19'b0010011110101010000: color_data = Z;
		19'b0010011110101010001: color_data = Z;
		19'b0010011110101010010: color_data = Z;
		19'b0010011110101010011: color_data = Z;
		19'b0010011110101010100: color_data = Z;
		19'b0010011110101010101: color_data = Z;
		19'b0010011110101010110: color_data = Z;
		19'b0010011110101010111: color_data = Z;
		19'b0010011110101011000: color_data = Z;
		19'b0010011110101011001: color_data = Z;
		19'b0010011110101011010: color_data = Z;
		19'b0010011110101011011: color_data = Z;
		19'b0010011110101011100: color_data = Z;
		19'b0010011110101011101: color_data = Z;
		19'b0010011110101011110: color_data = Z;
		19'b0010011110101011111: color_data = Z;
		19'b0010011110101100000: color_data = Z;
		19'b0010011110101100001: color_data = Z;
		19'b0010011110101100010: color_data = Z;
		19'b0010011110101100011: color_data = Z;
		19'b0010011110101100100: color_data = Z;
		19'b0010011110101100101: color_data = Z;
		19'b0010011110101100110: color_data = Z;
		19'b0010011110101100111: color_data = Z;
		19'b0010011110101101000: color_data = Z;
		19'b0010011110101101001: color_data = Z;
		19'b0010011110101101010: color_data = Z;
		19'b0010011110101101011: color_data = Z;
		19'b0010011110101101100: color_data = Z;
		19'b0010011110101101101: color_data = Z;
		19'b0010011110101101110: color_data = Z;
		19'b0010011110101101111: color_data = Z;
		19'b0010011110101110000: color_data = Z;
		19'b0010011110101110001: color_data = Z;
		19'b0010011110101110010: color_data = Z;
		19'b0010011110101110011: color_data = Z;
		19'b0010011110101110100: color_data = Z;
		19'b0010011110101110101: color_data = Z;
		19'b0010011110101110110: color_data = Z;
		19'b0010011110101110111: color_data = Z;
		19'b0010011110101111000: color_data = Z;
		19'b0010011110101111001: color_data = Z;
		19'b0010011110101111010: color_data = Z;
		19'b0010011110101111011: color_data = Z;
		19'b0010011110101111100: color_data = Z;
		19'b0010011110101111101: color_data = Z;
		19'b0010011110101111110: color_data = Z;
		19'b0010011110101111111: color_data = Z;
		19'b0010011110110000000: color_data = Z;
		19'b0010011110110000001: color_data = Z;
		19'b0010011110110000010: color_data = Z;
		19'b0010011110110000011: color_data = Z;
		19'b0010011110110000100: color_data = Z;
		19'b0010011110110000101: color_data = Z;
		19'b0010011110110000110: color_data = Z;
		19'b0010011110110000111: color_data = Z;
		19'b0010011110110001000: color_data = Z;
		19'b0010011110110001001: color_data = Z;
		19'b0010011110110001010: color_data = Z;
		19'b0010011110110001011: color_data = Z;
		19'b0010011110110001100: color_data = Z;
		19'b0010011110110001101: color_data = Z;
		19'b0010011110110001110: color_data = Z;
		19'b0010011110110001111: color_data = Z;
		19'b0010011110110010000: color_data = Z;
		19'b0010011110110010001: color_data = Z;
		19'b0010011110110010010: color_data = Z;
		19'b0010011110110010011: color_data = Z;
		19'b0010011110110010100: color_data = Z;
		19'b0010011110110010101: color_data = Z;
		19'b0010011110110010110: color_data = Z;
		19'b0010011110110010111: color_data = Z;
		19'b0010011110110011000: color_data = Z;
		19'b0010011110110011001: color_data = Z;
		19'b0010011110110011010: color_data = Z;
		19'b0010011110110011011: color_data = Z;
		19'b0010011110110011100: color_data = Z;
		19'b0010011110110011101: color_data = Z;
		19'b0010011110110011110: color_data = Z;
		19'b0010011110110011111: color_data = Z;
		19'b0010011110110100000: color_data = Z;
		19'b0010011110110100001: color_data = Z;
		19'b0010011110110100010: color_data = Z;
		19'b0010011110110100011: color_data = Z;
		19'b0010011110110100100: color_data = Z;
		19'b0010011110110100101: color_data = Z;
		19'b0010011110110100110: color_data = Z;
		19'b0010011110110100111: color_data = Z;
		19'b0010011110110101000: color_data = Z;
		19'b0010011110110101001: color_data = Z;
		19'b0010011110110101010: color_data = Z;
		19'b0010011110110101011: color_data = Z;
		19'b0010011110110101100: color_data = Z;
		19'b0010011110110101101: color_data = Z;
		19'b0010011110110101110: color_data = Z;
		19'b0010011110110110011: color_data = Z;
		19'b0010011110110110100: color_data = Z;
		19'b0010011110110110101: color_data = Z;
		19'b0010011110110110110: color_data = Z;
		19'b0010011110110110111: color_data = Z;
		19'b0010011110110111000: color_data = Z;
		19'b0010011110110111001: color_data = Z;
		19'b0010011110110111101: color_data = Z;
		19'b0010011110110111110: color_data = Z;
		19'b0010011110110111111: color_data = Z;
		19'b0010011110111000000: color_data = Z;
		19'b0010011110111000001: color_data = Z;
		19'b0010011110111000010: color_data = Z;
		19'b0010011110111000011: color_data = Z;
		19'b0010011110111000100: color_data = Z;
		19'b0010011110111000101: color_data = Z;
		19'b0010011110111000110: color_data = Z;
		19'b0010011110111000111: color_data = Z;
		19'b0010011110111001000: color_data = Z;
		19'b0010011110111001001: color_data = Z;
		19'b0010100000011001010: color_data = Z;
		19'b0010100000011001011: color_data = Z;
		19'b0010100000011001100: color_data = Z;
		19'b0010100000011001101: color_data = Z;
		19'b0010100000011001110: color_data = Z;
		19'b0010100000011001111: color_data = Z;
		19'b0010100000011010000: color_data = Z;
		19'b0010100000011010001: color_data = Z;
		19'b0010100000011010010: color_data = Z;
		19'b0010100000011010011: color_data = Z;
		19'b0010100000011010100: color_data = Z;
		19'b0010100000011010101: color_data = Z;
		19'b0010100000011010110: color_data = Z;
		19'b0010100000011010111: color_data = Z;
		19'b0010100000011011000: color_data = Z;
		19'b0010100000011011001: color_data = Z;
		19'b0010100000011011010: color_data = Z;
		19'b0010100000011011011: color_data = Z;
		19'b0010100000011011100: color_data = Z;
		19'b0010100000011011101: color_data = Z;
		19'b0010100000011011110: color_data = Z;
		19'b0010100000011011111: color_data = Z;
		19'b0010100000011100000: color_data = Z;
		19'b0010100000011100001: color_data = Z;
		19'b0010100000011100010: color_data = Z;
		19'b0010100000011100011: color_data = Z;
		19'b0010100000011100100: color_data = Z;
		19'b0010100000011100101: color_data = Z;
		19'b0010100000011100110: color_data = Z;
		19'b0010100000011100111: color_data = Z;
		19'b0010100000011101000: color_data = Z;
		19'b0010100000011101001: color_data = Z;
		19'b0010100000011101010: color_data = Z;
		19'b0010100000011101011: color_data = Z;
		19'b0010100000011101100: color_data = Z;
		19'b0010100000011101101: color_data = Z;
		19'b0010100000011101110: color_data = Z;
		19'b0010100000011101111: color_data = Z;
		19'b0010100000011110000: color_data = Z;
		19'b0010100000011110001: color_data = Z;
		19'b0010100000011110010: color_data = Z;
		19'b0010100000011110011: color_data = Z;
		19'b0010100000011110100: color_data = Z;
		19'b0010100000011110101: color_data = Z;
		19'b0010100000011110110: color_data = Z;
		19'b0010100000011110111: color_data = Z;
		19'b0010100000011111000: color_data = Z;
		19'b0010100000011111001: color_data = Z;
		19'b0010100000011111010: color_data = Z;
		19'b0010100000011111011: color_data = Z;
		19'b0010100000011111100: color_data = Z;
		19'b0010100000011111101: color_data = Z;
		19'b0010100000011111110: color_data = Z;
		19'b0010100000011111111: color_data = Z;
		19'b0010100000100000000: color_data = Z;
		19'b0010100000100000001: color_data = Z;
		19'b0010100000100000010: color_data = Z;
		19'b0010100000100000011: color_data = Z;
		19'b0010100000100000100: color_data = Z;
		19'b0010100000100000101: color_data = Z;
		19'b0010100000100000110: color_data = Z;
		19'b0010100000100000111: color_data = Z;
		19'b0010100000100001000: color_data = Z;
		19'b0010100000100001001: color_data = Z;
		19'b0010100000100001010: color_data = Z;
		19'b0010100000100001011: color_data = Z;
		19'b0010100000100001100: color_data = Z;
		19'b0010100000100001101: color_data = Z;
		19'b0010100000100001110: color_data = Z;
		19'b0010100000100001111: color_data = Z;
		19'b0010100000100010000: color_data = Z;
		19'b0010100000100010001: color_data = Z;
		19'b0010100000100010010: color_data = Z;
		19'b0010100000100010011: color_data = Z;
		19'b0010100000100010100: color_data = Z;
		19'b0010100000100010101: color_data = Z;
		19'b0010100000100010110: color_data = Z;
		19'b0010100000100010111: color_data = Z;
		19'b0010100000100011000: color_data = Z;
		19'b0010100000100011001: color_data = Z;
		19'b0010100000100011010: color_data = Z;
		19'b0010100000100011011: color_data = Z;
		19'b0010100000100011100: color_data = Z;
		19'b0010100000100011101: color_data = Z;
		19'b0010100000100011110: color_data = Z;
		19'b0010100000100011111: color_data = Z;
		19'b0010100000100100000: color_data = Z;
		19'b0010100000100100001: color_data = Z;
		19'b0010100000100100010: color_data = Z;
		19'b0010100000100100011: color_data = Z;
		19'b0010100000100100100: color_data = Z;
		19'b0010100000100100101: color_data = Z;
		19'b0010100000100100110: color_data = Z;
		19'b0010100000100100111: color_data = Z;
		19'b0010100000100101000: color_data = Z;
		19'b0010100000100101001: color_data = Z;
		19'b0010100000100101010: color_data = Z;
		19'b0010100000100101011: color_data = Z;
		19'b0010100000100101100: color_data = Z;
		19'b0010100000100101101: color_data = Z;
		19'b0010100000100101110: color_data = Z;
		19'b0010100000100101111: color_data = Z;
		19'b0010100000100110000: color_data = Z;
		19'b0010100000100110001: color_data = Z;
		19'b0010100000100110010: color_data = Z;
		19'b0010100000100110011: color_data = Z;
		19'b0010100000100110100: color_data = Z;
		19'b0010100000100110101: color_data = Z;
		19'b0010100000100110110: color_data = Z;
		19'b0010100000100110111: color_data = Z;
		19'b0010100000100111000: color_data = Z;
		19'b0010100000100111001: color_data = Z;
		19'b0010100000100111010: color_data = Z;
		19'b0010100000100111011: color_data = Z;
		19'b0010100000100111100: color_data = Z;
		19'b0010100000100111101: color_data = Z;
		19'b0010100000100111110: color_data = Z;
		19'b0010100000100111111: color_data = Z;
		19'b0010100000101000000: color_data = Z;
		19'b0010100000101000001: color_data = Z;
		19'b0010100000101000010: color_data = Z;
		19'b0010100000101000011: color_data = Z;
		19'b0010100000101000100: color_data = Z;
		19'b0010100000101000101: color_data = Z;
		19'b0010100000101000110: color_data = Z;
		19'b0010100000101000111: color_data = Z;
		19'b0010100000101001000: color_data = Z;
		19'b0010100000101001001: color_data = Z;
		19'b0010100000101001010: color_data = Z;
		19'b0010100000101001011: color_data = Z;
		19'b0010100000101001100: color_data = Z;
		19'b0010100000101001101: color_data = Z;
		19'b0010100000101001110: color_data = Z;
		19'b0010100000101001111: color_data = Z;
		19'b0010100000101010000: color_data = Z;
		19'b0010100000101010001: color_data = Z;
		19'b0010100000101010010: color_data = Z;
		19'b0010100000101010011: color_data = Z;
		19'b0010100000101010100: color_data = Z;
		19'b0010100000101010101: color_data = Z;
		19'b0010100000101010110: color_data = Z;
		19'b0010100000101010111: color_data = Z;
		19'b0010100000101011000: color_data = Z;
		19'b0010100000101011001: color_data = Z;
		19'b0010100000101011010: color_data = Z;
		19'b0010100000101011011: color_data = Z;
		19'b0010100000101011100: color_data = Z;
		19'b0010100000101011101: color_data = Z;
		19'b0010100000101011110: color_data = Z;
		19'b0010100000101011111: color_data = Z;
		19'b0010100000101100000: color_data = Z;
		19'b0010100000101100001: color_data = Z;
		19'b0010100000101100010: color_data = Z;
		19'b0010100000101100011: color_data = Z;
		19'b0010100000101100100: color_data = Z;
		19'b0010100000101100101: color_data = Z;
		19'b0010100000101100110: color_data = Z;
		19'b0010100000101100111: color_data = Z;
		19'b0010100000101101000: color_data = Z;
		19'b0010100000101101001: color_data = Z;
		19'b0010100000101101010: color_data = Z;
		19'b0010100000101101011: color_data = Z;
		19'b0010100000101101100: color_data = Z;
		19'b0010100000101101101: color_data = Z;
		19'b0010100000101101110: color_data = Z;
		19'b0010100000101101111: color_data = Z;
		19'b0010100000101110000: color_data = Z;
		19'b0010100000101110001: color_data = Z;
		19'b0010100000101110010: color_data = Z;
		19'b0010100000101110011: color_data = Z;
		19'b0010100000101110100: color_data = Z;
		19'b0010100000101110101: color_data = Z;
		19'b0010100000101110110: color_data = Z;
		19'b0010100000101110111: color_data = Z;
		19'b0010100000101111000: color_data = Z;
		19'b0010100000101111001: color_data = Z;
		19'b0010100000101111010: color_data = Z;
		19'b0010100000101111011: color_data = Z;
		19'b0010100000101111100: color_data = Z;
		19'b0010100000101111101: color_data = Z;
		19'b0010100000101111110: color_data = Z;
		19'b0010100000101111111: color_data = Z;
		19'b0010100000110000000: color_data = Z;
		19'b0010100000110000001: color_data = Z;
		19'b0010100000110000010: color_data = Z;
		19'b0010100000110000011: color_data = Z;
		19'b0010100000110000100: color_data = Z;
		19'b0010100000110000101: color_data = Z;
		19'b0010100000110000110: color_data = Z;
		19'b0010100000110000111: color_data = Z;
		19'b0010100000110001000: color_data = Z;
		19'b0010100000110001001: color_data = Z;
		19'b0010100000110001010: color_data = Z;
		19'b0010100000110001011: color_data = Z;
		19'b0010100000110001100: color_data = Z;
		19'b0010100000110001101: color_data = Z;
		19'b0010100000110001110: color_data = Z;
		19'b0010100000110001111: color_data = Z;
		19'b0010100000110010000: color_data = Z;
		19'b0010100000110010001: color_data = Z;
		19'b0010100000110010010: color_data = Z;
		19'b0010100000110010011: color_data = Z;
		19'b0010100000110010100: color_data = Z;
		19'b0010100000110010101: color_data = Z;
		19'b0010100000110010110: color_data = Z;
		19'b0010100000110010111: color_data = Z;
		19'b0010100000110011000: color_data = Z;
		19'b0010100000110011001: color_data = Z;
		19'b0010100000110011010: color_data = Z;
		19'b0010100000110011011: color_data = Z;
		19'b0010100000110011100: color_data = Z;
		19'b0010100000110011101: color_data = Z;
		19'b0010100000110011110: color_data = Z;
		19'b0010100000110011111: color_data = Z;
		19'b0010100000110100000: color_data = Z;
		19'b0010100000110100001: color_data = Z;
		19'b0010100000110100010: color_data = Z;
		19'b0010100000110100011: color_data = Z;
		19'b0010100000110100100: color_data = Z;
		19'b0010100000110100101: color_data = Z;
		19'b0010100000110100110: color_data = Z;
		19'b0010100000110100111: color_data = Z;
		19'b0010100000110101000: color_data = Z;
		19'b0010100000110101001: color_data = Z;
		19'b0010100000110101010: color_data = Z;
		19'b0010100000110101011: color_data = Z;
		19'b0010100000110101100: color_data = Z;
		19'b0010100000110101101: color_data = Z;
		19'b0010100000110101110: color_data = Z;
		19'b0010100000110101111: color_data = Z;
		19'b0010100000110110100: color_data = Z;
		19'b0010100000110110101: color_data = Z;
		19'b0010100000110110110: color_data = Z;
		19'b0010100000110110111: color_data = Z;
		19'b0010100000110111000: color_data = Z;
		19'b0010100000110111001: color_data = Z;
		19'b0010100000110111010: color_data = Z;
		19'b0010100000110111110: color_data = Z;
		19'b0010100000110111111: color_data = Z;
		19'b0010100000111000000: color_data = Z;
		19'b0010100000111000001: color_data = Z;
		19'b0010100000111000010: color_data = Z;
		19'b0010100000111000011: color_data = Z;
		19'b0010100000111000100: color_data = Z;
		19'b0010100000111000101: color_data = Z;
		19'b0010100000111000110: color_data = Z;
		19'b0010100000111000111: color_data = Z;
		19'b0010100000111001000: color_data = Z;
		19'b0010100000111001001: color_data = Z;
		19'b0010100010011001001: color_data = Z;
		19'b0010100010011001010: color_data = Z;
		19'b0010100010011001011: color_data = Z;
		19'b0010100010011001100: color_data = Z;
		19'b0010100010011001101: color_data = Z;
		19'b0010100010011001110: color_data = Z;
		19'b0010100010011001111: color_data = Z;
		19'b0010100010011010000: color_data = Z;
		19'b0010100010011010001: color_data = Z;
		19'b0010100010011010010: color_data = Z;
		19'b0010100010011010011: color_data = Z;
		19'b0010100010011010100: color_data = Z;
		19'b0010100010011010101: color_data = Z;
		19'b0010100010011010110: color_data = Z;
		19'b0010100010011010111: color_data = Z;
		19'b0010100010011011000: color_data = Z;
		19'b0010100010011011001: color_data = Z;
		19'b0010100010011011010: color_data = Z;
		19'b0010100010011011011: color_data = Z;
		19'b0010100010011011100: color_data = Z;
		19'b0010100010011011101: color_data = Z;
		19'b0010100010011011110: color_data = Z;
		19'b0010100010011011111: color_data = Z;
		19'b0010100010011100000: color_data = Z;
		19'b0010100010011100001: color_data = Z;
		19'b0010100010011100010: color_data = Z;
		19'b0010100010011100011: color_data = Z;
		19'b0010100010011100100: color_data = Z;
		19'b0010100010011100101: color_data = Z;
		19'b0010100010011100110: color_data = Z;
		19'b0010100010011100111: color_data = Z;
		19'b0010100010011101000: color_data = Z;
		19'b0010100010011101001: color_data = Z;
		19'b0010100010011101010: color_data = Z;
		19'b0010100010011101011: color_data = Z;
		19'b0010100010011101100: color_data = Z;
		19'b0010100010011101101: color_data = Z;
		19'b0010100010011101110: color_data = Z;
		19'b0010100010011101111: color_data = Z;
		19'b0010100010011110000: color_data = Z;
		19'b0010100010011110001: color_data = Z;
		19'b0010100010011110010: color_data = Z;
		19'b0010100010011110011: color_data = Z;
		19'b0010100010011110100: color_data = Z;
		19'b0010100010011110101: color_data = Z;
		19'b0010100010011110110: color_data = Z;
		19'b0010100010011110111: color_data = Z;
		19'b0010100010011111000: color_data = Z;
		19'b0010100010011111001: color_data = Z;
		19'b0010100010011111010: color_data = Z;
		19'b0010100010011111011: color_data = Z;
		19'b0010100010011111100: color_data = Z;
		19'b0010100010011111101: color_data = Z;
		19'b0010100010011111110: color_data = Z;
		19'b0010100010011111111: color_data = Z;
		19'b0010100010100000000: color_data = Z;
		19'b0010100010100000001: color_data = Z;
		19'b0010100010100000010: color_data = Z;
		19'b0010100010100000011: color_data = Z;
		19'b0010100010100000100: color_data = Z;
		19'b0010100010100000101: color_data = Z;
		19'b0010100010100000110: color_data = Z;
		19'b0010100010100000111: color_data = Z;
		19'b0010100010100001000: color_data = Z;
		19'b0010100010100001001: color_data = Z;
		19'b0010100010100001010: color_data = Z;
		19'b0010100010100001011: color_data = Z;
		19'b0010100010100001100: color_data = Z;
		19'b0010100010100001101: color_data = Z;
		19'b0010100010100001110: color_data = Z;
		19'b0010100010100001111: color_data = Z;
		19'b0010100010100010000: color_data = Z;
		19'b0010100010100010001: color_data = Z;
		19'b0010100010100010010: color_data = Z;
		19'b0010100010100010011: color_data = Z;
		19'b0010100010100010100: color_data = Z;
		19'b0010100010100010101: color_data = Z;
		19'b0010100010100010110: color_data = Z;
		19'b0010100010100010111: color_data = Z;
		19'b0010100010100011000: color_data = Z;
		19'b0010100010100011001: color_data = Z;
		19'b0010100010100011010: color_data = Z;
		19'b0010100010100011011: color_data = Z;
		19'b0010100010100011100: color_data = Z;
		19'b0010100010100011101: color_data = Z;
		19'b0010100010100011110: color_data = Z;
		19'b0010100010100011111: color_data = Z;
		19'b0010100010100100000: color_data = Z;
		19'b0010100010100100001: color_data = Z;
		19'b0010100010100100010: color_data = Z;
		19'b0010100010100100011: color_data = Z;
		19'b0010100010100100100: color_data = Z;
		19'b0010100010100100101: color_data = Z;
		19'b0010100010100100110: color_data = Z;
		19'b0010100010100100111: color_data = Z;
		19'b0010100010100101000: color_data = Z;
		19'b0010100010100101001: color_data = Z;
		19'b0010100010100101010: color_data = Z;
		19'b0010100010100101011: color_data = Z;
		19'b0010100010100101100: color_data = Z;
		19'b0010100010100101101: color_data = Z;
		19'b0010100010100101110: color_data = Z;
		19'b0010100010100101111: color_data = Z;
		19'b0010100010100110000: color_data = Z;
		19'b0010100010100110001: color_data = Z;
		19'b0010100010100110010: color_data = Z;
		19'b0010100010100110011: color_data = Z;
		19'b0010100010100110100: color_data = Z;
		19'b0010100010100110101: color_data = Z;
		19'b0010100010100110110: color_data = Z;
		19'b0010100010100110111: color_data = Z;
		19'b0010100010100111000: color_data = Z;
		19'b0010100010100111001: color_data = Z;
		19'b0010100010100111010: color_data = Z;
		19'b0010100010100111011: color_data = Z;
		19'b0010100010100111100: color_data = Z;
		19'b0010100010100111101: color_data = Z;
		19'b0010100010100111110: color_data = Z;
		19'b0010100010100111111: color_data = Z;
		19'b0010100010101000000: color_data = Z;
		19'b0010100010101000001: color_data = Z;
		19'b0010100010101000010: color_data = Z;
		19'b0010100010101000011: color_data = Z;
		19'b0010100010101000100: color_data = Z;
		19'b0010100010101000101: color_data = Z;
		19'b0010100010101000110: color_data = Z;
		19'b0010100010101000111: color_data = Z;
		19'b0010100010101001000: color_data = Z;
		19'b0010100010101001001: color_data = Z;
		19'b0010100010101001010: color_data = Z;
		19'b0010100010101001011: color_data = Z;
		19'b0010100010101001100: color_data = Z;
		19'b0010100010101001101: color_data = Z;
		19'b0010100010101001110: color_data = Z;
		19'b0010100010101001111: color_data = Z;
		19'b0010100010101010000: color_data = Z;
		19'b0010100010101010001: color_data = Z;
		19'b0010100010101010010: color_data = Z;
		19'b0010100010101010011: color_data = Z;
		19'b0010100010101010100: color_data = Z;
		19'b0010100010101010101: color_data = Z;
		19'b0010100010101010110: color_data = Z;
		19'b0010100010101010111: color_data = Z;
		19'b0010100010101011000: color_data = Z;
		19'b0010100010101011001: color_data = Z;
		19'b0010100010101011010: color_data = Z;
		19'b0010100010101011011: color_data = Z;
		19'b0010100010101011100: color_data = Z;
		19'b0010100010101011101: color_data = Z;
		19'b0010100010101011110: color_data = Z;
		19'b0010100010101011111: color_data = Z;
		19'b0010100010101100000: color_data = Z;
		19'b0010100010101100001: color_data = Z;
		19'b0010100010101100010: color_data = Z;
		19'b0010100010101100011: color_data = Z;
		19'b0010100010101100100: color_data = Z;
		19'b0010100010101100101: color_data = Z;
		19'b0010100010101100110: color_data = Z;
		19'b0010100010101100111: color_data = Z;
		19'b0010100010101101000: color_data = Z;
		19'b0010100010101101001: color_data = Z;
		19'b0010100010101101010: color_data = Z;
		19'b0010100010101101011: color_data = Z;
		19'b0010100010101101100: color_data = Z;
		19'b0010100010101101101: color_data = Z;
		19'b0010100010101101110: color_data = Z;
		19'b0010100010101101111: color_data = Z;
		19'b0010100010101110000: color_data = Z;
		19'b0010100010101110001: color_data = Z;
		19'b0010100010101110010: color_data = Z;
		19'b0010100010101110011: color_data = Z;
		19'b0010100010101110100: color_data = Z;
		19'b0010100010101110101: color_data = Z;
		19'b0010100010101110110: color_data = Z;
		19'b0010100010101110111: color_data = Z;
		19'b0010100010101111000: color_data = Z;
		19'b0010100010101111001: color_data = Z;
		19'b0010100010101111010: color_data = Z;
		19'b0010100010101111011: color_data = Z;
		19'b0010100010101111100: color_data = Z;
		19'b0010100010101111101: color_data = Z;
		19'b0010100010101111110: color_data = Z;
		19'b0010100010101111111: color_data = Z;
		19'b0010100010110000000: color_data = Z;
		19'b0010100010110000001: color_data = Z;
		19'b0010100010110000010: color_data = Z;
		19'b0010100010110000011: color_data = Z;
		19'b0010100010110000100: color_data = Z;
		19'b0010100010110000101: color_data = Z;
		19'b0010100010110000110: color_data = Z;
		19'b0010100010110000111: color_data = Z;
		19'b0010100010110001000: color_data = Z;
		19'b0010100010110001001: color_data = Z;
		19'b0010100010110001010: color_data = Z;
		19'b0010100010110001011: color_data = Z;
		19'b0010100010110001100: color_data = Z;
		19'b0010100010110001101: color_data = Z;
		19'b0010100010110001110: color_data = Z;
		19'b0010100010110001111: color_data = Z;
		19'b0010100010110010000: color_data = Z;
		19'b0010100010110010001: color_data = Z;
		19'b0010100010110010010: color_data = Z;
		19'b0010100010110010011: color_data = Z;
		19'b0010100010110010100: color_data = Z;
		19'b0010100010110010101: color_data = Z;
		19'b0010100010110010110: color_data = Z;
		19'b0010100010110010111: color_data = Z;
		19'b0010100010110011000: color_data = Z;
		19'b0010100010110011001: color_data = Z;
		19'b0010100010110011010: color_data = Z;
		19'b0010100010110011011: color_data = Z;
		19'b0010100010110011100: color_data = Z;
		19'b0010100010110011101: color_data = Z;
		19'b0010100010110011110: color_data = Z;
		19'b0010100010110011111: color_data = Z;
		19'b0010100010110100000: color_data = Z;
		19'b0010100010110100001: color_data = Z;
		19'b0010100010110100010: color_data = Z;
		19'b0010100010110100011: color_data = Z;
		19'b0010100010110100100: color_data = Z;
		19'b0010100010110100101: color_data = Z;
		19'b0010100010110100110: color_data = Z;
		19'b0010100010110100111: color_data = Z;
		19'b0010100010110101000: color_data = Z;
		19'b0010100010110101001: color_data = Z;
		19'b0010100010110101010: color_data = Z;
		19'b0010100010110101011: color_data = Z;
		19'b0010100010110101100: color_data = Z;
		19'b0010100010110101101: color_data = Z;
		19'b0010100010110101110: color_data = Z;
		19'b0010100010110101111: color_data = Z;
		19'b0010100010110110100: color_data = Z;
		19'b0010100010110110101: color_data = Z;
		19'b0010100010110110110: color_data = Z;
		19'b0010100010110110111: color_data = Z;
		19'b0010100010110111000: color_data = Z;
		19'b0010100010110111001: color_data = Z;
		19'b0010100010110111010: color_data = Z;
		19'b0010100010110111011: color_data = Z;
		19'b0010100010110111100: color_data = Z;
		19'b0010100010110111111: color_data = Z;
		19'b0010100010111000000: color_data = Z;
		19'b0010100010111000001: color_data = Z;
		19'b0010100010111000010: color_data = Z;
		19'b0010100010111000011: color_data = Z;
		19'b0010100010111000100: color_data = Z;
		19'b0010100010111000101: color_data = Z;
		19'b0010100010111000110: color_data = Z;
		19'b0010100010111000111: color_data = Z;
		19'b0010100010111001000: color_data = Z;
		19'b0010100010111001001: color_data = Z;
		19'b0010100100011001000: color_data = Z;
		19'b0010100100011001001: color_data = Z;
		19'b0010100100011001010: color_data = Z;
		19'b0010100100011001011: color_data = Z;
		19'b0010100100011001100: color_data = Z;
		19'b0010100100011001101: color_data = Z;
		19'b0010100100011001110: color_data = Z;
		19'b0010100100011001111: color_data = Z;
		19'b0010100100011010000: color_data = Z;
		19'b0010100100011010001: color_data = Z;
		19'b0010100100011010010: color_data = Z;
		19'b0010100100011010011: color_data = Z;
		19'b0010100100011010100: color_data = Z;
		19'b0010100100011010101: color_data = Z;
		19'b0010100100011010110: color_data = Z;
		19'b0010100100011010111: color_data = Z;
		19'b0010100100011011000: color_data = Z;
		19'b0010100100011011001: color_data = Z;
		19'b0010100100011011010: color_data = Z;
		19'b0010100100011011011: color_data = Z;
		19'b0010100100011011100: color_data = Z;
		19'b0010100100011011101: color_data = Z;
		19'b0010100100011011110: color_data = Z;
		19'b0010100100011011111: color_data = Z;
		19'b0010100100011100000: color_data = Z;
		19'b0010100100011100001: color_data = Z;
		19'b0010100100011100010: color_data = Z;
		19'b0010100100011100011: color_data = Z;
		19'b0010100100011100100: color_data = Z;
		19'b0010100100011100101: color_data = Z;
		19'b0010100100011100110: color_data = Z;
		19'b0010100100011100111: color_data = Z;
		19'b0010100100011101000: color_data = Z;
		19'b0010100100011101001: color_data = Z;
		19'b0010100100011101010: color_data = Z;
		19'b0010100100011101011: color_data = Z;
		19'b0010100100011101100: color_data = Z;
		19'b0010100100011101101: color_data = Z;
		19'b0010100100011101110: color_data = Z;
		19'b0010100100011101111: color_data = Z;
		19'b0010100100011110000: color_data = Z;
		19'b0010100100011110001: color_data = Z;
		19'b0010100100011110010: color_data = Z;
		19'b0010100100011110011: color_data = Z;
		19'b0010100100011110100: color_data = Z;
		19'b0010100100011110101: color_data = Z;
		19'b0010100100011110110: color_data = Z;
		19'b0010100100011110111: color_data = Z;
		19'b0010100100011111000: color_data = Z;
		19'b0010100100011111001: color_data = Z;
		19'b0010100100011111010: color_data = Z;
		19'b0010100100011111011: color_data = Z;
		19'b0010100100011111100: color_data = Z;
		19'b0010100100011111101: color_data = Z;
		19'b0010100100011111110: color_data = Z;
		19'b0010100100011111111: color_data = Z;
		19'b0010100100100000000: color_data = Z;
		19'b0010100100100000001: color_data = Z;
		19'b0010100100100000010: color_data = Z;
		19'b0010100100100000011: color_data = Z;
		19'b0010100100100000100: color_data = Z;
		19'b0010100100100000101: color_data = Z;
		19'b0010100100100000110: color_data = Z;
		19'b0010100100100000111: color_data = Z;
		19'b0010100100100001000: color_data = Z;
		19'b0010100100100001001: color_data = Z;
		19'b0010100100100001010: color_data = Z;
		19'b0010100100100001011: color_data = Z;
		19'b0010100100100001100: color_data = Z;
		19'b0010100100100001101: color_data = Z;
		19'b0010100100100001110: color_data = Z;
		19'b0010100100100001111: color_data = Z;
		19'b0010100100100010000: color_data = Z;
		19'b0010100100100010001: color_data = Z;
		19'b0010100100100010010: color_data = Z;
		19'b0010100100100010011: color_data = Z;
		19'b0010100100100010100: color_data = Z;
		19'b0010100100100010101: color_data = Z;
		19'b0010100100100010110: color_data = Z;
		19'b0010100100100010111: color_data = Z;
		19'b0010100100100011000: color_data = Z;
		19'b0010100100100011001: color_data = Z;
		19'b0010100100100011010: color_data = Z;
		19'b0010100100100011011: color_data = Z;
		19'b0010100100100011100: color_data = Z;
		19'b0010100100100011101: color_data = Z;
		19'b0010100100100011110: color_data = Z;
		19'b0010100100100011111: color_data = Z;
		19'b0010100100100100000: color_data = Z;
		19'b0010100100100100001: color_data = Z;
		19'b0010100100100100010: color_data = Z;
		19'b0010100100100100011: color_data = Z;
		19'b0010100100100100100: color_data = Z;
		19'b0010100100100100101: color_data = Z;
		19'b0010100100100100110: color_data = Z;
		19'b0010100100100100111: color_data = Z;
		19'b0010100100100101000: color_data = Z;
		19'b0010100100100101001: color_data = Z;
		19'b0010100100100101010: color_data = Z;
		19'b0010100100100101011: color_data = Z;
		19'b0010100100100101100: color_data = Z;
		19'b0010100100100101101: color_data = Z;
		19'b0010100100100101110: color_data = Z;
		19'b0010100100100101111: color_data = Z;
		19'b0010100100100110000: color_data = Z;
		19'b0010100100100110001: color_data = Z;
		19'b0010100100100110010: color_data = Z;
		19'b0010100100100110011: color_data = Z;
		19'b0010100100100110100: color_data = Z;
		19'b0010100100100110101: color_data = Z;
		19'b0010100100100110110: color_data = Z;
		19'b0010100100100110111: color_data = Z;
		19'b0010100100100111000: color_data = Z;
		19'b0010100100100111001: color_data = Z;
		19'b0010100100100111010: color_data = Z;
		19'b0010100100100111011: color_data = Z;
		19'b0010100100100111100: color_data = Z;
		19'b0010100100100111101: color_data = Z;
		19'b0010100100100111110: color_data = Z;
		19'b0010100100100111111: color_data = Z;
		19'b0010100100101000000: color_data = Z;
		19'b0010100100101000001: color_data = Z;
		19'b0010100100101000010: color_data = Z;
		19'b0010100100101000011: color_data = Z;
		19'b0010100100101000100: color_data = Z;
		19'b0010100100101000101: color_data = Z;
		19'b0010100100101000110: color_data = Z;
		19'b0010100100101000111: color_data = Z;
		19'b0010100100101001000: color_data = Z;
		19'b0010100100101001001: color_data = Z;
		19'b0010100100101001010: color_data = Z;
		19'b0010100100101001011: color_data = Z;
		19'b0010100100101001100: color_data = Z;
		19'b0010100100101001101: color_data = Z;
		19'b0010100100101001110: color_data = Z;
		19'b0010100100101001111: color_data = Z;
		19'b0010100100101010000: color_data = Z;
		19'b0010100100101010001: color_data = Z;
		19'b0010100100101010010: color_data = Z;
		19'b0010100100101010011: color_data = Z;
		19'b0010100100101010100: color_data = Z;
		19'b0010100100101010101: color_data = Z;
		19'b0010100100101010110: color_data = Z;
		19'b0010100100101010111: color_data = Z;
		19'b0010100100101011000: color_data = Z;
		19'b0010100100101011001: color_data = Z;
		19'b0010100100101011010: color_data = Z;
		19'b0010100100101011011: color_data = Z;
		19'b0010100100101011100: color_data = Z;
		19'b0010100100101011101: color_data = Z;
		19'b0010100100101011110: color_data = Z;
		19'b0010100100101011111: color_data = Z;
		19'b0010100100101100000: color_data = Z;
		19'b0010100100101100001: color_data = Z;
		19'b0010100100101100010: color_data = Z;
		19'b0010100100101100011: color_data = Z;
		19'b0010100100101100100: color_data = Z;
		19'b0010100100101100101: color_data = Z;
		19'b0010100100101100110: color_data = Z;
		19'b0010100100101100111: color_data = Z;
		19'b0010100100101101000: color_data = Z;
		19'b0010100100101101001: color_data = Z;
		19'b0010100100101101010: color_data = Z;
		19'b0010100100101101011: color_data = Z;
		19'b0010100100101101100: color_data = Z;
		19'b0010100100101101101: color_data = Z;
		19'b0010100100101101110: color_data = Z;
		19'b0010100100101101111: color_data = Z;
		19'b0010100100101110000: color_data = Z;
		19'b0010100100101110001: color_data = Z;
		19'b0010100100101110010: color_data = Z;
		19'b0010100100101110011: color_data = Z;
		19'b0010100100101110100: color_data = Z;
		19'b0010100100101110101: color_data = Z;
		19'b0010100100101110110: color_data = Z;
		19'b0010100100101110111: color_data = Z;
		19'b0010100100101111000: color_data = Z;
		19'b0010100100101111001: color_data = Z;
		19'b0010100100101111010: color_data = Z;
		19'b0010100100101111011: color_data = Z;
		19'b0010100100101111100: color_data = Z;
		19'b0010100100101111101: color_data = Z;
		19'b0010100100101111110: color_data = Z;
		19'b0010100100101111111: color_data = Z;
		19'b0010100100110000000: color_data = Z;
		19'b0010100100110000001: color_data = Z;
		19'b0010100100110000010: color_data = Z;
		19'b0010100100110000011: color_data = Z;
		19'b0010100100110000100: color_data = Z;
		19'b0010100100110000101: color_data = Z;
		19'b0010100100110000110: color_data = Z;
		19'b0010100100110000111: color_data = Z;
		19'b0010100100110001000: color_data = Z;
		19'b0010100100110001001: color_data = Z;
		19'b0010100100110001010: color_data = Z;
		19'b0010100100110001011: color_data = Z;
		19'b0010100100110001100: color_data = Z;
		19'b0010100100110001101: color_data = Z;
		19'b0010100100110001110: color_data = Z;
		19'b0010100100110001111: color_data = Z;
		19'b0010100100110010000: color_data = Z;
		19'b0010100100110010001: color_data = Z;
		19'b0010100100110010010: color_data = Z;
		19'b0010100100110010011: color_data = Z;
		19'b0010100100110010100: color_data = Z;
		19'b0010100100110010101: color_data = Z;
		19'b0010100100110010110: color_data = Z;
		19'b0010100100110010111: color_data = Z;
		19'b0010100100110011000: color_data = Z;
		19'b0010100100110011001: color_data = Z;
		19'b0010100100110011010: color_data = Z;
		19'b0010100100110011011: color_data = Z;
		19'b0010100100110011100: color_data = Z;
		19'b0010100100110011101: color_data = Z;
		19'b0010100100110011110: color_data = Z;
		19'b0010100100110011111: color_data = Z;
		19'b0010100100110100000: color_data = Z;
		19'b0010100100110100001: color_data = Z;
		19'b0010100100110100010: color_data = Z;
		19'b0010100100110100011: color_data = Z;
		19'b0010100100110100100: color_data = Z;
		19'b0010100100110100101: color_data = Z;
		19'b0010100100110100110: color_data = Z;
		19'b0010100100110100111: color_data = Z;
		19'b0010100100110101000: color_data = Z;
		19'b0010100100110101001: color_data = Z;
		19'b0010100100110101010: color_data = Z;
		19'b0010100100110101011: color_data = Z;
		19'b0010100100110101100: color_data = Z;
		19'b0010100100110101101: color_data = Z;
		19'b0010100100110101110: color_data = Z;
		19'b0010100100110101111: color_data = Z;
		19'b0010100100110110000: color_data = Z;
		19'b0010100100110110101: color_data = Z;
		19'b0010100100110110110: color_data = Z;
		19'b0010100100110110111: color_data = Z;
		19'b0010100100110111000: color_data = Z;
		19'b0010100100110111001: color_data = Z;
		19'b0010100100110111010: color_data = Z;
		19'b0010100100110111011: color_data = Z;
		19'b0010100100110111100: color_data = Z;
		19'b0010100100110111101: color_data = Z;
		19'b0010100100111000000: color_data = Z;
		19'b0010100100111000001: color_data = Z;
		19'b0010100100111000010: color_data = Z;
		19'b0010100100111000011: color_data = Z;
		19'b0010100100111000100: color_data = Z;
		19'b0010100100111000101: color_data = Z;
		19'b0010100100111000110: color_data = Z;
		19'b0010100100111000111: color_data = Z;
		19'b0010100100111001000: color_data = Z;
		19'b0010100100111001001: color_data = Z;
		19'b0010100100111001010: color_data = Z;
		19'b0010100110011001000: color_data = Z;
		19'b0010100110011001001: color_data = Z;
		19'b0010100110011001010: color_data = Z;
		19'b0010100110011001011: color_data = Z;
		19'b0010100110011001100: color_data = Z;
		19'b0010100110011001101: color_data = Z;
		19'b0010100110011001110: color_data = Z;
		19'b0010100110011001111: color_data = Z;
		19'b0010100110011010000: color_data = Z;
		19'b0010100110011010001: color_data = Z;
		19'b0010100110011010010: color_data = Z;
		19'b0010100110011010011: color_data = Z;
		19'b0010100110011010100: color_data = Z;
		19'b0010100110011010101: color_data = Z;
		19'b0010100110011010110: color_data = Z;
		19'b0010100110011010111: color_data = Z;
		19'b0010100110011011000: color_data = Z;
		19'b0010100110011011001: color_data = Z;
		19'b0010100110011011010: color_data = Z;
		19'b0010100110011011011: color_data = Z;
		19'b0010100110011011100: color_data = Z;
		19'b0010100110011011101: color_data = Z;
		19'b0010100110011011110: color_data = Z;
		19'b0010100110011011111: color_data = Z;
		19'b0010100110011100000: color_data = Z;
		19'b0010100110011100001: color_data = Z;
		19'b0010100110011100010: color_data = Z;
		19'b0010100110011100011: color_data = Z;
		19'b0010100110011100100: color_data = Z;
		19'b0010100110011100101: color_data = Z;
		19'b0010100110011100110: color_data = Z;
		19'b0010100110011100111: color_data = Z;
		19'b0010100110011101000: color_data = Z;
		19'b0010100110011101001: color_data = Z;
		19'b0010100110011101010: color_data = Z;
		19'b0010100110011101011: color_data = Z;
		19'b0010100110011101100: color_data = Z;
		19'b0010100110011101101: color_data = Z;
		19'b0010100110011101110: color_data = Z;
		19'b0010100110011101111: color_data = Z;
		19'b0010100110011110000: color_data = Z;
		19'b0010100110011110001: color_data = Z;
		19'b0010100110011110010: color_data = Z;
		19'b0010100110011110011: color_data = Z;
		19'b0010100110011110100: color_data = Z;
		19'b0010100110011110101: color_data = Z;
		19'b0010100110011110110: color_data = Z;
		19'b0010100110011110111: color_data = Z;
		19'b0010100110011111000: color_data = Z;
		19'b0010100110011111001: color_data = Z;
		19'b0010100110011111010: color_data = Z;
		19'b0010100110011111011: color_data = Z;
		19'b0010100110011111100: color_data = Z;
		19'b0010100110011111101: color_data = Z;
		19'b0010100110011111110: color_data = Z;
		19'b0010100110011111111: color_data = Z;
		19'b0010100110100000000: color_data = Z;
		19'b0010100110100000001: color_data = Z;
		19'b0010100110100000010: color_data = Z;
		19'b0010100110100000011: color_data = Z;
		19'b0010100110100000100: color_data = Z;
		19'b0010100110100000101: color_data = Z;
		19'b0010100110100000110: color_data = Z;
		19'b0010100110100000111: color_data = Z;
		19'b0010100110100001000: color_data = Z;
		19'b0010100110100001001: color_data = Z;
		19'b0010100110100001010: color_data = Z;
		19'b0010100110100001011: color_data = Z;
		19'b0010100110100001100: color_data = Z;
		19'b0010100110100001101: color_data = Z;
		19'b0010100110100001110: color_data = Z;
		19'b0010100110100001111: color_data = Z;
		19'b0010100110100010000: color_data = Z;
		19'b0010100110100010001: color_data = Z;
		19'b0010100110100010010: color_data = Z;
		19'b0010100110100010011: color_data = Z;
		19'b0010100110100010100: color_data = Z;
		19'b0010100110100010101: color_data = Z;
		19'b0010100110100010110: color_data = Z;
		19'b0010100110100010111: color_data = Z;
		19'b0010100110100011000: color_data = Z;
		19'b0010100110100011001: color_data = Z;
		19'b0010100110100011010: color_data = Z;
		19'b0010100110100011011: color_data = Z;
		19'b0010100110100011100: color_data = Z;
		19'b0010100110100011101: color_data = Z;
		19'b0010100110100011110: color_data = Z;
		19'b0010100110100011111: color_data = Z;
		19'b0010100110100100000: color_data = Z;
		19'b0010100110100100001: color_data = Z;
		19'b0010100110100100010: color_data = Z;
		19'b0010100110100100011: color_data = Z;
		19'b0010100110100100100: color_data = Z;
		19'b0010100110100100101: color_data = Z;
		19'b0010100110100100110: color_data = Z;
		19'b0010100110100100111: color_data = Z;
		19'b0010100110100101000: color_data = Z;
		19'b0010100110100101001: color_data = Z;
		19'b0010100110100101010: color_data = Z;
		19'b0010100110100101011: color_data = Z;
		19'b0010100110100101100: color_data = Z;
		19'b0010100110100101101: color_data = Z;
		19'b0010100110100101110: color_data = Z;
		19'b0010100110100101111: color_data = Z;
		19'b0010100110100110000: color_data = Z;
		19'b0010100110100110001: color_data = Z;
		19'b0010100110100110010: color_data = Z;
		19'b0010100110100110011: color_data = Z;
		19'b0010100110100110100: color_data = Z;
		19'b0010100110100110101: color_data = Z;
		19'b0010100110100110110: color_data = Z;
		19'b0010100110100110111: color_data = Z;
		19'b0010100110100111000: color_data = Z;
		19'b0010100110100111001: color_data = Z;
		19'b0010100110100111010: color_data = Z;
		19'b0010100110100111011: color_data = Z;
		19'b0010100110100111100: color_data = Z;
		19'b0010100110100111101: color_data = Z;
		19'b0010100110100111110: color_data = Z;
		19'b0010100110100111111: color_data = Z;
		19'b0010100110101000000: color_data = Z;
		19'b0010100110101000001: color_data = Z;
		19'b0010100110101000010: color_data = Z;
		19'b0010100110101000011: color_data = Z;
		19'b0010100110101000100: color_data = Z;
		19'b0010100110101000101: color_data = Z;
		19'b0010100110101000110: color_data = Z;
		19'b0010100110101000111: color_data = Z;
		19'b0010100110101001000: color_data = Z;
		19'b0010100110101001001: color_data = Z;
		19'b0010100110101001010: color_data = Z;
		19'b0010100110101001011: color_data = Z;
		19'b0010100110101001100: color_data = Z;
		19'b0010100110101001101: color_data = Z;
		19'b0010100110101001110: color_data = Z;
		19'b0010100110101001111: color_data = Z;
		19'b0010100110101010000: color_data = Z;
		19'b0010100110101010001: color_data = Z;
		19'b0010100110101010010: color_data = Z;
		19'b0010100110101010011: color_data = Z;
		19'b0010100110101010100: color_data = Z;
		19'b0010100110101010101: color_data = Z;
		19'b0010100110101010110: color_data = Z;
		19'b0010100110101010111: color_data = Z;
		19'b0010100110101011000: color_data = Z;
		19'b0010100110101011001: color_data = Z;
		19'b0010100110101011010: color_data = Z;
		19'b0010100110101011011: color_data = Z;
		19'b0010100110101011100: color_data = Z;
		19'b0010100110101011101: color_data = Z;
		19'b0010100110101011110: color_data = Z;
		19'b0010100110101011111: color_data = Z;
		19'b0010100110101100000: color_data = Z;
		19'b0010100110101100001: color_data = Z;
		19'b0010100110101100010: color_data = Z;
		19'b0010100110101100011: color_data = Z;
		19'b0010100110101100100: color_data = Z;
		19'b0010100110101100101: color_data = Z;
		19'b0010100110101100110: color_data = Z;
		19'b0010100110101100111: color_data = Z;
		19'b0010100110101101000: color_data = Z;
		19'b0010100110101101001: color_data = Z;
		19'b0010100110101101010: color_data = Z;
		19'b0010100110101101011: color_data = Z;
		19'b0010100110101101100: color_data = Z;
		19'b0010100110101101101: color_data = Z;
		19'b0010100110101101110: color_data = Z;
		19'b0010100110101101111: color_data = Z;
		19'b0010100110101110000: color_data = Z;
		19'b0010100110101110001: color_data = Z;
		19'b0010100110101110010: color_data = Z;
		19'b0010100110101110011: color_data = Z;
		19'b0010100110101110100: color_data = Z;
		19'b0010100110101110101: color_data = Z;
		19'b0010100110101110110: color_data = Z;
		19'b0010100110101110111: color_data = Z;
		19'b0010100110101111000: color_data = Z;
		19'b0010100110101111001: color_data = Z;
		19'b0010100110101111010: color_data = Z;
		19'b0010100110101111011: color_data = Z;
		19'b0010100110101111100: color_data = Z;
		19'b0010100110101111101: color_data = Z;
		19'b0010100110101111110: color_data = Z;
		19'b0010100110101111111: color_data = Z;
		19'b0010100110110000000: color_data = Z;
		19'b0010100110110000001: color_data = Z;
		19'b0010100110110000010: color_data = Z;
		19'b0010100110110000011: color_data = Z;
		19'b0010100110110000100: color_data = Z;
		19'b0010100110110000101: color_data = Z;
		19'b0010100110110000110: color_data = Z;
		19'b0010100110110000111: color_data = Z;
		19'b0010100110110001000: color_data = Z;
		19'b0010100110110001001: color_data = Z;
		19'b0010100110110001010: color_data = Z;
		19'b0010100110110001011: color_data = Z;
		19'b0010100110110001100: color_data = Z;
		19'b0010100110110001101: color_data = Z;
		19'b0010100110110001110: color_data = Z;
		19'b0010100110110001111: color_data = Z;
		19'b0010100110110010000: color_data = Z;
		19'b0010100110110010001: color_data = Z;
		19'b0010100110110010010: color_data = Z;
		19'b0010100110110010011: color_data = Z;
		19'b0010100110110010100: color_data = Z;
		19'b0010100110110010101: color_data = Z;
		19'b0010100110110010110: color_data = Z;
		19'b0010100110110010111: color_data = Z;
		19'b0010100110110011000: color_data = Z;
		19'b0010100110110011001: color_data = Z;
		19'b0010100110110011010: color_data = Z;
		19'b0010100110110011011: color_data = Z;
		19'b0010100110110011100: color_data = Z;
		19'b0010100110110011101: color_data = Z;
		19'b0010100110110011110: color_data = Z;
		19'b0010100110110011111: color_data = Z;
		19'b0010100110110100000: color_data = Z;
		19'b0010100110110100001: color_data = Z;
		19'b0010100110110100010: color_data = Z;
		19'b0010100110110100011: color_data = Z;
		19'b0010100110110100100: color_data = Z;
		19'b0010100110110100101: color_data = Z;
		19'b0010100110110100110: color_data = Z;
		19'b0010100110110100111: color_data = Z;
		19'b0010100110110101000: color_data = Z;
		19'b0010100110110101001: color_data = Z;
		19'b0010100110110101010: color_data = Z;
		19'b0010100110110101011: color_data = Z;
		19'b0010100110110101100: color_data = Z;
		19'b0010100110110101101: color_data = Z;
		19'b0010100110110101110: color_data = Z;
		19'b0010100110110101111: color_data = Z;
		19'b0010100110110110000: color_data = Z;
		19'b0010100110110110101: color_data = Z;
		19'b0010100110110110110: color_data = Z;
		19'b0010100110110110111: color_data = Z;
		19'b0010100110110111000: color_data = Z;
		19'b0010100110110111001: color_data = Z;
		19'b0010100110110111010: color_data = Z;
		19'b0010100110110111011: color_data = Z;
		19'b0010100110110111100: color_data = Z;
		19'b0010100110110111101: color_data = Z;
		19'b0010100110110111110: color_data = Z;
		19'b0010100110111000000: color_data = Z;
		19'b0010100110111000001: color_data = Z;
		19'b0010100110111000010: color_data = Z;
		19'b0010100110111000011: color_data = Z;
		19'b0010100110111000100: color_data = Z;
		19'b0010100110111000101: color_data = Z;
		19'b0010100110111000110: color_data = Z;
		19'b0010100110111000111: color_data = Z;
		19'b0010100110111001000: color_data = Z;
		19'b0010100110111001001: color_data = Z;
		19'b0010100110111001010: color_data = Z;
		19'b0010101000011000111: color_data = Z;
		19'b0010101000011001000: color_data = Z;
		19'b0010101000011001001: color_data = Z;
		19'b0010101000011001010: color_data = Z;
		19'b0010101000011001011: color_data = Z;
		19'b0010101000011001100: color_data = Z;
		19'b0010101000011001101: color_data = Z;
		19'b0010101000011001110: color_data = Z;
		19'b0010101000011001111: color_data = Z;
		19'b0010101000011010000: color_data = Z;
		19'b0010101000011010001: color_data = Z;
		19'b0010101000011010010: color_data = Z;
		19'b0010101000011010011: color_data = Z;
		19'b0010101000011010100: color_data = Z;
		19'b0010101000011010101: color_data = Z;
		19'b0010101000011010110: color_data = Z;
		19'b0010101000011010111: color_data = Z;
		19'b0010101000011011000: color_data = Z;
		19'b0010101000011011001: color_data = Z;
		19'b0010101000011011010: color_data = Z;
		19'b0010101000011011011: color_data = Z;
		19'b0010101000011011100: color_data = Z;
		19'b0010101000011011101: color_data = Z;
		19'b0010101000011011110: color_data = Z;
		19'b0010101000011011111: color_data = Z;
		19'b0010101000011100000: color_data = Z;
		19'b0010101000011100001: color_data = Z;
		19'b0010101000011100010: color_data = Z;
		19'b0010101000011100011: color_data = Z;
		19'b0010101000011100100: color_data = Z;
		19'b0010101000011100101: color_data = Z;
		19'b0010101000011100110: color_data = Z;
		19'b0010101000011100111: color_data = Z;
		19'b0010101000011101000: color_data = Z;
		19'b0010101000011101001: color_data = Z;
		19'b0010101000011101010: color_data = Z;
		19'b0010101000011101011: color_data = Z;
		19'b0010101000011101100: color_data = Z;
		19'b0010101000011101101: color_data = Z;
		19'b0010101000011101110: color_data = Z;
		19'b0010101000011101111: color_data = Z;
		19'b0010101000011110000: color_data = Z;
		19'b0010101000011110001: color_data = Z;
		19'b0010101000011110010: color_data = Z;
		19'b0010101000011110011: color_data = Z;
		19'b0010101000011110100: color_data = Z;
		19'b0010101000011110101: color_data = Z;
		19'b0010101000011110110: color_data = Z;
		19'b0010101000011110111: color_data = Z;
		19'b0010101000011111000: color_data = Z;
		19'b0010101000011111001: color_data = Z;
		19'b0010101000011111010: color_data = Z;
		19'b0010101000011111011: color_data = Z;
		19'b0010101000011111100: color_data = Z;
		19'b0010101000011111101: color_data = Z;
		19'b0010101000011111110: color_data = Z;
		19'b0010101000011111111: color_data = Z;
		19'b0010101000100000000: color_data = Z;
		19'b0010101000100000001: color_data = Z;
		19'b0010101000100000010: color_data = Z;
		19'b0010101000100000011: color_data = Z;
		19'b0010101000100000100: color_data = Z;
		19'b0010101000100000101: color_data = Z;
		19'b0010101000100000110: color_data = Z;
		19'b0010101000100000111: color_data = Z;
		19'b0010101000100001000: color_data = Z;
		19'b0010101000100001001: color_data = Z;
		19'b0010101000100001010: color_data = Z;
		19'b0010101000100001011: color_data = Z;
		19'b0010101000100001100: color_data = Z;
		19'b0010101000100001101: color_data = Z;
		19'b0010101000100001110: color_data = Z;
		19'b0010101000100001111: color_data = Z;
		19'b0010101000100010000: color_data = Z;
		19'b0010101000100010001: color_data = Z;
		19'b0010101000100010010: color_data = Z;
		19'b0010101000100010011: color_data = Z;
		19'b0010101000100010100: color_data = Z;
		19'b0010101000100010101: color_data = Z;
		19'b0010101000100010110: color_data = Z;
		19'b0010101000100010111: color_data = Z;
		19'b0010101000100011000: color_data = Z;
		19'b0010101000100011001: color_data = Z;
		19'b0010101000100011010: color_data = Z;
		19'b0010101000100011011: color_data = Z;
		19'b0010101000100011100: color_data = Z;
		19'b0010101000100011101: color_data = Z;
		19'b0010101000100011110: color_data = Z;
		19'b0010101000100011111: color_data = Z;
		19'b0010101000100100000: color_data = Z;
		19'b0010101000100100001: color_data = Z;
		19'b0010101000100100010: color_data = Z;
		19'b0010101000100100011: color_data = Z;
		19'b0010101000100100100: color_data = Z;
		19'b0010101000100100101: color_data = Z;
		19'b0010101000100100110: color_data = Z;
		19'b0010101000100100111: color_data = Z;
		19'b0010101000100101000: color_data = Z;
		19'b0010101000100101001: color_data = Z;
		19'b0010101000100101010: color_data = Z;
		19'b0010101000100101011: color_data = Z;
		19'b0010101000100101100: color_data = Z;
		19'b0010101000100101101: color_data = Z;
		19'b0010101000100101110: color_data = Z;
		19'b0010101000100101111: color_data = Z;
		19'b0010101000100110000: color_data = Z;
		19'b0010101000100110001: color_data = Z;
		19'b0010101000100110010: color_data = Z;
		19'b0010101000100110011: color_data = Z;
		19'b0010101000100110100: color_data = Z;
		19'b0010101000100110101: color_data = Z;
		19'b0010101000100110110: color_data = Z;
		19'b0010101000100110111: color_data = Z;
		19'b0010101000100111000: color_data = Z;
		19'b0010101000100111001: color_data = Z;
		19'b0010101000100111010: color_data = Z;
		19'b0010101000100111011: color_data = Z;
		19'b0010101000100111100: color_data = Z;
		19'b0010101000100111101: color_data = Z;
		19'b0010101000100111110: color_data = Z;
		19'b0010101000100111111: color_data = Z;
		19'b0010101000101000000: color_data = Z;
		19'b0010101000101000001: color_data = Z;
		19'b0010101000101000010: color_data = Z;
		19'b0010101000101000011: color_data = Z;
		19'b0010101000101000100: color_data = Z;
		19'b0010101000101000101: color_data = Z;
		19'b0010101000101000110: color_data = Z;
		19'b0010101000101000111: color_data = Z;
		19'b0010101000101001000: color_data = Z;
		19'b0010101000101001001: color_data = Z;
		19'b0010101000101001010: color_data = Z;
		19'b0010101000101001011: color_data = Z;
		19'b0010101000101001100: color_data = Z;
		19'b0010101000101001101: color_data = Z;
		19'b0010101000101001110: color_data = Z;
		19'b0010101000101001111: color_data = Z;
		19'b0010101000101010000: color_data = Z;
		19'b0010101000101010001: color_data = Z;
		19'b0010101000101010010: color_data = Z;
		19'b0010101000101010011: color_data = Z;
		19'b0010101000101010100: color_data = Z;
		19'b0010101000101010101: color_data = Z;
		19'b0010101000101010110: color_data = Z;
		19'b0010101000101010111: color_data = Z;
		19'b0010101000101011000: color_data = Z;
		19'b0010101000101011001: color_data = Z;
		19'b0010101000101011010: color_data = Z;
		19'b0010101000101011011: color_data = Z;
		19'b0010101000101011100: color_data = Z;
		19'b0010101000101011101: color_data = Z;
		19'b0010101000101011110: color_data = Z;
		19'b0010101000101011111: color_data = Z;
		19'b0010101000101100000: color_data = Z;
		19'b0010101000101100001: color_data = Z;
		19'b0010101000101100010: color_data = Z;
		19'b0010101000101100011: color_data = Z;
		19'b0010101000101100100: color_data = Z;
		19'b0010101000101100101: color_data = Z;
		19'b0010101000101100110: color_data = Z;
		19'b0010101000101100111: color_data = Z;
		19'b0010101000101101000: color_data = Z;
		19'b0010101000101101001: color_data = Z;
		19'b0010101000101101010: color_data = Z;
		19'b0010101000101101011: color_data = Z;
		19'b0010101000101101100: color_data = Z;
		19'b0010101000101101101: color_data = Z;
		19'b0010101000101101110: color_data = Z;
		19'b0010101000101101111: color_data = Z;
		19'b0010101000101110000: color_data = Z;
		19'b0010101000101110001: color_data = Z;
		19'b0010101000101110010: color_data = Z;
		19'b0010101000101110011: color_data = Z;
		19'b0010101000101110100: color_data = Z;
		19'b0010101000101110101: color_data = Z;
		19'b0010101000101110110: color_data = Z;
		19'b0010101000101110111: color_data = Z;
		19'b0010101000101111000: color_data = Z;
		19'b0010101000101111001: color_data = Z;
		19'b0010101000101111010: color_data = Z;
		19'b0010101000101111011: color_data = Z;
		19'b0010101000101111100: color_data = Z;
		19'b0010101000101111101: color_data = Z;
		19'b0010101000101111110: color_data = Z;
		19'b0010101000101111111: color_data = Z;
		19'b0010101000110000000: color_data = Z;
		19'b0010101000110000001: color_data = Z;
		19'b0010101000110000010: color_data = Z;
		19'b0010101000110000011: color_data = Z;
		19'b0010101000110000100: color_data = Z;
		19'b0010101000110000101: color_data = Z;
		19'b0010101000110000110: color_data = Z;
		19'b0010101000110000111: color_data = Z;
		19'b0010101000110001000: color_data = Z;
		19'b0010101000110001001: color_data = Z;
		19'b0010101000110001010: color_data = Z;
		19'b0010101000110001011: color_data = Z;
		19'b0010101000110001100: color_data = Z;
		19'b0010101000110001101: color_data = Z;
		19'b0010101000110001110: color_data = Z;
		19'b0010101000110001111: color_data = Z;
		19'b0010101000110010000: color_data = Z;
		19'b0010101000110010001: color_data = Z;
		19'b0010101000110010010: color_data = Z;
		19'b0010101000110010011: color_data = Z;
		19'b0010101000110010100: color_data = Z;
		19'b0010101000110010101: color_data = Z;
		19'b0010101000110010110: color_data = Z;
		19'b0010101000110010111: color_data = Z;
		19'b0010101000110011000: color_data = Z;
		19'b0010101000110011001: color_data = Z;
		19'b0010101000110011010: color_data = Z;
		19'b0010101000110011011: color_data = Z;
		19'b0010101000110011100: color_data = Z;
		19'b0010101000110011101: color_data = Z;
		19'b0010101000110011110: color_data = Z;
		19'b0010101000110011111: color_data = Z;
		19'b0010101000110100000: color_data = Z;
		19'b0010101000110100001: color_data = Z;
		19'b0010101000110100010: color_data = Z;
		19'b0010101000110100011: color_data = Z;
		19'b0010101000110100100: color_data = Z;
		19'b0010101000110100101: color_data = Z;
		19'b0010101000110100110: color_data = Z;
		19'b0010101000110100111: color_data = Z;
		19'b0010101000110101000: color_data = Z;
		19'b0010101000110101001: color_data = Z;
		19'b0010101000110101010: color_data = Z;
		19'b0010101000110101011: color_data = Z;
		19'b0010101000110101100: color_data = Z;
		19'b0010101000110101101: color_data = Z;
		19'b0010101000110101110: color_data = Z;
		19'b0010101000110101111: color_data = Z;
		19'b0010101000110110000: color_data = Z;
		19'b0010101000110111000: color_data = Z;
		19'b0010101000110111001: color_data = Z;
		19'b0010101000110111010: color_data = Z;
		19'b0010101000110111011: color_data = Z;
		19'b0010101000110111100: color_data = Z;
		19'b0010101000110111101: color_data = Z;
		19'b0010101000110111110: color_data = Z;
		19'b0010101000110111111: color_data = Z;
		19'b0010101000111000000: color_data = Z;
		19'b0010101000111000001: color_data = Z;
		19'b0010101000111000010: color_data = Z;
		19'b0010101000111000011: color_data = Z;
		19'b0010101000111000100: color_data = Z;
		19'b0010101000111000101: color_data = Z;
		19'b0010101000111000110: color_data = Z;
		19'b0010101000111000111: color_data = Z;
		19'b0010101000111001000: color_data = Z;
		19'b0010101000111001001: color_data = Z;
		19'b0010101000111001010: color_data = Z;
		19'b0010101000111001011: color_data = Z;
		19'b0010101010011000101: color_data = Z;
		19'b0010101010011000110: color_data = Z;
		19'b0010101010011000111: color_data = Z;
		19'b0010101010011001000: color_data = Z;
		19'b0010101010011001001: color_data = Z;
		19'b0010101010011001010: color_data = Z;
		19'b0010101010011001011: color_data = Z;
		19'b0010101010011001100: color_data = Z;
		19'b0010101010011001101: color_data = Z;
		19'b0010101010011001110: color_data = Z;
		19'b0010101010011001111: color_data = Z;
		19'b0010101010011010000: color_data = Z;
		19'b0010101010011010001: color_data = Z;
		19'b0010101010011010010: color_data = Z;
		19'b0010101010011010011: color_data = Z;
		19'b0010101010011010100: color_data = Z;
		19'b0010101010011010101: color_data = Z;
		19'b0010101010011010110: color_data = Z;
		19'b0010101010011010111: color_data = Z;
		19'b0010101010011011000: color_data = Z;
		19'b0010101010011011001: color_data = Z;
		19'b0010101010011011010: color_data = Z;
		19'b0010101010011011011: color_data = Z;
		19'b0010101010011011100: color_data = Z;
		19'b0010101010011011101: color_data = Z;
		19'b0010101010011011110: color_data = Z;
		19'b0010101010011011111: color_data = Z;
		19'b0010101010011100000: color_data = Z;
		19'b0010101010011100001: color_data = Z;
		19'b0010101010011100010: color_data = Z;
		19'b0010101010011100011: color_data = Z;
		19'b0010101010011100100: color_data = Z;
		19'b0010101010011100101: color_data = Z;
		19'b0010101010011100110: color_data = Z;
		19'b0010101010011100111: color_data = Z;
		19'b0010101010011101000: color_data = Z;
		19'b0010101010011101001: color_data = Z;
		19'b0010101010011101010: color_data = Z;
		19'b0010101010011101011: color_data = Z;
		19'b0010101010011101100: color_data = Z;
		19'b0010101010011101101: color_data = Z;
		19'b0010101010011101110: color_data = Z;
		19'b0010101010011101111: color_data = Z;
		19'b0010101010011110000: color_data = Z;
		19'b0010101010011110001: color_data = Z;
		19'b0010101010011110010: color_data = Z;
		19'b0010101010011110011: color_data = Z;
		19'b0010101010011110100: color_data = Z;
		19'b0010101010011110101: color_data = Z;
		19'b0010101010011110110: color_data = Z;
		19'b0010101010011110111: color_data = Z;
		19'b0010101010011111000: color_data = Z;
		19'b0010101010011111001: color_data = Z;
		19'b0010101010011111010: color_data = Z;
		19'b0010101010011111011: color_data = Z;
		19'b0010101010011111100: color_data = Z;
		19'b0010101010011111101: color_data = Z;
		19'b0010101010011111110: color_data = Z;
		19'b0010101010011111111: color_data = Z;
		19'b0010101010100000000: color_data = Z;
		19'b0010101010100000001: color_data = Z;
		19'b0010101010100000010: color_data = Z;
		19'b0010101010100000011: color_data = Z;
		19'b0010101010100000100: color_data = Z;
		19'b0010101010100000101: color_data = Z;
		19'b0010101010100000110: color_data = Z;
		19'b0010101010100000111: color_data = Z;
		19'b0010101010100001000: color_data = Z;
		19'b0010101010100001001: color_data = Z;
		19'b0010101010100001010: color_data = Z;
		19'b0010101010100001011: color_data = Z;
		19'b0010101010100001100: color_data = Z;
		19'b0010101010100001101: color_data = Z;
		19'b0010101010100001110: color_data = Z;
		19'b0010101010100001111: color_data = Z;
		19'b0010101010100010000: color_data = Z;
		19'b0010101010100010001: color_data = Z;
		19'b0010101010100010010: color_data = Z;
		19'b0010101010100010011: color_data = Z;
		19'b0010101010100010100: color_data = Z;
		19'b0010101010100010101: color_data = Z;
		19'b0010101010100010110: color_data = Z;
		19'b0010101010100010111: color_data = Z;
		19'b0010101010100011000: color_data = Z;
		19'b0010101010100011001: color_data = Z;
		19'b0010101010100011010: color_data = Z;
		19'b0010101010100011011: color_data = Z;
		19'b0010101010100011100: color_data = Z;
		19'b0010101010100011101: color_data = Z;
		19'b0010101010100011110: color_data = Z;
		19'b0010101010100011111: color_data = Z;
		19'b0010101010100100000: color_data = Z;
		19'b0010101010100100001: color_data = Z;
		19'b0010101010100100010: color_data = Z;
		19'b0010101010100100011: color_data = Z;
		19'b0010101010100100100: color_data = Z;
		19'b0010101010100100101: color_data = Z;
		19'b0010101010100100110: color_data = Z;
		19'b0010101010100100111: color_data = Z;
		19'b0010101010100101000: color_data = Z;
		19'b0010101010100101001: color_data = Z;
		19'b0010101010100101010: color_data = Z;
		19'b0010101010100101011: color_data = Z;
		19'b0010101010100101100: color_data = Z;
		19'b0010101010100101101: color_data = Z;
		19'b0010101010100101110: color_data = Z;
		19'b0010101010100101111: color_data = Z;
		19'b0010101010100110000: color_data = Z;
		19'b0010101010100110001: color_data = Z;
		19'b0010101010100110010: color_data = Z;
		19'b0010101010100110011: color_data = Z;
		19'b0010101010100110100: color_data = Z;
		19'b0010101010100110101: color_data = Z;
		19'b0010101010100110110: color_data = Z;
		19'b0010101010100110111: color_data = Z;
		19'b0010101010100111000: color_data = Z;
		19'b0010101010100111001: color_data = Z;
		19'b0010101010100111010: color_data = Z;
		19'b0010101010100111011: color_data = Z;
		19'b0010101010100111100: color_data = Z;
		19'b0010101010100111101: color_data = Z;
		19'b0010101010100111110: color_data = Z;
		19'b0010101010100111111: color_data = Z;
		19'b0010101010101000000: color_data = Z;
		19'b0010101010101000001: color_data = Z;
		19'b0010101010101000010: color_data = Z;
		19'b0010101010101000011: color_data = Z;
		19'b0010101010101000100: color_data = Z;
		19'b0010101010101000101: color_data = Z;
		19'b0010101010101000110: color_data = Z;
		19'b0010101010101000111: color_data = Z;
		19'b0010101010101001000: color_data = Z;
		19'b0010101010101001001: color_data = Z;
		19'b0010101010101001010: color_data = Z;
		19'b0010101010101001011: color_data = Z;
		19'b0010101010101001100: color_data = Z;
		19'b0010101010101001101: color_data = Z;
		19'b0010101010101001110: color_data = Z;
		19'b0010101010101001111: color_data = Z;
		19'b0010101010101010000: color_data = Z;
		19'b0010101010101010001: color_data = Z;
		19'b0010101010101010010: color_data = Z;
		19'b0010101010101010011: color_data = Z;
		19'b0010101010101010100: color_data = Z;
		19'b0010101010101010101: color_data = Z;
		19'b0010101010101010110: color_data = Z;
		19'b0010101010101010111: color_data = Z;
		19'b0010101010101011000: color_data = Z;
		19'b0010101010101011001: color_data = Z;
		19'b0010101010101011010: color_data = Z;
		19'b0010101010101011011: color_data = Z;
		19'b0010101010101011100: color_data = Z;
		19'b0010101010101011101: color_data = Z;
		19'b0010101010101011110: color_data = Z;
		19'b0010101010101011111: color_data = Z;
		19'b0010101010101100000: color_data = Z;
		19'b0010101010101100001: color_data = Z;
		19'b0010101010101100010: color_data = Z;
		19'b0010101010101100011: color_data = Z;
		19'b0010101010101100100: color_data = Z;
		19'b0010101010101100101: color_data = Z;
		19'b0010101010101100110: color_data = Z;
		19'b0010101010101100111: color_data = Z;
		19'b0010101010101101000: color_data = Z;
		19'b0010101010101101001: color_data = Z;
		19'b0010101010101101010: color_data = Z;
		19'b0010101010101101011: color_data = Z;
		19'b0010101010101101100: color_data = Z;
		19'b0010101010101101101: color_data = Z;
		19'b0010101010101101110: color_data = Z;
		19'b0010101010101101111: color_data = Z;
		19'b0010101010101110000: color_data = Z;
		19'b0010101010101110001: color_data = Z;
		19'b0010101010101110010: color_data = Z;
		19'b0010101010101110011: color_data = Z;
		19'b0010101010101110100: color_data = Z;
		19'b0010101010101110101: color_data = Z;
		19'b0010101010101110110: color_data = Z;
		19'b0010101010101110111: color_data = Z;
		19'b0010101010101111000: color_data = Z;
		19'b0010101010101111001: color_data = Z;
		19'b0010101010101111010: color_data = Z;
		19'b0010101010101111011: color_data = Z;
		19'b0010101010101111100: color_data = Z;
		19'b0010101010101111101: color_data = Z;
		19'b0010101010101111110: color_data = Z;
		19'b0010101010101111111: color_data = Z;
		19'b0010101010110000000: color_data = Z;
		19'b0010101010110000001: color_data = Z;
		19'b0010101010110000010: color_data = Z;
		19'b0010101010110000011: color_data = Z;
		19'b0010101010110000100: color_data = Z;
		19'b0010101010110000101: color_data = Z;
		19'b0010101010110000110: color_data = Z;
		19'b0010101010110000111: color_data = Z;
		19'b0010101010110001000: color_data = Z;
		19'b0010101010110001001: color_data = Z;
		19'b0010101010110001010: color_data = Z;
		19'b0010101010110001011: color_data = Z;
		19'b0010101010110001100: color_data = Z;
		19'b0010101010110001101: color_data = Z;
		19'b0010101010110001110: color_data = Z;
		19'b0010101010110001111: color_data = Z;
		19'b0010101010110010000: color_data = Z;
		19'b0010101010110010001: color_data = Z;
		19'b0010101010110010010: color_data = Z;
		19'b0010101010110010011: color_data = Z;
		19'b0010101010110010100: color_data = Z;
		19'b0010101010110010101: color_data = Z;
		19'b0010101010110010110: color_data = Z;
		19'b0010101010110010111: color_data = Z;
		19'b0010101010110011000: color_data = Z;
		19'b0010101010110011001: color_data = Z;
		19'b0010101010110011010: color_data = Z;
		19'b0010101010110011011: color_data = Z;
		19'b0010101010110011100: color_data = Z;
		19'b0010101010110011101: color_data = Z;
		19'b0010101010110011110: color_data = Z;
		19'b0010101010110011111: color_data = Z;
		19'b0010101010110100000: color_data = Z;
		19'b0010101010110100001: color_data = Z;
		19'b0010101010110100010: color_data = Z;
		19'b0010101010110100011: color_data = Z;
		19'b0010101010110100100: color_data = Z;
		19'b0010101010110100101: color_data = Z;
		19'b0010101010110100110: color_data = Z;
		19'b0010101010110100111: color_data = Z;
		19'b0010101010110101000: color_data = Z;
		19'b0010101010110101001: color_data = Z;
		19'b0010101010110101010: color_data = Z;
		19'b0010101010110101011: color_data = Z;
		19'b0010101010110101100: color_data = Z;
		19'b0010101010110101101: color_data = Z;
		19'b0010101010110101110: color_data = Z;
		19'b0010101010110101111: color_data = Z;
		19'b0010101010110110000: color_data = Z;
		19'b0010101010110111010: color_data = Z;
		19'b0010101010110111011: color_data = Z;
		19'b0010101010110111100: color_data = Z;
		19'b0010101010110111101: color_data = Z;
		19'b0010101010110111110: color_data = Z;
		19'b0010101010110111111: color_data = Z;
		19'b0010101010111000000: color_data = Z;
		19'b0010101010111000001: color_data = Z;
		19'b0010101010111000010: color_data = Z;
		19'b0010101010111000011: color_data = Z;
		19'b0010101010111000100: color_data = Z;
		19'b0010101010111000101: color_data = Z;
		19'b0010101010111000110: color_data = Z;
		19'b0010101010111000111: color_data = Z;
		19'b0010101010111001000: color_data = Z;
		19'b0010101010111001001: color_data = Z;
		19'b0010101010111001010: color_data = Z;
		19'b0010101010111001011: color_data = Z;
		19'b0010101100011000100: color_data = Z;
		19'b0010101100011000101: color_data = Z;
		19'b0010101100011000110: color_data = Z;
		19'b0010101100011000111: color_data = Z;
		19'b0010101100011001000: color_data = Z;
		19'b0010101100011001001: color_data = Z;
		19'b0010101100011001010: color_data = Z;
		19'b0010101100011001011: color_data = Z;
		19'b0010101100011001100: color_data = Z;
		19'b0010101100011001101: color_data = Z;
		19'b0010101100011001110: color_data = Z;
		19'b0010101100011001111: color_data = Z;
		19'b0010101100011010000: color_data = Z;
		19'b0010101100011010001: color_data = Z;
		19'b0010101100011010010: color_data = Z;
		19'b0010101100011010011: color_data = Z;
		19'b0010101100011010100: color_data = Z;
		19'b0010101100011010101: color_data = Z;
		19'b0010101100011010110: color_data = Z;
		19'b0010101100011010111: color_data = Z;
		19'b0010101100011011000: color_data = Z;
		19'b0010101100011011001: color_data = Z;
		19'b0010101100011011010: color_data = Z;
		19'b0010101100011011011: color_data = Z;
		19'b0010101100011011100: color_data = Z;
		19'b0010101100011011101: color_data = Z;
		19'b0010101100011011110: color_data = Z;
		19'b0010101100011011111: color_data = Z;
		19'b0010101100011100000: color_data = Z;
		19'b0010101100011100001: color_data = Z;
		19'b0010101100011100010: color_data = Z;
		19'b0010101100011100011: color_data = Z;
		19'b0010101100011100100: color_data = Z;
		19'b0010101100011100101: color_data = Z;
		19'b0010101100011100110: color_data = Z;
		19'b0010101100011100111: color_data = Z;
		19'b0010101100011101000: color_data = Z;
		19'b0010101100011101001: color_data = Z;
		19'b0010101100011101010: color_data = Z;
		19'b0010101100011101011: color_data = Z;
		19'b0010101100011101100: color_data = Z;
		19'b0010101100011101101: color_data = Z;
		19'b0010101100011101110: color_data = Z;
		19'b0010101100011101111: color_data = Z;
		19'b0010101100011110000: color_data = Z;
		19'b0010101100011110001: color_data = Z;
		19'b0010101100011110010: color_data = Z;
		19'b0010101100011110011: color_data = Z;
		19'b0010101100011110100: color_data = Z;
		19'b0010101100011110101: color_data = Z;
		19'b0010101100011110110: color_data = Z;
		19'b0010101100011110111: color_data = Z;
		19'b0010101100011111000: color_data = Z;
		19'b0010101100011111001: color_data = Z;
		19'b0010101100011111010: color_data = Z;
		19'b0010101100011111011: color_data = Z;
		19'b0010101100011111100: color_data = Z;
		19'b0010101100011111101: color_data = Z;
		19'b0010101100011111110: color_data = Z;
		19'b0010101100011111111: color_data = Z;
		19'b0010101100100000000: color_data = Z;
		19'b0010101100100000001: color_data = Z;
		19'b0010101100100000010: color_data = Z;
		19'b0010101100100000011: color_data = Z;
		19'b0010101100100000100: color_data = Z;
		19'b0010101100100000101: color_data = Z;
		19'b0010101100100000110: color_data = Z;
		19'b0010101100100000111: color_data = Z;
		19'b0010101100100001000: color_data = Z;
		19'b0010101100100001001: color_data = Z;
		19'b0010101100100001010: color_data = Z;
		19'b0010101100100001011: color_data = Z;
		19'b0010101100100001100: color_data = Z;
		19'b0010101100100001101: color_data = Z;
		19'b0010101100100001110: color_data = Z;
		19'b0010101100100001111: color_data = Z;
		19'b0010101100100010000: color_data = Z;
		19'b0010101100100010001: color_data = Z;
		19'b0010101100100010010: color_data = Z;
		19'b0010101100100010011: color_data = Z;
		19'b0010101100100010100: color_data = Z;
		19'b0010101100100010101: color_data = Z;
		19'b0010101100100010110: color_data = Z;
		19'b0010101100100010111: color_data = Z;
		19'b0010101100100011000: color_data = Z;
		19'b0010101100100011001: color_data = Z;
		19'b0010101100100011010: color_data = Z;
		19'b0010101100100011011: color_data = Z;
		19'b0010101100100011100: color_data = Z;
		19'b0010101100100011101: color_data = Z;
		19'b0010101100100011110: color_data = Z;
		19'b0010101100100011111: color_data = Z;
		19'b0010101100100100000: color_data = Z;
		19'b0010101100100100001: color_data = Z;
		19'b0010101100100100010: color_data = Z;
		19'b0010101100100100011: color_data = Z;
		19'b0010101100100100100: color_data = Z;
		19'b0010101100100100101: color_data = Z;
		19'b0010101100100100110: color_data = Z;
		19'b0010101100100100111: color_data = Z;
		19'b0010101100100101000: color_data = Z;
		19'b0010101100100101001: color_data = Z;
		19'b0010101100100101010: color_data = Z;
		19'b0010101100100101011: color_data = Z;
		19'b0010101100100101100: color_data = Z;
		19'b0010101100100101101: color_data = Z;
		19'b0010101100100101110: color_data = Z;
		19'b0010101100100101111: color_data = Z;
		19'b0010101100100110000: color_data = Z;
		19'b0010101100100110001: color_data = Z;
		19'b0010101100100110010: color_data = Z;
		19'b0010101100100110011: color_data = Z;
		19'b0010101100100110100: color_data = Z;
		19'b0010101100100110101: color_data = Z;
		19'b0010101100100110110: color_data = Z;
		19'b0010101100100110111: color_data = Z;
		19'b0010101100100111000: color_data = Z;
		19'b0010101100100111001: color_data = Z;
		19'b0010101100100111010: color_data = Z;
		19'b0010101100100111011: color_data = Z;
		19'b0010101100100111100: color_data = Z;
		19'b0010101100100111101: color_data = Z;
		19'b0010101100100111110: color_data = Z;
		19'b0010101100100111111: color_data = Z;
		19'b0010101100101000000: color_data = Z;
		19'b0010101100101000001: color_data = Z;
		19'b0010101100101000010: color_data = Z;
		19'b0010101100101000011: color_data = Z;
		19'b0010101100101000100: color_data = Z;
		19'b0010101100101000101: color_data = Z;
		19'b0010101100101000110: color_data = Z;
		19'b0010101100101000111: color_data = Z;
		19'b0010101100101001000: color_data = Z;
		19'b0010101100101001001: color_data = Z;
		19'b0010101100101001010: color_data = Z;
		19'b0010101100101001011: color_data = Z;
		19'b0010101100101001100: color_data = Z;
		19'b0010101100101001101: color_data = Z;
		19'b0010101100101001110: color_data = Z;
		19'b0010101100101001111: color_data = Z;
		19'b0010101100101010000: color_data = Z;
		19'b0010101100101010001: color_data = Z;
		19'b0010101100101010010: color_data = Z;
		19'b0010101100101010011: color_data = Z;
		19'b0010101100101010100: color_data = Z;
		19'b0010101100101010101: color_data = Z;
		19'b0010101100101010110: color_data = Z;
		19'b0010101100101010111: color_data = Z;
		19'b0010101100101011000: color_data = Z;
		19'b0010101100101011001: color_data = Z;
		19'b0010101100101011010: color_data = Z;
		19'b0010101100101011011: color_data = Z;
		19'b0010101100101011100: color_data = Z;
		19'b0010101100101011101: color_data = Z;
		19'b0010101100101011110: color_data = Z;
		19'b0010101100101011111: color_data = Z;
		19'b0010101100101100000: color_data = Z;
		19'b0010101100101100001: color_data = Z;
		19'b0010101100101100010: color_data = Z;
		19'b0010101100101100011: color_data = Z;
		19'b0010101100101100100: color_data = Z;
		19'b0010101100101100101: color_data = Z;
		19'b0010101100101100110: color_data = Z;
		19'b0010101100101100111: color_data = Z;
		19'b0010101100101101000: color_data = Z;
		19'b0010101100101101001: color_data = Z;
		19'b0010101100101101010: color_data = Z;
		19'b0010101100101101011: color_data = Z;
		19'b0010101100101101100: color_data = Z;
		19'b0010101100101101101: color_data = Z;
		19'b0010101100101101110: color_data = Z;
		19'b0010101100101101111: color_data = Z;
		19'b0010101100101110000: color_data = Z;
		19'b0010101100101110001: color_data = Z;
		19'b0010101100101110010: color_data = Z;
		19'b0010101100101110011: color_data = Z;
		19'b0010101100101110100: color_data = Z;
		19'b0010101100101110101: color_data = Z;
		19'b0010101100101110110: color_data = Z;
		19'b0010101100101110111: color_data = Z;
		19'b0010101100101111000: color_data = Z;
		19'b0010101100101111001: color_data = Z;
		19'b0010101100101111010: color_data = Z;
		19'b0010101100101111011: color_data = Z;
		19'b0010101100101111100: color_data = Z;
		19'b0010101100101111101: color_data = Z;
		19'b0010101100101111110: color_data = Z;
		19'b0010101100101111111: color_data = Z;
		19'b0010101100110000000: color_data = Z;
		19'b0010101100110000001: color_data = Z;
		19'b0010101100110000010: color_data = Z;
		19'b0010101100110000011: color_data = Z;
		19'b0010101100110000100: color_data = Z;
		19'b0010101100110000101: color_data = Z;
		19'b0010101100110000110: color_data = Z;
		19'b0010101100110000111: color_data = Z;
		19'b0010101100110001000: color_data = Z;
		19'b0010101100110001001: color_data = Z;
		19'b0010101100110001010: color_data = Z;
		19'b0010101100110001011: color_data = Z;
		19'b0010101100110001100: color_data = Z;
		19'b0010101100110001101: color_data = Z;
		19'b0010101100110001110: color_data = Z;
		19'b0010101100110001111: color_data = Z;
		19'b0010101100110010000: color_data = Z;
		19'b0010101100110010001: color_data = Z;
		19'b0010101100110010010: color_data = Z;
		19'b0010101100110010011: color_data = Z;
		19'b0010101100110010100: color_data = Z;
		19'b0010101100110010101: color_data = Z;
		19'b0010101100110010110: color_data = Z;
		19'b0010101100110010111: color_data = Z;
		19'b0010101100110011000: color_data = Z;
		19'b0010101100110011001: color_data = Z;
		19'b0010101100110011010: color_data = Z;
		19'b0010101100110011011: color_data = Z;
		19'b0010101100110011100: color_data = Z;
		19'b0010101100110011101: color_data = Z;
		19'b0010101100110011110: color_data = Z;
		19'b0010101100110011111: color_data = Z;
		19'b0010101100110100000: color_data = Z;
		19'b0010101100110100001: color_data = Z;
		19'b0010101100110100010: color_data = Z;
		19'b0010101100110100011: color_data = Z;
		19'b0010101100110100100: color_data = Z;
		19'b0010101100110100101: color_data = Z;
		19'b0010101100110100110: color_data = Z;
		19'b0010101100110100111: color_data = Z;
		19'b0010101100110101000: color_data = Z;
		19'b0010101100110101001: color_data = Z;
		19'b0010101100110101010: color_data = Z;
		19'b0010101100110101011: color_data = Z;
		19'b0010101100110101100: color_data = Z;
		19'b0010101100110101101: color_data = Z;
		19'b0010101100110101110: color_data = Z;
		19'b0010101100110101111: color_data = Z;
		19'b0010101100110110000: color_data = Z;
		19'b0010101100110110001: color_data = Z;
		19'b0010101100110111101: color_data = Z;
		19'b0010101100110111110: color_data = Z;
		19'b0010101100110111111: color_data = Z;
		19'b0010101100111000000: color_data = Z;
		19'b0010101100111000001: color_data = Z;
		19'b0010101100111000010: color_data = Z;
		19'b0010101100111000011: color_data = Z;
		19'b0010101100111000100: color_data = Z;
		19'b0010101100111000101: color_data = Z;
		19'b0010101100111000110: color_data = Z;
		19'b0010101100111000111: color_data = Z;
		19'b0010101100111001000: color_data = Z;
		19'b0010101100111001001: color_data = Z;
		19'b0010101100111001010: color_data = Z;
		19'b0010101100111001011: color_data = Z;
		19'b0010101100111001100: color_data = Z;
		19'b0010101110011000011: color_data = Z;
		19'b0010101110011000100: color_data = Z;
		19'b0010101110011000101: color_data = Z;
		19'b0010101110011000110: color_data = Z;
		19'b0010101110011000111: color_data = Z;
		19'b0010101110011001000: color_data = Z;
		19'b0010101110011001001: color_data = Z;
		19'b0010101110011001010: color_data = Z;
		19'b0010101110011001011: color_data = Z;
		19'b0010101110011001100: color_data = Z;
		19'b0010101110011001101: color_data = Z;
		19'b0010101110011001110: color_data = Z;
		19'b0010101110011001111: color_data = Z;
		19'b0010101110011010000: color_data = Z;
		19'b0010101110011010001: color_data = Z;
		19'b0010101110011010010: color_data = Z;
		19'b0010101110011010011: color_data = Z;
		19'b0010101110011010100: color_data = Z;
		19'b0010101110011010101: color_data = Z;
		19'b0010101110011010110: color_data = Z;
		19'b0010101110011010111: color_data = Z;
		19'b0010101110011011000: color_data = Z;
		19'b0010101110011011001: color_data = Z;
		19'b0010101110011011010: color_data = Z;
		19'b0010101110011011011: color_data = Z;
		19'b0010101110011011100: color_data = Z;
		19'b0010101110011011101: color_data = Z;
		19'b0010101110011011110: color_data = Z;
		19'b0010101110011011111: color_data = Z;
		19'b0010101110011100000: color_data = Z;
		19'b0010101110011100001: color_data = Z;
		19'b0010101110011100010: color_data = Z;
		19'b0010101110011100011: color_data = Z;
		19'b0010101110011100100: color_data = Z;
		19'b0010101110011100101: color_data = Z;
		19'b0010101110011100110: color_data = Z;
		19'b0010101110011100111: color_data = Z;
		19'b0010101110011101000: color_data = Z;
		19'b0010101110011101001: color_data = Z;
		19'b0010101110011101010: color_data = Z;
		19'b0010101110011101011: color_data = Z;
		19'b0010101110011101100: color_data = Z;
		19'b0010101110011101101: color_data = Z;
		19'b0010101110011101110: color_data = Z;
		19'b0010101110011101111: color_data = Z;
		19'b0010101110011110000: color_data = Z;
		19'b0010101110011110001: color_data = Z;
		19'b0010101110011110010: color_data = Z;
		19'b0010101110011110011: color_data = Z;
		19'b0010101110011110100: color_data = Z;
		19'b0010101110011110101: color_data = Z;
		19'b0010101110011110110: color_data = Z;
		19'b0010101110011110111: color_data = Z;
		19'b0010101110011111000: color_data = Z;
		19'b0010101110011111001: color_data = Z;
		19'b0010101110011111010: color_data = Z;
		19'b0010101110011111011: color_data = Z;
		19'b0010101110011111100: color_data = Z;
		19'b0010101110011111101: color_data = Z;
		19'b0010101110011111110: color_data = Z;
		19'b0010101110011111111: color_data = Z;
		19'b0010101110100000000: color_data = Z;
		19'b0010101110100000001: color_data = Z;
		19'b0010101110100000010: color_data = Z;
		19'b0010101110100000011: color_data = Z;
		19'b0010101110100000100: color_data = Z;
		19'b0010101110100000101: color_data = Z;
		19'b0010101110100000110: color_data = Z;
		19'b0010101110100000111: color_data = Z;
		19'b0010101110100001000: color_data = Z;
		19'b0010101110100001001: color_data = Z;
		19'b0010101110100001010: color_data = Z;
		19'b0010101110100001011: color_data = Z;
		19'b0010101110100001100: color_data = Z;
		19'b0010101110100001101: color_data = Z;
		19'b0010101110100001110: color_data = Z;
		19'b0010101110100001111: color_data = Z;
		19'b0010101110100010000: color_data = Z;
		19'b0010101110100010001: color_data = Z;
		19'b0010101110100010010: color_data = Z;
		19'b0010101110100010011: color_data = Z;
		19'b0010101110100010100: color_data = Z;
		19'b0010101110100010101: color_data = Z;
		19'b0010101110100010110: color_data = Z;
		19'b0010101110100010111: color_data = Z;
		19'b0010101110100011000: color_data = Z;
		19'b0010101110100011001: color_data = Z;
		19'b0010101110100011010: color_data = Z;
		19'b0010101110100011011: color_data = Z;
		19'b0010101110100011100: color_data = Z;
		19'b0010101110100011101: color_data = Z;
		19'b0010101110100011110: color_data = Z;
		19'b0010101110100011111: color_data = Z;
		19'b0010101110100100000: color_data = Z;
		19'b0010101110100100001: color_data = Z;
		19'b0010101110100100010: color_data = Z;
		19'b0010101110100100011: color_data = Z;
		19'b0010101110100100100: color_data = Z;
		19'b0010101110100100101: color_data = Z;
		19'b0010101110100100110: color_data = Z;
		19'b0010101110100100111: color_data = Z;
		19'b0010101110100101000: color_data = Z;
		19'b0010101110100101001: color_data = Z;
		19'b0010101110100101010: color_data = Z;
		19'b0010101110100101011: color_data = Z;
		19'b0010101110100101100: color_data = Z;
		19'b0010101110100101101: color_data = Z;
		19'b0010101110100101110: color_data = Z;
		19'b0010101110100101111: color_data = Z;
		19'b0010101110100110000: color_data = Z;
		19'b0010101110100110001: color_data = Z;
		19'b0010101110100110010: color_data = Z;
		19'b0010101110100110011: color_data = Z;
		19'b0010101110100110100: color_data = Z;
		19'b0010101110100110101: color_data = Z;
		19'b0010101110100110110: color_data = Z;
		19'b0010101110100110111: color_data = Z;
		19'b0010101110100111000: color_data = Z;
		19'b0010101110100111001: color_data = Z;
		19'b0010101110100111010: color_data = Z;
		19'b0010101110100111011: color_data = Z;
		19'b0010101110100111100: color_data = Z;
		19'b0010101110100111101: color_data = Z;
		19'b0010101110100111110: color_data = Z;
		19'b0010101110100111111: color_data = Z;
		19'b0010101110101000000: color_data = Z;
		19'b0010101110101000001: color_data = Z;
		19'b0010101110101000010: color_data = Z;
		19'b0010101110101000011: color_data = Z;
		19'b0010101110101000100: color_data = Z;
		19'b0010101110101000101: color_data = Z;
		19'b0010101110101000110: color_data = Z;
		19'b0010101110101000111: color_data = Z;
		19'b0010101110101001000: color_data = Z;
		19'b0010101110101001001: color_data = Z;
		19'b0010101110101001010: color_data = Z;
		19'b0010101110101001011: color_data = Z;
		19'b0010101110101001100: color_data = Z;
		19'b0010101110101001101: color_data = Z;
		19'b0010101110101001110: color_data = Z;
		19'b0010101110101001111: color_data = Z;
		19'b0010101110101010000: color_data = Z;
		19'b0010101110101010001: color_data = Z;
		19'b0010101110101010010: color_data = Z;
		19'b0010101110101010011: color_data = Z;
		19'b0010101110101010100: color_data = Z;
		19'b0010101110101010101: color_data = Z;
		19'b0010101110101010110: color_data = Z;
		19'b0010101110101010111: color_data = Z;
		19'b0010101110101011000: color_data = Z;
		19'b0010101110101011001: color_data = Z;
		19'b0010101110101011010: color_data = Z;
		19'b0010101110101011011: color_data = Z;
		19'b0010101110101011100: color_data = Z;
		19'b0010101110101011101: color_data = Z;
		19'b0010101110101011110: color_data = Z;
		19'b0010101110101011111: color_data = Z;
		19'b0010101110101100000: color_data = Z;
		19'b0010101110101100001: color_data = Z;
		19'b0010101110101100010: color_data = Z;
		19'b0010101110101100011: color_data = Z;
		19'b0010101110101100100: color_data = Z;
		19'b0010101110101100101: color_data = Z;
		19'b0010101110101100110: color_data = Z;
		19'b0010101110101100111: color_data = Z;
		19'b0010101110101101000: color_data = Z;
		19'b0010101110101101001: color_data = Z;
		19'b0010101110101101010: color_data = Z;
		19'b0010101110101101011: color_data = Z;
		19'b0010101110101101100: color_data = Z;
		19'b0010101110101101101: color_data = Z;
		19'b0010101110101101110: color_data = Z;
		19'b0010101110101101111: color_data = Z;
		19'b0010101110101110000: color_data = Z;
		19'b0010101110101110001: color_data = Z;
		19'b0010101110101110010: color_data = Z;
		19'b0010101110101110011: color_data = Z;
		19'b0010101110101110100: color_data = Z;
		19'b0010101110101110101: color_data = Z;
		19'b0010101110101110110: color_data = Z;
		19'b0010101110101110111: color_data = Z;
		19'b0010101110101111000: color_data = Z;
		19'b0010101110101111001: color_data = Z;
		19'b0010101110101111010: color_data = Z;
		19'b0010101110101111011: color_data = Z;
		19'b0010101110101111100: color_data = Z;
		19'b0010101110101111101: color_data = Z;
		19'b0010101110101111110: color_data = Z;
		19'b0010101110101111111: color_data = Z;
		19'b0010101110110000000: color_data = Z;
		19'b0010101110110000001: color_data = Z;
		19'b0010101110110000010: color_data = Z;
		19'b0010101110110000011: color_data = Z;
		19'b0010101110110000100: color_data = Z;
		19'b0010101110110000101: color_data = Z;
		19'b0010101110110000110: color_data = Z;
		19'b0010101110110000111: color_data = Z;
		19'b0010101110110001000: color_data = Z;
		19'b0010101110110001001: color_data = Z;
		19'b0010101110110001010: color_data = Z;
		19'b0010101110110001011: color_data = Z;
		19'b0010101110110001100: color_data = Z;
		19'b0010101110110001101: color_data = Z;
		19'b0010101110110001110: color_data = Z;
		19'b0010101110110001111: color_data = Z;
		19'b0010101110110010000: color_data = Z;
		19'b0010101110110010001: color_data = Z;
		19'b0010101110110010010: color_data = Z;
		19'b0010101110110010011: color_data = Z;
		19'b0010101110110010100: color_data = Z;
		19'b0010101110110010101: color_data = Z;
		19'b0010101110110010110: color_data = Z;
		19'b0010101110110010111: color_data = Z;
		19'b0010101110110011000: color_data = Z;
		19'b0010101110110011001: color_data = Z;
		19'b0010101110110011010: color_data = Z;
		19'b0010101110110011011: color_data = Z;
		19'b0010101110110011100: color_data = Z;
		19'b0010101110110011101: color_data = Z;
		19'b0010101110110011110: color_data = Z;
		19'b0010101110110011111: color_data = Z;
		19'b0010101110110100000: color_data = Z;
		19'b0010101110110100001: color_data = Z;
		19'b0010101110110100010: color_data = Z;
		19'b0010101110110100011: color_data = Z;
		19'b0010101110110100100: color_data = Z;
		19'b0010101110110100101: color_data = Z;
		19'b0010101110110100110: color_data = Z;
		19'b0010101110110100111: color_data = Z;
		19'b0010101110110101000: color_data = Z;
		19'b0010101110110101001: color_data = Z;
		19'b0010101110110101010: color_data = Z;
		19'b0010101110110101011: color_data = Z;
		19'b0010101110110101100: color_data = Z;
		19'b0010101110110101101: color_data = Z;
		19'b0010101110110101110: color_data = Z;
		19'b0010101110110101111: color_data = Z;
		19'b0010101110110110000: color_data = Z;
		19'b0010101110110110001: color_data = Z;
		19'b0010101110110111111: color_data = Z;
		19'b0010101110111000000: color_data = Z;
		19'b0010101110111000001: color_data = Z;
		19'b0010101110111000010: color_data = Z;
		19'b0010101110111000011: color_data = Z;
		19'b0010101110111000100: color_data = Z;
		19'b0010101110111000101: color_data = Z;
		19'b0010101110111000110: color_data = Z;
		19'b0010101110111000111: color_data = Z;
		19'b0010101110111001000: color_data = Z;
		19'b0010101110111001001: color_data = Z;
		19'b0010101110111001010: color_data = Z;
		19'b0010101110111001011: color_data = Z;
		19'b0010101110111001100: color_data = Z;
		19'b0010110000011000010: color_data = Z;
		19'b0010110000011000011: color_data = Z;
		19'b0010110000011000100: color_data = Z;
		19'b0010110000011000101: color_data = Z;
		19'b0010110000011000110: color_data = Z;
		19'b0010110000011000111: color_data = Z;
		19'b0010110000011001000: color_data = Z;
		19'b0010110000011001001: color_data = Z;
		19'b0010110000011001010: color_data = Z;
		19'b0010110000011001011: color_data = Z;
		19'b0010110000011001100: color_data = Z;
		19'b0010110000011001101: color_data = Z;
		19'b0010110000011001110: color_data = Z;
		19'b0010110000011001111: color_data = Z;
		19'b0010110000011010000: color_data = Z;
		19'b0010110000011010001: color_data = Z;
		19'b0010110000011010010: color_data = Z;
		19'b0010110000011010011: color_data = Z;
		19'b0010110000011010100: color_data = Z;
		19'b0010110000011010101: color_data = Z;
		19'b0010110000011010110: color_data = Z;
		19'b0010110000011010111: color_data = Z;
		19'b0010110000011011000: color_data = Z;
		19'b0010110000011011001: color_data = Z;
		19'b0010110000011011010: color_data = Z;
		19'b0010110000011011011: color_data = Z;
		19'b0010110000011011100: color_data = Z;
		19'b0010110000011011101: color_data = Z;
		19'b0010110000011011110: color_data = Z;
		19'b0010110000011011111: color_data = Z;
		19'b0010110000011100000: color_data = Z;
		19'b0010110000011100001: color_data = Z;
		19'b0010110000011100010: color_data = Z;
		19'b0010110000011100011: color_data = Z;
		19'b0010110000011100100: color_data = Z;
		19'b0010110000011100101: color_data = Z;
		19'b0010110000011100110: color_data = Z;
		19'b0010110000011100111: color_data = Z;
		19'b0010110000011101000: color_data = Z;
		19'b0010110000011101001: color_data = Z;
		19'b0010110000011101010: color_data = Z;
		19'b0010110000011101011: color_data = Z;
		19'b0010110000011101100: color_data = Z;
		19'b0010110000011101101: color_data = Z;
		19'b0010110000011101110: color_data = Z;
		19'b0010110000011101111: color_data = Z;
		19'b0010110000011110000: color_data = Z;
		19'b0010110000011110001: color_data = Z;
		19'b0010110000011110010: color_data = Z;
		19'b0010110000011110011: color_data = Z;
		19'b0010110000011110100: color_data = Z;
		19'b0010110000011110101: color_data = Z;
		19'b0010110000011110110: color_data = Z;
		19'b0010110000011110111: color_data = Z;
		19'b0010110000011111000: color_data = Z;
		19'b0010110000011111001: color_data = Z;
		19'b0010110000011111010: color_data = Z;
		19'b0010110000011111011: color_data = Z;
		19'b0010110000011111100: color_data = Z;
		19'b0010110000011111101: color_data = Z;
		19'b0010110000011111110: color_data = Z;
		19'b0010110000011111111: color_data = Z;
		19'b0010110000100000000: color_data = Z;
		19'b0010110000100000001: color_data = Z;
		19'b0010110000100000010: color_data = Z;
		19'b0010110000100000011: color_data = Z;
		19'b0010110000100000100: color_data = Z;
		19'b0010110000100000101: color_data = Z;
		19'b0010110000100000110: color_data = Z;
		19'b0010110000100000111: color_data = Z;
		19'b0010110000100001000: color_data = Z;
		19'b0010110000100001001: color_data = Z;
		19'b0010110000100001010: color_data = Z;
		19'b0010110000100001011: color_data = Z;
		19'b0010110000100001100: color_data = Z;
		19'b0010110000100001101: color_data = Z;
		19'b0010110000100001110: color_data = Z;
		19'b0010110000100001111: color_data = Z;
		19'b0010110000100010000: color_data = Z;
		19'b0010110000100010001: color_data = Z;
		19'b0010110000100010010: color_data = Z;
		19'b0010110000100010011: color_data = Z;
		19'b0010110000100010100: color_data = Z;
		19'b0010110000100010101: color_data = Z;
		19'b0010110000100010110: color_data = Z;
		19'b0010110000100010111: color_data = Z;
		19'b0010110000100011000: color_data = Z;
		19'b0010110000100011001: color_data = Z;
		19'b0010110000100011010: color_data = Z;
		19'b0010110000100011011: color_data = Z;
		19'b0010110000100011100: color_data = Z;
		19'b0010110000100011101: color_data = Z;
		19'b0010110000100011110: color_data = Z;
		19'b0010110000100011111: color_data = Z;
		19'b0010110000100100000: color_data = Z;
		19'b0010110000100100001: color_data = Z;
		19'b0010110000100100010: color_data = Z;
		19'b0010110000100100011: color_data = Z;
		19'b0010110000100100100: color_data = Z;
		19'b0010110000100100101: color_data = Z;
		19'b0010110000100100110: color_data = Z;
		19'b0010110000100100111: color_data = Z;
		19'b0010110000100101000: color_data = Z;
		19'b0010110000100101001: color_data = Z;
		19'b0010110000100101010: color_data = Z;
		19'b0010110000100101011: color_data = Z;
		19'b0010110000100101100: color_data = Z;
		19'b0010110000100101101: color_data = Z;
		19'b0010110000100101110: color_data = Z;
		19'b0010110000100101111: color_data = Z;
		19'b0010110000100110000: color_data = Z;
		19'b0010110000100110001: color_data = Z;
		19'b0010110000100110010: color_data = Z;
		19'b0010110000100110011: color_data = Z;
		19'b0010110000100110100: color_data = Z;
		19'b0010110000100110101: color_data = Z;
		19'b0010110000100110110: color_data = Z;
		19'b0010110000100110111: color_data = Z;
		19'b0010110000100111000: color_data = Z;
		19'b0010110000100111001: color_data = Z;
		19'b0010110000100111010: color_data = Z;
		19'b0010110000100111011: color_data = Z;
		19'b0010110000100111100: color_data = Z;
		19'b0010110000100111101: color_data = Z;
		19'b0010110000100111110: color_data = Z;
		19'b0010110000100111111: color_data = Z;
		19'b0010110000101000000: color_data = Z;
		19'b0010110000101000001: color_data = Z;
		19'b0010110000101000010: color_data = Z;
		19'b0010110000101000011: color_data = Z;
		19'b0010110000101000100: color_data = Z;
		19'b0010110000101000101: color_data = Z;
		19'b0010110000101000110: color_data = Z;
		19'b0010110000101000111: color_data = Z;
		19'b0010110000101001000: color_data = Z;
		19'b0010110000101001001: color_data = Z;
		19'b0010110000101001010: color_data = Z;
		19'b0010110000101001011: color_data = Z;
		19'b0010110000101001100: color_data = Z;
		19'b0010110000101001101: color_data = Z;
		19'b0010110000101001110: color_data = Z;
		19'b0010110000101001111: color_data = Z;
		19'b0010110000101010000: color_data = Z;
		19'b0010110000101010001: color_data = Z;
		19'b0010110000101010010: color_data = Z;
		19'b0010110000101010011: color_data = Z;
		19'b0010110000101010100: color_data = Z;
		19'b0010110000101010101: color_data = Z;
		19'b0010110000101010110: color_data = Z;
		19'b0010110000101010111: color_data = Z;
		19'b0010110000101011000: color_data = Z;
		19'b0010110000101011001: color_data = Z;
		19'b0010110000101011010: color_data = Z;
		19'b0010110000101011011: color_data = Z;
		19'b0010110000101011100: color_data = Z;
		19'b0010110000101011101: color_data = Z;
		19'b0010110000101011110: color_data = Z;
		19'b0010110000101011111: color_data = Z;
		19'b0010110000101100000: color_data = Z;
		19'b0010110000101100001: color_data = Z;
		19'b0010110000101100010: color_data = Z;
		19'b0010110000101100011: color_data = Z;
		19'b0010110000101100100: color_data = Z;
		19'b0010110000101100101: color_data = Z;
		19'b0010110000101100110: color_data = Z;
		19'b0010110000101100111: color_data = Z;
		19'b0010110000101101000: color_data = Z;
		19'b0010110000101101001: color_data = Z;
		19'b0010110000101101010: color_data = Z;
		19'b0010110000101101011: color_data = Z;
		19'b0010110000101101100: color_data = Z;
		19'b0010110000101101101: color_data = Z;
		19'b0010110000101101110: color_data = Z;
		19'b0010110000101101111: color_data = Z;
		19'b0010110000101110000: color_data = Z;
		19'b0010110000101110001: color_data = Z;
		19'b0010110000101110010: color_data = Z;
		19'b0010110000101110011: color_data = Z;
		19'b0010110000101110100: color_data = Z;
		19'b0010110000101110101: color_data = Z;
		19'b0010110000101110110: color_data = Z;
		19'b0010110000101110111: color_data = Z;
		19'b0010110000101111000: color_data = Z;
		19'b0010110000101111001: color_data = Z;
		19'b0010110000101111010: color_data = Z;
		19'b0010110000101111011: color_data = Z;
		19'b0010110000101111100: color_data = Z;
		19'b0010110000101111101: color_data = Z;
		19'b0010110000101111110: color_data = Z;
		19'b0010110000101111111: color_data = Z;
		19'b0010110000110000000: color_data = Z;
		19'b0010110000110000001: color_data = Z;
		19'b0010110000110000010: color_data = Z;
		19'b0010110000110000011: color_data = Z;
		19'b0010110000110000100: color_data = Z;
		19'b0010110000110000101: color_data = Z;
		19'b0010110000110000110: color_data = Z;
		19'b0010110000110000111: color_data = Z;
		19'b0010110000110001000: color_data = Z;
		19'b0010110000110001001: color_data = Z;
		19'b0010110000110001010: color_data = Z;
		19'b0010110000110001011: color_data = Z;
		19'b0010110000110001100: color_data = Z;
		19'b0010110000110001101: color_data = Z;
		19'b0010110000110001110: color_data = Z;
		19'b0010110000110001111: color_data = Z;
		19'b0010110000110010000: color_data = Z;
		19'b0010110000110010001: color_data = Z;
		19'b0010110000110010010: color_data = Z;
		19'b0010110000110010011: color_data = Z;
		19'b0010110000110010100: color_data = Z;
		19'b0010110000110010101: color_data = Z;
		19'b0010110000110010110: color_data = Z;
		19'b0010110000110010111: color_data = Z;
		19'b0010110000110011000: color_data = Z;
		19'b0010110000110011001: color_data = Z;
		19'b0010110000110011010: color_data = Z;
		19'b0010110000110011011: color_data = Z;
		19'b0010110000110011100: color_data = Z;
		19'b0010110000110011101: color_data = Z;
		19'b0010110000110011110: color_data = Z;
		19'b0010110000110011111: color_data = Z;
		19'b0010110000110100000: color_data = Z;
		19'b0010110000110100001: color_data = Z;
		19'b0010110000110100010: color_data = Z;
		19'b0010110000110100011: color_data = Z;
		19'b0010110000110100100: color_data = Z;
		19'b0010110000110100101: color_data = Z;
		19'b0010110000110100110: color_data = Z;
		19'b0010110000110100111: color_data = Z;
		19'b0010110000110101000: color_data = Z;
		19'b0010110000110101001: color_data = Z;
		19'b0010110000110101010: color_data = Z;
		19'b0010110000110101011: color_data = Z;
		19'b0010110000110101100: color_data = Z;
		19'b0010110000110101101: color_data = Z;
		19'b0010110000110101110: color_data = Z;
		19'b0010110000110101111: color_data = Z;
		19'b0010110000110110000: color_data = Z;
		19'b0010110000110110001: color_data = Z;
		19'b0010110000110111011: color_data = Z;
		19'b0010110000110111100: color_data = Z;
		19'b0010110000110111101: color_data = Z;
		19'b0010110000110111110: color_data = Z;
		19'b0010110000110111111: color_data = Z;
		19'b0010110000111000001: color_data = Z;
		19'b0010110000111000010: color_data = Z;
		19'b0010110000111000011: color_data = Z;
		19'b0010110000111000100: color_data = Z;
		19'b0010110000111000101: color_data = Z;
		19'b0010110000111000110: color_data = Z;
		19'b0010110000111000111: color_data = Z;
		19'b0010110000111001000: color_data = Z;
		19'b0010110000111001001: color_data = Z;
		19'b0010110000111001010: color_data = Z;
		19'b0010110000111001011: color_data = Z;
		19'b0010110000111001100: color_data = Z;
		19'b0010110010011000001: color_data = Z;
		19'b0010110010011000010: color_data = Z;
		19'b0010110010011000011: color_data = Z;
		19'b0010110010011000100: color_data = Z;
		19'b0010110010011000101: color_data = Z;
		19'b0010110010011000110: color_data = Z;
		19'b0010110010011000111: color_data = Z;
		19'b0010110010011001000: color_data = Z;
		19'b0010110010011001001: color_data = Z;
		19'b0010110010011001010: color_data = Z;
		19'b0010110010011001011: color_data = Z;
		19'b0010110010011001100: color_data = Z;
		19'b0010110010011001101: color_data = Z;
		19'b0010110010011001110: color_data = Z;
		19'b0010110010011001111: color_data = Z;
		19'b0010110010011010000: color_data = Z;
		19'b0010110010011010001: color_data = Z;
		19'b0010110010011010010: color_data = Z;
		19'b0010110010011010011: color_data = Z;
		19'b0010110010011010100: color_data = Z;
		19'b0010110010011010101: color_data = Z;
		19'b0010110010011010110: color_data = Z;
		19'b0010110010011010111: color_data = Z;
		19'b0010110010011011000: color_data = Z;
		19'b0010110010011011001: color_data = Z;
		19'b0010110010011011010: color_data = Z;
		19'b0010110010011011011: color_data = Z;
		19'b0010110010011011100: color_data = Z;
		19'b0010110010011011101: color_data = Z;
		19'b0010110010011011110: color_data = Z;
		19'b0010110010011011111: color_data = Z;
		19'b0010110010011100000: color_data = Z;
		19'b0010110010011100001: color_data = Z;
		19'b0010110010011100010: color_data = Z;
		19'b0010110010011100011: color_data = Z;
		19'b0010110010011100100: color_data = Z;
		19'b0010110010011100101: color_data = Z;
		19'b0010110010011100110: color_data = Z;
		19'b0010110010011100111: color_data = Z;
		19'b0010110010011101000: color_data = Z;
		19'b0010110010011101001: color_data = Z;
		19'b0010110010011101010: color_data = Z;
		19'b0010110010011101011: color_data = Z;
		19'b0010110010011101100: color_data = Z;
		19'b0010110010011101101: color_data = Z;
		19'b0010110010011101110: color_data = Z;
		19'b0010110010011101111: color_data = Z;
		19'b0010110010011110000: color_data = Z;
		19'b0010110010011110001: color_data = Z;
		19'b0010110010011110010: color_data = Z;
		19'b0010110010011110011: color_data = Z;
		19'b0010110010011110100: color_data = Z;
		19'b0010110010011110101: color_data = Z;
		19'b0010110010011110110: color_data = Z;
		19'b0010110010011110111: color_data = Z;
		19'b0010110010011111000: color_data = Z;
		19'b0010110010011111001: color_data = Z;
		19'b0010110010011111010: color_data = Z;
		19'b0010110010011111011: color_data = Z;
		19'b0010110010011111100: color_data = Z;
		19'b0010110010011111101: color_data = Z;
		19'b0010110010011111110: color_data = Z;
		19'b0010110010011111111: color_data = Z;
		19'b0010110010100000000: color_data = Z;
		19'b0010110010100000001: color_data = Z;
		19'b0010110010100000010: color_data = Z;
		19'b0010110010100000011: color_data = Z;
		19'b0010110010100000100: color_data = Z;
		19'b0010110010100000101: color_data = Z;
		19'b0010110010100000110: color_data = Z;
		19'b0010110010100000111: color_data = Z;
		19'b0010110010100001000: color_data = Z;
		19'b0010110010100001001: color_data = Z;
		19'b0010110010100001010: color_data = Z;
		19'b0010110010100001011: color_data = Z;
		19'b0010110010100001100: color_data = Z;
		19'b0010110010100001101: color_data = Z;
		19'b0010110010100001110: color_data = Z;
		19'b0010110010100001111: color_data = Z;
		19'b0010110010100010000: color_data = Z;
		19'b0010110010100010001: color_data = Z;
		19'b0010110010100010010: color_data = Z;
		19'b0010110010100010011: color_data = Z;
		19'b0010110010100010100: color_data = Z;
		19'b0010110010100010101: color_data = Z;
		19'b0010110010100010110: color_data = Z;
		19'b0010110010100010111: color_data = Z;
		19'b0010110010100011000: color_data = Z;
		19'b0010110010100011001: color_data = Z;
		19'b0010110010100011010: color_data = Z;
		19'b0010110010100011011: color_data = Z;
		19'b0010110010100011100: color_data = Z;
		19'b0010110010100011101: color_data = Z;
		19'b0010110010100011110: color_data = Z;
		19'b0010110010100011111: color_data = Z;
		19'b0010110010100100000: color_data = Z;
		19'b0010110010100100001: color_data = Z;
		19'b0010110010100100010: color_data = Z;
		19'b0010110010100100011: color_data = Z;
		19'b0010110010100100100: color_data = Z;
		19'b0010110010100100101: color_data = Z;
		19'b0010110010100100110: color_data = Z;
		19'b0010110010100100111: color_data = Z;
		19'b0010110010100101000: color_data = Z;
		19'b0010110010100101001: color_data = Z;
		19'b0010110010100101010: color_data = Z;
		19'b0010110010100101011: color_data = Z;
		19'b0010110010100101100: color_data = Z;
		19'b0010110010100101101: color_data = Z;
		19'b0010110010100101110: color_data = Z;
		19'b0010110010100101111: color_data = Z;
		19'b0010110010100110000: color_data = Z;
		19'b0010110010100110001: color_data = Z;
		19'b0010110010100110010: color_data = Z;
		19'b0010110010100110011: color_data = Z;
		19'b0010110010100110100: color_data = Z;
		19'b0010110010100110101: color_data = Z;
		19'b0010110010100110110: color_data = Z;
		19'b0010110010100110111: color_data = Z;
		19'b0010110010100111000: color_data = Z;
		19'b0010110010100111001: color_data = Z;
		19'b0010110010100111010: color_data = Z;
		19'b0010110010100111011: color_data = Z;
		19'b0010110010100111100: color_data = Z;
		19'b0010110010100111101: color_data = Z;
		19'b0010110010100111110: color_data = Z;
		19'b0010110010100111111: color_data = Z;
		19'b0010110010101000000: color_data = Z;
		19'b0010110010101000001: color_data = Z;
		19'b0010110010101000010: color_data = Z;
		19'b0010110010101000011: color_data = Z;
		19'b0010110010101000100: color_data = Z;
		19'b0010110010101000101: color_data = Z;
		19'b0010110010101000110: color_data = Z;
		19'b0010110010101000111: color_data = Z;
		19'b0010110010101001000: color_data = Z;
		19'b0010110010101001001: color_data = Z;
		19'b0010110010101001010: color_data = Z;
		19'b0010110010101001011: color_data = Z;
		19'b0010110010101001100: color_data = Z;
		19'b0010110010101001101: color_data = Z;
		19'b0010110010101001110: color_data = Z;
		19'b0010110010101001111: color_data = Z;
		19'b0010110010101010000: color_data = Z;
		19'b0010110010101010001: color_data = Z;
		19'b0010110010101010010: color_data = Z;
		19'b0010110010101010011: color_data = Z;
		19'b0010110010101010100: color_data = Z;
		19'b0010110010101010101: color_data = Z;
		19'b0010110010101010110: color_data = Z;
		19'b0010110010101010111: color_data = Z;
		19'b0010110010101011000: color_data = Z;
		19'b0010110010101011001: color_data = Z;
		19'b0010110010101011010: color_data = Z;
		19'b0010110010101011011: color_data = Z;
		19'b0010110010101011100: color_data = Z;
		19'b0010110010101011101: color_data = Z;
		19'b0010110010101011110: color_data = Z;
		19'b0010110010101011111: color_data = Z;
		19'b0010110010101100000: color_data = Z;
		19'b0010110010101100001: color_data = Z;
		19'b0010110010101100010: color_data = Z;
		19'b0010110010101100011: color_data = Z;
		19'b0010110010101100100: color_data = Z;
		19'b0010110010101100101: color_data = Z;
		19'b0010110010101100110: color_data = Z;
		19'b0010110010101100111: color_data = Z;
		19'b0010110010101101000: color_data = Z;
		19'b0010110010101101001: color_data = Z;
		19'b0010110010101101010: color_data = Z;
		19'b0010110010101101011: color_data = Z;
		19'b0010110010101101100: color_data = Z;
		19'b0010110010101101101: color_data = Z;
		19'b0010110010101101110: color_data = Z;
		19'b0010110010101101111: color_data = Z;
		19'b0010110010101110000: color_data = Z;
		19'b0010110010101110001: color_data = Z;
		19'b0010110010101110010: color_data = Z;
		19'b0010110010101110011: color_data = Z;
		19'b0010110010101110100: color_data = Z;
		19'b0010110010101110101: color_data = Z;
		19'b0010110010101110110: color_data = Z;
		19'b0010110010101110111: color_data = Z;
		19'b0010110010101111000: color_data = Z;
		19'b0010110010101111001: color_data = Z;
		19'b0010110010101111010: color_data = Z;
		19'b0010110010101111011: color_data = Z;
		19'b0010110010101111100: color_data = Z;
		19'b0010110010101111101: color_data = Z;
		19'b0010110010101111110: color_data = Z;
		19'b0010110010101111111: color_data = Z;
		19'b0010110010110000000: color_data = Z;
		19'b0010110010110000001: color_data = Z;
		19'b0010110010110000010: color_data = Z;
		19'b0010110010110000011: color_data = Z;
		19'b0010110010110000100: color_data = Z;
		19'b0010110010110000101: color_data = Z;
		19'b0010110010110000110: color_data = Z;
		19'b0010110010110000111: color_data = Z;
		19'b0010110010110001000: color_data = Z;
		19'b0010110010110001001: color_data = Z;
		19'b0010110010110001010: color_data = Z;
		19'b0010110010110001011: color_data = Z;
		19'b0010110010110001100: color_data = Z;
		19'b0010110010110001101: color_data = Z;
		19'b0010110010110001110: color_data = Z;
		19'b0010110010110001111: color_data = Z;
		19'b0010110010110010000: color_data = Z;
		19'b0010110010110010001: color_data = Z;
		19'b0010110010110010010: color_data = Z;
		19'b0010110010110010011: color_data = Z;
		19'b0010110010110010100: color_data = Z;
		19'b0010110010110010101: color_data = Z;
		19'b0010110010110010110: color_data = Z;
		19'b0010110010110010111: color_data = Z;
		19'b0010110010110011000: color_data = Z;
		19'b0010110010110011001: color_data = Z;
		19'b0010110010110011010: color_data = Z;
		19'b0010110010110011011: color_data = Z;
		19'b0010110010110011100: color_data = Z;
		19'b0010110010110011101: color_data = Z;
		19'b0010110010110011110: color_data = Z;
		19'b0010110010110011111: color_data = Z;
		19'b0010110010110100000: color_data = Z;
		19'b0010110010110100001: color_data = Z;
		19'b0010110010110100010: color_data = Z;
		19'b0010110010110100011: color_data = Z;
		19'b0010110010110100100: color_data = Z;
		19'b0010110010110100101: color_data = Z;
		19'b0010110010110100110: color_data = Z;
		19'b0010110010110100111: color_data = Z;
		19'b0010110010110101000: color_data = Z;
		19'b0010110010110101001: color_data = Z;
		19'b0010110010110101010: color_data = Z;
		19'b0010110010110101011: color_data = Z;
		19'b0010110010110101100: color_data = Z;
		19'b0010110010110101101: color_data = Z;
		19'b0010110010110101110: color_data = Z;
		19'b0010110010110101111: color_data = Z;
		19'b0010110010110110000: color_data = Z;
		19'b0010110010110110001: color_data = Z;
		19'b0010110010110110010: color_data = Z;
		19'b0010110010110111011: color_data = Z;
		19'b0010110010110111100: color_data = Z;
		19'b0010110010111000001: color_data = Z;
		19'b0010110010111000010: color_data = Z;
		19'b0010110010111000011: color_data = Z;
		19'b0010110010111000100: color_data = Z;
		19'b0010110010111000101: color_data = Z;
		19'b0010110010111000110: color_data = Z;
		19'b0010110010111000111: color_data = Z;
		19'b0010110010111001000: color_data = Z;
		19'b0010110010111001001: color_data = Z;
		19'b0010110010111001010: color_data = Z;
		19'b0010110010111001011: color_data = Z;
		19'b0010110010111001100: color_data = Z;
		19'b0010110010111001101: color_data = Z;
		19'b0010110100011000001: color_data = Z;
		19'b0010110100011000010: color_data = Z;
		19'b0010110100011000011: color_data = Z;
		19'b0010110100011000100: color_data = Z;
		19'b0010110100011000101: color_data = Z;
		19'b0010110100011000110: color_data = Z;
		19'b0010110100011000111: color_data = Z;
		19'b0010110100011001000: color_data = Z;
		19'b0010110100011001001: color_data = Z;
		19'b0010110100011001010: color_data = Z;
		19'b0010110100011001011: color_data = Z;
		19'b0010110100011001100: color_data = Z;
		19'b0010110100011001101: color_data = Z;
		19'b0010110100011001110: color_data = Z;
		19'b0010110100011001111: color_data = Z;
		19'b0010110100011010000: color_data = Z;
		19'b0010110100011010001: color_data = Z;
		19'b0010110100011010010: color_data = Z;
		19'b0010110100011010011: color_data = Z;
		19'b0010110100011010100: color_data = Z;
		19'b0010110100011010101: color_data = Z;
		19'b0010110100011010110: color_data = Z;
		19'b0010110100011010111: color_data = Z;
		19'b0010110100011011000: color_data = Z;
		19'b0010110100011011001: color_data = Z;
		19'b0010110100011011010: color_data = Z;
		19'b0010110100011011011: color_data = Z;
		19'b0010110100011011100: color_data = Z;
		19'b0010110100011011101: color_data = Z;
		19'b0010110100011011110: color_data = Z;
		19'b0010110100011011111: color_data = Z;
		19'b0010110100011100000: color_data = Z;
		19'b0010110100011100001: color_data = Z;
		19'b0010110100011100010: color_data = Z;
		19'b0010110100011100011: color_data = Z;
		19'b0010110100011100100: color_data = Z;
		19'b0010110100011100101: color_data = Z;
		19'b0010110100011100110: color_data = Z;
		19'b0010110100011100111: color_data = Z;
		19'b0010110100011101000: color_data = Z;
		19'b0010110100011101001: color_data = Z;
		19'b0010110100011101010: color_data = Z;
		19'b0010110100011101011: color_data = Z;
		19'b0010110100011101100: color_data = Z;
		19'b0010110100011101101: color_data = Z;
		19'b0010110100011101110: color_data = Z;
		19'b0010110100011101111: color_data = Z;
		19'b0010110100011110000: color_data = Z;
		19'b0010110100011110001: color_data = Z;
		19'b0010110100011110010: color_data = Z;
		19'b0010110100011110011: color_data = Z;
		19'b0010110100011110100: color_data = Z;
		19'b0010110100011110101: color_data = Z;
		19'b0010110100011110110: color_data = Z;
		19'b0010110100011110111: color_data = Z;
		19'b0010110100011111000: color_data = Z;
		19'b0010110100011111001: color_data = Z;
		19'b0010110100011111010: color_data = Z;
		19'b0010110100011111011: color_data = Z;
		19'b0010110100011111100: color_data = Z;
		19'b0010110100011111101: color_data = Z;
		19'b0010110100011111110: color_data = Z;
		19'b0010110100011111111: color_data = Z;
		19'b0010110100100000000: color_data = Z;
		19'b0010110100100000001: color_data = Z;
		19'b0010110100100000010: color_data = Z;
		19'b0010110100100000011: color_data = Z;
		19'b0010110100100000100: color_data = Z;
		19'b0010110100100000101: color_data = Z;
		19'b0010110100100000110: color_data = Z;
		19'b0010110100100000111: color_data = Z;
		19'b0010110100100001000: color_data = Z;
		19'b0010110100100001001: color_data = Z;
		19'b0010110100100001010: color_data = Z;
		19'b0010110100100001011: color_data = Z;
		19'b0010110100100001100: color_data = Z;
		19'b0010110100100001101: color_data = Z;
		19'b0010110100100001110: color_data = Z;
		19'b0010110100100001111: color_data = Z;
		19'b0010110100100010000: color_data = Z;
		19'b0010110100100010001: color_data = Z;
		19'b0010110100100010010: color_data = Z;
		19'b0010110100100010011: color_data = Z;
		19'b0010110100100010100: color_data = Z;
		19'b0010110100100010101: color_data = Z;
		19'b0010110100100010110: color_data = Z;
		19'b0010110100100010111: color_data = Z;
		19'b0010110100100011000: color_data = Z;
		19'b0010110100100011001: color_data = Z;
		19'b0010110100100011010: color_data = Z;
		19'b0010110100100011011: color_data = Z;
		19'b0010110100100011100: color_data = Z;
		19'b0010110100100011101: color_data = Z;
		19'b0010110100100011110: color_data = Z;
		19'b0010110100100011111: color_data = Z;
		19'b0010110100100100000: color_data = Z;
		19'b0010110100100100001: color_data = Z;
		19'b0010110100100100010: color_data = Z;
		19'b0010110100100100011: color_data = Z;
		19'b0010110100100100100: color_data = Z;
		19'b0010110100100100101: color_data = Z;
		19'b0010110100100100110: color_data = Z;
		19'b0010110100100100111: color_data = Z;
		19'b0010110100100101000: color_data = Z;
		19'b0010110100100101001: color_data = Z;
		19'b0010110100100101010: color_data = Z;
		19'b0010110100100101011: color_data = Z;
		19'b0010110100100101100: color_data = Z;
		19'b0010110100100101101: color_data = Z;
		19'b0010110100100101110: color_data = Z;
		19'b0010110100100101111: color_data = Z;
		19'b0010110100100110000: color_data = Z;
		19'b0010110100100110001: color_data = Z;
		19'b0010110100100110010: color_data = Z;
		19'b0010110100100110011: color_data = Z;
		19'b0010110100100110100: color_data = Z;
		19'b0010110100100110101: color_data = Z;
		19'b0010110100100110110: color_data = Z;
		19'b0010110100100110111: color_data = Z;
		19'b0010110100100111000: color_data = Z;
		19'b0010110100100111001: color_data = Z;
		19'b0010110100100111010: color_data = Z;
		19'b0010110100100111011: color_data = Z;
		19'b0010110100100111100: color_data = Z;
		19'b0010110100100111101: color_data = Z;
		19'b0010110100100111110: color_data = Z;
		19'b0010110100100111111: color_data = Z;
		19'b0010110100101000000: color_data = Z;
		19'b0010110100101000001: color_data = Z;
		19'b0010110100101000010: color_data = Z;
		19'b0010110100101000011: color_data = Z;
		19'b0010110100101000100: color_data = Z;
		19'b0010110100101000101: color_data = Z;
		19'b0010110100101000110: color_data = Z;
		19'b0010110100101000111: color_data = Z;
		19'b0010110100101001000: color_data = Z;
		19'b0010110100101001001: color_data = Z;
		19'b0010110100101001010: color_data = Z;
		19'b0010110100101001011: color_data = Z;
		19'b0010110100101001100: color_data = Z;
		19'b0010110100101001101: color_data = Z;
		19'b0010110100101001110: color_data = Z;
		19'b0010110100101001111: color_data = Z;
		19'b0010110100101010000: color_data = Z;
		19'b0010110100101010001: color_data = Z;
		19'b0010110100101010010: color_data = Z;
		19'b0010110100101010011: color_data = Z;
		19'b0010110100101010100: color_data = Z;
		19'b0010110100101010101: color_data = Z;
		19'b0010110100101010110: color_data = Z;
		19'b0010110100101010111: color_data = Z;
		19'b0010110100101011000: color_data = Z;
		19'b0010110100101011001: color_data = Z;
		19'b0010110100101011010: color_data = Z;
		19'b0010110100101011011: color_data = Z;
		19'b0010110100101011100: color_data = Z;
		19'b0010110100101011101: color_data = Z;
		19'b0010110100101011110: color_data = Z;
		19'b0010110100101011111: color_data = Z;
		19'b0010110100101100000: color_data = Z;
		19'b0010110100101100001: color_data = Z;
		19'b0010110100101100010: color_data = Z;
		19'b0010110100101100011: color_data = Z;
		19'b0010110100101100100: color_data = Z;
		19'b0010110100101100101: color_data = Z;
		19'b0010110100101100110: color_data = Z;
		19'b0010110100101100111: color_data = Z;
		19'b0010110100101101000: color_data = Z;
		19'b0010110100101101001: color_data = Z;
		19'b0010110100101101010: color_data = Z;
		19'b0010110100101101011: color_data = Z;
		19'b0010110100101101100: color_data = Z;
		19'b0010110100101101101: color_data = Z;
		19'b0010110100101101110: color_data = Z;
		19'b0010110100101101111: color_data = Z;
		19'b0010110100101110000: color_data = Z;
		19'b0010110100101110001: color_data = Z;
		19'b0010110100101110010: color_data = Z;
		19'b0010110100101110011: color_data = Z;
		19'b0010110100101110100: color_data = Z;
		19'b0010110100101110101: color_data = Z;
		19'b0010110100101110110: color_data = Z;
		19'b0010110100101110111: color_data = Z;
		19'b0010110100101111000: color_data = Z;
		19'b0010110100101111001: color_data = Z;
		19'b0010110100101111010: color_data = Z;
		19'b0010110100101111011: color_data = Z;
		19'b0010110100101111100: color_data = Z;
		19'b0010110100101111101: color_data = Z;
		19'b0010110100101111110: color_data = Z;
		19'b0010110100101111111: color_data = Z;
		19'b0010110100110000000: color_data = Z;
		19'b0010110100110000001: color_data = Z;
		19'b0010110100110000010: color_data = Z;
		19'b0010110100110000011: color_data = Z;
		19'b0010110100110000100: color_data = Z;
		19'b0010110100110000101: color_data = Z;
		19'b0010110100110000110: color_data = Z;
		19'b0010110100110000111: color_data = Z;
		19'b0010110100110001000: color_data = Z;
		19'b0010110100110001001: color_data = Z;
		19'b0010110100110001010: color_data = Z;
		19'b0010110100110001011: color_data = Z;
		19'b0010110100110001100: color_data = Z;
		19'b0010110100110001101: color_data = Z;
		19'b0010110100110001110: color_data = Z;
		19'b0010110100110001111: color_data = Z;
		19'b0010110100110010000: color_data = Z;
		19'b0010110100110010001: color_data = Z;
		19'b0010110100110010010: color_data = Z;
		19'b0010110100110010011: color_data = Z;
		19'b0010110100110010100: color_data = Z;
		19'b0010110100110010101: color_data = Z;
		19'b0010110100110010110: color_data = Z;
		19'b0010110100110010111: color_data = Z;
		19'b0010110100110011000: color_data = Z;
		19'b0010110100110011001: color_data = Z;
		19'b0010110100110011010: color_data = Z;
		19'b0010110100110011011: color_data = Z;
		19'b0010110100110011100: color_data = Z;
		19'b0010110100110011101: color_data = Z;
		19'b0010110100110011110: color_data = Z;
		19'b0010110100110011111: color_data = Z;
		19'b0010110100110100000: color_data = Z;
		19'b0010110100110100001: color_data = Z;
		19'b0010110100110100010: color_data = Z;
		19'b0010110100110100011: color_data = Z;
		19'b0010110100110100100: color_data = Z;
		19'b0010110100110100101: color_data = Z;
		19'b0010110100110100110: color_data = Z;
		19'b0010110100110100111: color_data = Z;
		19'b0010110100110101000: color_data = Z;
		19'b0010110100110101001: color_data = Z;
		19'b0010110100110101010: color_data = Z;
		19'b0010110100110101011: color_data = Z;
		19'b0010110100110101100: color_data = Z;
		19'b0010110100110101101: color_data = Z;
		19'b0010110100110101110: color_data = Z;
		19'b0010110100110101111: color_data = Z;
		19'b0010110100110110000: color_data = Z;
		19'b0010110100110110001: color_data = Z;
		19'b0010110100110110010: color_data = Z;
		19'b0010110100110111011: color_data = Z;
		19'b0010110100111000010: color_data = Z;
		19'b0010110100111000011: color_data = Z;
		19'b0010110100111000100: color_data = Z;
		19'b0010110100111000101: color_data = Z;
		19'b0010110100111000110: color_data = Z;
		19'b0010110100111000111: color_data = Z;
		19'b0010110100111001000: color_data = Z;
		19'b0010110100111001001: color_data = Z;
		19'b0010110100111001010: color_data = Z;
		19'b0010110100111001011: color_data = Z;
		19'b0010110100111001100: color_data = Z;
		19'b0010110100111001101: color_data = Z;
		19'b0010110100111001110: color_data = Z;
		19'b0010110110011000000: color_data = Z;
		19'b0010110110011000001: color_data = Z;
		19'b0010110110011000010: color_data = Z;
		19'b0010110110011000011: color_data = Z;
		19'b0010110110011000100: color_data = Z;
		19'b0010110110011000101: color_data = Z;
		19'b0010110110011000110: color_data = Z;
		19'b0010110110011000111: color_data = Z;
		19'b0010110110011001000: color_data = Z;
		19'b0010110110011001001: color_data = Z;
		19'b0010110110011001010: color_data = Z;
		19'b0010110110011001011: color_data = Z;
		19'b0010110110011001100: color_data = Z;
		19'b0010110110011001101: color_data = Z;
		19'b0010110110011001110: color_data = Z;
		19'b0010110110011001111: color_data = Z;
		19'b0010110110011010000: color_data = Z;
		19'b0010110110011010001: color_data = Z;
		19'b0010110110011010010: color_data = Z;
		19'b0010110110011010011: color_data = Z;
		19'b0010110110011010100: color_data = Z;
		19'b0010110110011010101: color_data = Z;
		19'b0010110110011010110: color_data = Z;
		19'b0010110110011010111: color_data = Z;
		19'b0010110110011011000: color_data = Z;
		19'b0010110110011011001: color_data = Z;
		19'b0010110110011011010: color_data = Z;
		19'b0010110110011011011: color_data = Z;
		19'b0010110110011011100: color_data = Z;
		19'b0010110110011011101: color_data = Z;
		19'b0010110110011011110: color_data = Z;
		19'b0010110110011011111: color_data = Z;
		19'b0010110110011100000: color_data = Z;
		19'b0010110110011100001: color_data = Z;
		19'b0010110110011100010: color_data = Z;
		19'b0010110110011100011: color_data = Z;
		19'b0010110110011100100: color_data = Z;
		19'b0010110110011100101: color_data = Z;
		19'b0010110110011100110: color_data = Z;
		19'b0010110110011100111: color_data = Z;
		19'b0010110110011101000: color_data = Z;
		19'b0010110110011101001: color_data = Z;
		19'b0010110110011101010: color_data = Z;
		19'b0010110110011101011: color_data = Z;
		19'b0010110110011101100: color_data = Z;
		19'b0010110110011101101: color_data = Z;
		19'b0010110110011101110: color_data = Z;
		19'b0010110110011101111: color_data = Z;
		19'b0010110110011110000: color_data = Z;
		19'b0010110110011110001: color_data = Z;
		19'b0010110110011110010: color_data = Z;
		19'b0010110110011110011: color_data = Z;
		19'b0010110110011110100: color_data = Z;
		19'b0010110110011110101: color_data = Z;
		19'b0010110110011110110: color_data = Z;
		19'b0010110110011110111: color_data = Z;
		19'b0010110110011111000: color_data = Z;
		19'b0010110110011111001: color_data = Z;
		19'b0010110110011111010: color_data = Z;
		19'b0010110110011111011: color_data = Z;
		19'b0010110110011111100: color_data = Z;
		19'b0010110110011111101: color_data = Z;
		19'b0010110110011111110: color_data = Z;
		19'b0010110110011111111: color_data = Z;
		19'b0010110110100000000: color_data = Z;
		19'b0010110110100000001: color_data = Z;
		19'b0010110110100000010: color_data = Z;
		19'b0010110110100000011: color_data = Z;
		19'b0010110110100000100: color_data = Z;
		19'b0010110110100000101: color_data = Z;
		19'b0010110110100000110: color_data = Z;
		19'b0010110110100000111: color_data = Z;
		19'b0010110110100001000: color_data = Z;
		19'b0010110110100001001: color_data = Z;
		19'b0010110110100001010: color_data = Z;
		19'b0010110110100001011: color_data = Z;
		19'b0010110110100001100: color_data = Z;
		19'b0010110110100001101: color_data = Z;
		19'b0010110110100001110: color_data = Z;
		19'b0010110110100001111: color_data = Z;
		19'b0010110110100010000: color_data = Z;
		19'b0010110110100010001: color_data = Z;
		19'b0010110110100010010: color_data = Z;
		19'b0010110110100010011: color_data = Z;
		19'b0010110110100010100: color_data = Z;
		19'b0010110110100010101: color_data = Z;
		19'b0010110110100010110: color_data = Z;
		19'b0010110110100010111: color_data = Z;
		19'b0010110110100011000: color_data = Z;
		19'b0010110110100011001: color_data = Z;
		19'b0010110110100011010: color_data = Z;
		19'b0010110110100011011: color_data = Z;
		19'b0010110110100011100: color_data = Z;
		19'b0010110110100011101: color_data = Z;
		19'b0010110110100011110: color_data = Z;
		19'b0010110110100011111: color_data = Z;
		19'b0010110110100100000: color_data = Z;
		19'b0010110110100100001: color_data = Z;
		19'b0010110110100100010: color_data = Z;
		19'b0010110110100100011: color_data = Z;
		19'b0010110110100100100: color_data = Z;
		19'b0010110110100100101: color_data = Z;
		19'b0010110110100100110: color_data = Z;
		19'b0010110110100100111: color_data = Z;
		19'b0010110110100101000: color_data = Z;
		19'b0010110110100101001: color_data = Z;
		19'b0010110110100101010: color_data = Z;
		19'b0010110110100101011: color_data = Z;
		19'b0010110110100101100: color_data = Z;
		19'b0010110110100101101: color_data = Z;
		19'b0010110110100101110: color_data = Z;
		19'b0010110110100101111: color_data = Z;
		19'b0010110110100110000: color_data = Z;
		19'b0010110110100110001: color_data = Z;
		19'b0010110110100110010: color_data = Z;
		19'b0010110110100110011: color_data = Z;
		19'b0010110110100110100: color_data = Z;
		19'b0010110110100110101: color_data = Z;
		19'b0010110110100110110: color_data = Z;
		19'b0010110110100110111: color_data = Z;
		19'b0010110110100111000: color_data = Z;
		19'b0010110110100111001: color_data = Z;
		19'b0010110110100111010: color_data = Z;
		19'b0010110110100111011: color_data = Z;
		19'b0010110110100111100: color_data = Z;
		19'b0010110110100111101: color_data = Z;
		19'b0010110110100111110: color_data = Z;
		19'b0010110110100111111: color_data = Z;
		19'b0010110110101000000: color_data = Z;
		19'b0010110110101000001: color_data = Z;
		19'b0010110110101000010: color_data = Z;
		19'b0010110110101000011: color_data = Z;
		19'b0010110110101000100: color_data = Z;
		19'b0010110110101000101: color_data = Z;
		19'b0010110110101000110: color_data = Z;
		19'b0010110110101000111: color_data = Z;
		19'b0010110110101001000: color_data = Z;
		19'b0010110110101001001: color_data = Z;
		19'b0010110110101001010: color_data = Z;
		19'b0010110110101001011: color_data = Z;
		19'b0010110110101001100: color_data = Z;
		19'b0010110110101001101: color_data = Z;
		19'b0010110110101001110: color_data = Z;
		19'b0010110110101001111: color_data = Z;
		19'b0010110110101010000: color_data = Z;
		19'b0010110110101010001: color_data = Z;
		19'b0010110110101010010: color_data = Z;
		19'b0010110110101010011: color_data = Z;
		19'b0010110110101010100: color_data = Z;
		19'b0010110110101010101: color_data = Z;
		19'b0010110110101010110: color_data = Z;
		19'b0010110110101010111: color_data = Z;
		19'b0010110110101011000: color_data = Z;
		19'b0010110110101011001: color_data = Z;
		19'b0010110110101011010: color_data = Z;
		19'b0010110110101011011: color_data = Z;
		19'b0010110110101011100: color_data = Z;
		19'b0010110110101011101: color_data = Z;
		19'b0010110110101011110: color_data = Z;
		19'b0010110110101011111: color_data = Z;
		19'b0010110110101100000: color_data = Z;
		19'b0010110110101100001: color_data = Z;
		19'b0010110110101100010: color_data = Z;
		19'b0010110110101100011: color_data = Z;
		19'b0010110110101100100: color_data = Z;
		19'b0010110110101100101: color_data = Z;
		19'b0010110110101100110: color_data = Z;
		19'b0010110110101100111: color_data = Z;
		19'b0010110110101101000: color_data = Z;
		19'b0010110110101101001: color_data = Z;
		19'b0010110110101101010: color_data = Z;
		19'b0010110110101101011: color_data = Z;
		19'b0010110110101101100: color_data = Z;
		19'b0010110110101101101: color_data = Z;
		19'b0010110110101101110: color_data = Z;
		19'b0010110110101101111: color_data = Z;
		19'b0010110110101110000: color_data = Z;
		19'b0010110110101110001: color_data = Z;
		19'b0010110110101110010: color_data = Z;
		19'b0010110110101110011: color_data = Z;
		19'b0010110110101110100: color_data = Z;
		19'b0010110110101110101: color_data = Z;
		19'b0010110110101110110: color_data = Z;
		19'b0010110110101110111: color_data = Z;
		19'b0010110110101111000: color_data = Z;
		19'b0010110110101111001: color_data = Z;
		19'b0010110110101111010: color_data = Z;
		19'b0010110110101111011: color_data = Z;
		19'b0010110110101111100: color_data = Z;
		19'b0010110110101111101: color_data = Z;
		19'b0010110110101111110: color_data = Z;
		19'b0010110110101111111: color_data = Z;
		19'b0010110110110000000: color_data = Z;
		19'b0010110110110000001: color_data = Z;
		19'b0010110110110000010: color_data = Z;
		19'b0010110110110000011: color_data = Z;
		19'b0010110110110000100: color_data = Z;
		19'b0010110110110000101: color_data = Z;
		19'b0010110110110000110: color_data = Z;
		19'b0010110110110000111: color_data = Z;
		19'b0010110110110001000: color_data = Z;
		19'b0010110110110001001: color_data = Z;
		19'b0010110110110001010: color_data = Z;
		19'b0010110110110001011: color_data = Z;
		19'b0010110110110001100: color_data = Z;
		19'b0010110110110001101: color_data = Z;
		19'b0010110110110001110: color_data = Z;
		19'b0010110110110001111: color_data = Z;
		19'b0010110110110010000: color_data = Z;
		19'b0010110110110010001: color_data = Z;
		19'b0010110110110010010: color_data = Z;
		19'b0010110110110010011: color_data = Z;
		19'b0010110110110010100: color_data = Z;
		19'b0010110110110010101: color_data = Z;
		19'b0010110110110010110: color_data = Z;
		19'b0010110110110010111: color_data = Z;
		19'b0010110110110011000: color_data = Z;
		19'b0010110110110011001: color_data = Z;
		19'b0010110110110011010: color_data = Z;
		19'b0010110110110011011: color_data = Z;
		19'b0010110110110011100: color_data = Z;
		19'b0010110110110011101: color_data = Z;
		19'b0010110110110011110: color_data = Z;
		19'b0010110110110011111: color_data = Z;
		19'b0010110110110100000: color_data = Z;
		19'b0010110110110100001: color_data = Z;
		19'b0010110110110100010: color_data = Z;
		19'b0010110110110100011: color_data = Z;
		19'b0010110110110100100: color_data = Z;
		19'b0010110110110100101: color_data = Z;
		19'b0010110110110100110: color_data = Z;
		19'b0010110110110100111: color_data = Z;
		19'b0010110110110101000: color_data = Z;
		19'b0010110110110101001: color_data = Z;
		19'b0010110110110101010: color_data = Z;
		19'b0010110110110101011: color_data = Z;
		19'b0010110110110101100: color_data = Z;
		19'b0010110110110101101: color_data = Z;
		19'b0010110110110101110: color_data = Z;
		19'b0010110110110101111: color_data = Z;
		19'b0010110110110110000: color_data = Z;
		19'b0010110110110110001: color_data = Z;
		19'b0010110110110110010: color_data = Z;
		19'b0010110110110110011: color_data = Z;
		19'b0010110110110111011: color_data = Z;
		19'b0010110110111000011: color_data = Z;
		19'b0010110110111000100: color_data = Z;
		19'b0010110110111000101: color_data = Z;
		19'b0010110110111000110: color_data = Z;
		19'b0010110110111000111: color_data = Z;
		19'b0010110110111001000: color_data = Z;
		19'b0010110110111001001: color_data = Z;
		19'b0010110110111001010: color_data = Z;
		19'b0010110110111001011: color_data = Z;
		19'b0010110110111001100: color_data = Z;
		19'b0010110110111001101: color_data = Z;
		19'b0010110110111001110: color_data = Z;
		19'b0010111000010111111: color_data = Z;
		19'b0010111000011000000: color_data = Z;
		19'b0010111000011000001: color_data = Z;
		19'b0010111000011000010: color_data = Z;
		19'b0010111000011000011: color_data = Z;
		19'b0010111000011000100: color_data = Z;
		19'b0010111000011000101: color_data = Z;
		19'b0010111000011000110: color_data = Z;
		19'b0010111000011000111: color_data = Z;
		19'b0010111000011001000: color_data = Z;
		19'b0010111000011001001: color_data = Z;
		19'b0010111000011001010: color_data = Z;
		19'b0010111000011001011: color_data = Z;
		19'b0010111000011001100: color_data = Z;
		19'b0010111000011001101: color_data = Z;
		19'b0010111000011001110: color_data = Z;
		19'b0010111000011001111: color_data = Z;
		19'b0010111000011010000: color_data = Z;
		19'b0010111000011010001: color_data = Z;
		19'b0010111000011010010: color_data = Z;
		19'b0010111000011010011: color_data = Z;
		19'b0010111000011010100: color_data = Z;
		19'b0010111000011010101: color_data = Z;
		19'b0010111000011010110: color_data = Z;
		19'b0010111000011010111: color_data = Z;
		19'b0010111000011011000: color_data = Z;
		19'b0010111000011011001: color_data = Z;
		19'b0010111000011011010: color_data = Z;
		19'b0010111000011011011: color_data = Z;
		19'b0010111000011011100: color_data = Z;
		19'b0010111000011011101: color_data = Z;
		19'b0010111000011011110: color_data = Z;
		19'b0010111000011011111: color_data = Z;
		19'b0010111000011100000: color_data = Z;
		19'b0010111000011100001: color_data = Z;
		19'b0010111000011100010: color_data = Z;
		19'b0010111000011100011: color_data = Z;
		19'b0010111000011100100: color_data = Z;
		19'b0010111000011100101: color_data = Z;
		19'b0010111000011100110: color_data = Z;
		19'b0010111000011100111: color_data = Z;
		19'b0010111000011101000: color_data = Z;
		19'b0010111000011101001: color_data = Z;
		19'b0010111000011101010: color_data = Z;
		19'b0010111000011101011: color_data = Z;
		19'b0010111000011101100: color_data = Z;
		19'b0010111000011101101: color_data = Z;
		19'b0010111000011101110: color_data = Z;
		19'b0010111000011101111: color_data = Z;
		19'b0010111000011110000: color_data = Z;
		19'b0010111000011110001: color_data = Z;
		19'b0010111000011110010: color_data = Z;
		19'b0010111000011110011: color_data = Z;
		19'b0010111000011110100: color_data = Z;
		19'b0010111000011110101: color_data = Z;
		19'b0010111000011110110: color_data = Z;
		19'b0010111000011110111: color_data = Z;
		19'b0010111000011111000: color_data = Z;
		19'b0010111000011111001: color_data = Z;
		19'b0010111000011111010: color_data = Z;
		19'b0010111000011111011: color_data = Z;
		19'b0010111000011111100: color_data = Z;
		19'b0010111000011111101: color_data = Z;
		19'b0010111000011111110: color_data = Z;
		19'b0010111000011111111: color_data = Z;
		19'b0010111000100000000: color_data = Z;
		19'b0010111000100000001: color_data = Z;
		19'b0010111000100000010: color_data = Z;
		19'b0010111000100000011: color_data = Z;
		19'b0010111000100000100: color_data = Z;
		19'b0010111000100000101: color_data = Z;
		19'b0010111000100000110: color_data = Z;
		19'b0010111000100000111: color_data = Z;
		19'b0010111000100001000: color_data = Z;
		19'b0010111000100001001: color_data = Z;
		19'b0010111000100001010: color_data = Z;
		19'b0010111000100001011: color_data = Z;
		19'b0010111000100001100: color_data = Z;
		19'b0010111000100001101: color_data = Z;
		19'b0010111000100001110: color_data = Z;
		19'b0010111000100001111: color_data = Z;
		19'b0010111000100010000: color_data = Z;
		19'b0010111000100010001: color_data = Z;
		19'b0010111000100010010: color_data = Z;
		19'b0010111000100010011: color_data = Z;
		19'b0010111000100010100: color_data = Z;
		19'b0010111000100010101: color_data = Z;
		19'b0010111000100010110: color_data = Z;
		19'b0010111000100010111: color_data = Z;
		19'b0010111000100011000: color_data = Z;
		19'b0010111000100011001: color_data = Z;
		19'b0010111000100011010: color_data = Z;
		19'b0010111000100011011: color_data = Z;
		19'b0010111000100011100: color_data = Z;
		19'b0010111000100011101: color_data = Z;
		19'b0010111000100011110: color_data = Z;
		19'b0010111000100011111: color_data = Z;
		19'b0010111000100100000: color_data = Z;
		19'b0010111000100100001: color_data = Z;
		19'b0010111000100100010: color_data = Z;
		19'b0010111000100100011: color_data = Z;
		19'b0010111000100100100: color_data = Z;
		19'b0010111000100100101: color_data = Z;
		19'b0010111000100100110: color_data = Z;
		19'b0010111000100100111: color_data = Z;
		19'b0010111000100101000: color_data = Z;
		19'b0010111000100101001: color_data = Z;
		19'b0010111000100101010: color_data = Z;
		19'b0010111000100101011: color_data = Z;
		19'b0010111000100101100: color_data = Z;
		19'b0010111000100101101: color_data = Z;
		19'b0010111000100101110: color_data = Z;
		19'b0010111000100101111: color_data = Z;
		19'b0010111000100110000: color_data = Z;
		19'b0010111000100110001: color_data = Z;
		19'b0010111000100110010: color_data = Z;
		19'b0010111000100110011: color_data = Z;
		19'b0010111000100110100: color_data = Z;
		19'b0010111000100110101: color_data = Z;
		19'b0010111000100110110: color_data = Z;
		19'b0010111000100110111: color_data = Z;
		19'b0010111000100111000: color_data = Z;
		19'b0010111000100111001: color_data = Z;
		19'b0010111000100111010: color_data = Z;
		19'b0010111000100111011: color_data = Z;
		19'b0010111000100111100: color_data = Z;
		19'b0010111000100111101: color_data = Z;
		19'b0010111000100111110: color_data = Z;
		19'b0010111000100111111: color_data = Z;
		19'b0010111000101000000: color_data = Z;
		19'b0010111000101000001: color_data = Z;
		19'b0010111000101000010: color_data = Z;
		19'b0010111000101000011: color_data = Z;
		19'b0010111000101000100: color_data = Z;
		19'b0010111000101000101: color_data = Z;
		19'b0010111000101000110: color_data = Z;
		19'b0010111000101000111: color_data = Z;
		19'b0010111000101001000: color_data = Z;
		19'b0010111000101001001: color_data = Z;
		19'b0010111000101001010: color_data = Z;
		19'b0010111000101001011: color_data = Z;
		19'b0010111000101001100: color_data = Z;
		19'b0010111000101001101: color_data = Z;
		19'b0010111000101001110: color_data = Z;
		19'b0010111000101001111: color_data = Z;
		19'b0010111000101010000: color_data = Z;
		19'b0010111000101010001: color_data = Z;
		19'b0010111000101010010: color_data = Z;
		19'b0010111000101010011: color_data = Z;
		19'b0010111000101010100: color_data = Z;
		19'b0010111000101010101: color_data = Z;
		19'b0010111000101010110: color_data = Z;
		19'b0010111000101010111: color_data = Z;
		19'b0010111000101011000: color_data = Z;
		19'b0010111000101011001: color_data = Z;
		19'b0010111000101011010: color_data = Z;
		19'b0010111000101011011: color_data = Z;
		19'b0010111000101011100: color_data = Z;
		19'b0010111000101011101: color_data = Z;
		19'b0010111000101011110: color_data = Z;
		19'b0010111000101011111: color_data = Z;
		19'b0010111000101100000: color_data = Z;
		19'b0010111000101100001: color_data = Z;
		19'b0010111000101100010: color_data = Z;
		19'b0010111000101100011: color_data = Z;
		19'b0010111000101100100: color_data = Z;
		19'b0010111000101100101: color_data = Z;
		19'b0010111000101100110: color_data = Z;
		19'b0010111000101100111: color_data = Z;
		19'b0010111000101101000: color_data = Z;
		19'b0010111000101101001: color_data = Z;
		19'b0010111000101101010: color_data = Z;
		19'b0010111000101101011: color_data = Z;
		19'b0010111000101101100: color_data = Z;
		19'b0010111000101101101: color_data = Z;
		19'b0010111000101101110: color_data = Z;
		19'b0010111000101101111: color_data = Z;
		19'b0010111000101110000: color_data = Z;
		19'b0010111000101110001: color_data = Z;
		19'b0010111000101110010: color_data = Z;
		19'b0010111000101110011: color_data = Z;
		19'b0010111000101110100: color_data = Z;
		19'b0010111000101110101: color_data = Z;
		19'b0010111000101110110: color_data = Z;
		19'b0010111000101110111: color_data = Z;
		19'b0010111000101111000: color_data = Z;
		19'b0010111000101111001: color_data = Z;
		19'b0010111000101111010: color_data = Z;
		19'b0010111000101111011: color_data = Z;
		19'b0010111000101111100: color_data = Z;
		19'b0010111000101111101: color_data = Z;
		19'b0010111000101111110: color_data = Z;
		19'b0010111000101111111: color_data = Z;
		19'b0010111000110000000: color_data = Z;
		19'b0010111000110000001: color_data = Z;
		19'b0010111000110000010: color_data = Z;
		19'b0010111000110000011: color_data = Z;
		19'b0010111000110000100: color_data = Z;
		19'b0010111000110000101: color_data = Z;
		19'b0010111000110000110: color_data = Z;
		19'b0010111000110000111: color_data = Z;
		19'b0010111000110001000: color_data = Z;
		19'b0010111000110001001: color_data = Z;
		19'b0010111000110001010: color_data = Z;
		19'b0010111000110001011: color_data = Z;
		19'b0010111000110001100: color_data = Z;
		19'b0010111000110001101: color_data = Z;
		19'b0010111000110001110: color_data = Z;
		19'b0010111000110001111: color_data = Z;
		19'b0010111000110010000: color_data = Z;
		19'b0010111000110010001: color_data = Z;
		19'b0010111000110010010: color_data = Z;
		19'b0010111000110010011: color_data = Z;
		19'b0010111000110010100: color_data = Z;
		19'b0010111000110010101: color_data = Z;
		19'b0010111000110010110: color_data = Z;
		19'b0010111000110010111: color_data = Z;
		19'b0010111000110011000: color_data = Z;
		19'b0010111000110011001: color_data = Z;
		19'b0010111000110011010: color_data = Z;
		19'b0010111000110011011: color_data = Z;
		19'b0010111000110011100: color_data = Z;
		19'b0010111000110011101: color_data = Z;
		19'b0010111000110011110: color_data = Z;
		19'b0010111000110011111: color_data = Z;
		19'b0010111000110100000: color_data = Z;
		19'b0010111000110100001: color_data = Z;
		19'b0010111000110100010: color_data = Z;
		19'b0010111000110100011: color_data = Z;
		19'b0010111000110100100: color_data = Z;
		19'b0010111000110100101: color_data = Z;
		19'b0010111000110100110: color_data = Z;
		19'b0010111000110100111: color_data = Z;
		19'b0010111000110101000: color_data = Z;
		19'b0010111000110101001: color_data = Z;
		19'b0010111000110101010: color_data = Z;
		19'b0010111000110101011: color_data = Z;
		19'b0010111000110101100: color_data = Z;
		19'b0010111000110101101: color_data = Z;
		19'b0010111000110101110: color_data = Z;
		19'b0010111000110101111: color_data = Z;
		19'b0010111000110110000: color_data = Z;
		19'b0010111000110110001: color_data = Z;
		19'b0010111000110110010: color_data = Z;
		19'b0010111000110110011: color_data = Z;
		19'b0010111000111000011: color_data = Z;
		19'b0010111000111000100: color_data = Z;
		19'b0010111000111000101: color_data = Z;
		19'b0010111000111000110: color_data = Z;
		19'b0010111000111000111: color_data = Z;
		19'b0010111000111001000: color_data = Z;
		19'b0010111000111001001: color_data = Z;
		19'b0010111000111001010: color_data = Z;
		19'b0010111000111001011: color_data = Z;
		19'b0010111000111001100: color_data = Z;
		19'b0010111000111001101: color_data = Z;
		19'b0010111000111001110: color_data = Z;
		19'b0010111010010111110: color_data = Z;
		19'b0010111010010111111: color_data = Z;
		19'b0010111010011000000: color_data = Z;
		19'b0010111010011000001: color_data = Z;
		19'b0010111010011000010: color_data = Z;
		19'b0010111010011000011: color_data = Z;
		19'b0010111010011000100: color_data = Z;
		19'b0010111010011000101: color_data = Z;
		19'b0010111010011000110: color_data = Z;
		19'b0010111010011000111: color_data = Z;
		19'b0010111010011001000: color_data = Z;
		19'b0010111010011001001: color_data = Z;
		19'b0010111010011001010: color_data = Z;
		19'b0010111010011001011: color_data = Z;
		19'b0010111010011001100: color_data = Z;
		19'b0010111010011001101: color_data = Z;
		19'b0010111010011001110: color_data = Z;
		19'b0010111010011001111: color_data = Z;
		19'b0010111010011010000: color_data = Z;
		19'b0010111010011010001: color_data = Z;
		19'b0010111010011010010: color_data = Z;
		19'b0010111010011010011: color_data = Z;
		19'b0010111010011010100: color_data = Z;
		19'b0010111010011010101: color_data = Z;
		19'b0010111010011010110: color_data = Z;
		19'b0010111010011010111: color_data = Z;
		19'b0010111010011011000: color_data = Z;
		19'b0010111010011011001: color_data = Z;
		19'b0010111010011011010: color_data = Z;
		19'b0010111010011011011: color_data = Z;
		19'b0010111010011011100: color_data = Z;
		19'b0010111010011011101: color_data = Z;
		19'b0010111010011011110: color_data = Z;
		19'b0010111010011011111: color_data = Z;
		19'b0010111010011100000: color_data = Z;
		19'b0010111010011100001: color_data = Z;
		19'b0010111010011100010: color_data = Z;
		19'b0010111010011100011: color_data = Z;
		19'b0010111010011100100: color_data = Z;
		19'b0010111010011100101: color_data = Z;
		19'b0010111010011100110: color_data = Z;
		19'b0010111010011100111: color_data = Z;
		19'b0010111010011101000: color_data = Z;
		19'b0010111010011101001: color_data = Z;
		19'b0010111010011101010: color_data = Z;
		19'b0010111010011101011: color_data = Z;
		19'b0010111010011101100: color_data = Z;
		19'b0010111010011101101: color_data = Z;
		19'b0010111010011101110: color_data = Z;
		19'b0010111010011101111: color_data = Z;
		19'b0010111010011110000: color_data = Z;
		19'b0010111010011110001: color_data = Z;
		19'b0010111010011110010: color_data = Z;
		19'b0010111010011110011: color_data = Z;
		19'b0010111010011110100: color_data = Z;
		19'b0010111010011110101: color_data = Z;
		19'b0010111010011110110: color_data = Z;
		19'b0010111010011110111: color_data = Z;
		19'b0010111010011111000: color_data = Z;
		19'b0010111010011111001: color_data = Z;
		19'b0010111010011111010: color_data = Z;
		19'b0010111010011111011: color_data = Z;
		19'b0010111010011111100: color_data = Z;
		19'b0010111010011111101: color_data = Z;
		19'b0010111010011111110: color_data = Z;
		19'b0010111010011111111: color_data = Z;
		19'b0010111010100000000: color_data = Z;
		19'b0010111010100000001: color_data = Z;
		19'b0010111010100000010: color_data = Z;
		19'b0010111010100000011: color_data = Z;
		19'b0010111010100000100: color_data = Z;
		19'b0010111010100000101: color_data = Z;
		19'b0010111010100000110: color_data = Z;
		19'b0010111010100000111: color_data = Z;
		19'b0010111010100001000: color_data = Z;
		19'b0010111010100001001: color_data = Z;
		19'b0010111010100001010: color_data = Z;
		19'b0010111010100001011: color_data = Z;
		19'b0010111010100001100: color_data = Z;
		19'b0010111010100001101: color_data = Z;
		19'b0010111010100001110: color_data = Z;
		19'b0010111010100001111: color_data = Z;
		19'b0010111010100010000: color_data = Z;
		19'b0010111010100010001: color_data = Z;
		19'b0010111010100010010: color_data = Z;
		19'b0010111010100010011: color_data = Z;
		19'b0010111010100010100: color_data = Z;
		19'b0010111010100010101: color_data = Z;
		19'b0010111010100010110: color_data = Z;
		19'b0010111010100010111: color_data = Z;
		19'b0010111010100011000: color_data = Z;
		19'b0010111010100011001: color_data = Z;
		19'b0010111010100011010: color_data = Z;
		19'b0010111010100011011: color_data = Z;
		19'b0010111010100011100: color_data = Z;
		19'b0010111010100011101: color_data = Z;
		19'b0010111010100011110: color_data = Z;
		19'b0010111010100011111: color_data = Z;
		19'b0010111010100100000: color_data = Z;
		19'b0010111010100100001: color_data = Z;
		19'b0010111010100100010: color_data = Z;
		19'b0010111010100100011: color_data = Z;
		19'b0010111010100100100: color_data = Z;
		19'b0010111010100100101: color_data = Z;
		19'b0010111010100100110: color_data = Z;
		19'b0010111010100100111: color_data = Z;
		19'b0010111010100101000: color_data = Z;
		19'b0010111010100101001: color_data = Z;
		19'b0010111010100101010: color_data = Z;
		19'b0010111010100101011: color_data = Z;
		19'b0010111010100101100: color_data = Z;
		19'b0010111010100101101: color_data = Z;
		19'b0010111010100101110: color_data = Z;
		19'b0010111010100101111: color_data = Z;
		19'b0010111010100110000: color_data = Z;
		19'b0010111010100110001: color_data = Z;
		19'b0010111010100110010: color_data = Z;
		19'b0010111010100110011: color_data = Z;
		19'b0010111010100110100: color_data = Z;
		19'b0010111010100110101: color_data = Z;
		19'b0010111010100110110: color_data = Z;
		19'b0010111010100110111: color_data = Z;
		19'b0010111010100111000: color_data = Z;
		19'b0010111010100111001: color_data = Z;
		19'b0010111010100111010: color_data = Z;
		19'b0010111010100111011: color_data = Z;
		19'b0010111010100111100: color_data = Z;
		19'b0010111010100111101: color_data = Z;
		19'b0010111010100111110: color_data = Z;
		19'b0010111010100111111: color_data = Z;
		19'b0010111010101000000: color_data = Z;
		19'b0010111010101000001: color_data = Z;
		19'b0010111010101000010: color_data = Z;
		19'b0010111010101000011: color_data = Z;
		19'b0010111010101000100: color_data = Z;
		19'b0010111010101000101: color_data = Z;
		19'b0010111010101000110: color_data = Z;
		19'b0010111010101000111: color_data = Z;
		19'b0010111010101001000: color_data = Z;
		19'b0010111010101001001: color_data = Z;
		19'b0010111010101001010: color_data = Z;
		19'b0010111010101001011: color_data = Z;
		19'b0010111010101001100: color_data = Z;
		19'b0010111010101001101: color_data = Z;
		19'b0010111010101001110: color_data = Z;
		19'b0010111010101001111: color_data = Z;
		19'b0010111010101010000: color_data = Z;
		19'b0010111010101010001: color_data = Z;
		19'b0010111010101010010: color_data = Z;
		19'b0010111010101010011: color_data = Z;
		19'b0010111010101010100: color_data = Z;
		19'b0010111010101010101: color_data = Z;
		19'b0010111010101010110: color_data = Z;
		19'b0010111010101010111: color_data = Z;
		19'b0010111010101011000: color_data = Z;
		19'b0010111010101011001: color_data = Z;
		19'b0010111010101011010: color_data = Z;
		19'b0010111010101011011: color_data = Z;
		19'b0010111010101011100: color_data = Z;
		19'b0010111010101011101: color_data = Z;
		19'b0010111010101011110: color_data = Z;
		19'b0010111010101011111: color_data = Z;
		19'b0010111010101100000: color_data = Z;
		19'b0010111010101100001: color_data = Z;
		19'b0010111010101100010: color_data = Z;
		19'b0010111010101100011: color_data = Z;
		19'b0010111010101100100: color_data = Z;
		19'b0010111010101100101: color_data = Z;
		19'b0010111010101100110: color_data = Z;
		19'b0010111010101100111: color_data = Z;
		19'b0010111010101101000: color_data = Z;
		19'b0010111010101101001: color_data = Z;
		19'b0010111010101101010: color_data = Z;
		19'b0010111010101101011: color_data = Z;
		19'b0010111010101101100: color_data = Z;
		19'b0010111010101101101: color_data = Z;
		19'b0010111010101101110: color_data = Z;
		19'b0010111010101101111: color_data = Z;
		19'b0010111010101110000: color_data = Z;
		19'b0010111010101110001: color_data = Z;
		19'b0010111010101110010: color_data = Z;
		19'b0010111010101110011: color_data = Z;
		19'b0010111010101110100: color_data = Z;
		19'b0010111010101110101: color_data = Z;
		19'b0010111010101110110: color_data = Z;
		19'b0010111010101110111: color_data = Z;
		19'b0010111010101111000: color_data = Z;
		19'b0010111010101111001: color_data = Z;
		19'b0010111010101111010: color_data = Z;
		19'b0010111010101111011: color_data = Z;
		19'b0010111010101111100: color_data = Z;
		19'b0010111010101111101: color_data = Z;
		19'b0010111010101111110: color_data = Z;
		19'b0010111010101111111: color_data = Z;
		19'b0010111010110000000: color_data = Z;
		19'b0010111010110000001: color_data = Z;
		19'b0010111010110000010: color_data = Z;
		19'b0010111010110000011: color_data = Z;
		19'b0010111010110000100: color_data = Z;
		19'b0010111010110000101: color_data = Z;
		19'b0010111010110000110: color_data = Z;
		19'b0010111010110000111: color_data = Z;
		19'b0010111010110001000: color_data = Z;
		19'b0010111010110001001: color_data = Z;
		19'b0010111010110001010: color_data = Z;
		19'b0010111010110001011: color_data = Z;
		19'b0010111010110001100: color_data = Z;
		19'b0010111010110001101: color_data = Z;
		19'b0010111010110001110: color_data = Z;
		19'b0010111010110001111: color_data = Z;
		19'b0010111010110010000: color_data = Z;
		19'b0010111010110010001: color_data = Z;
		19'b0010111010110010010: color_data = Z;
		19'b0010111010110010011: color_data = Z;
		19'b0010111010110010100: color_data = Z;
		19'b0010111010110010101: color_data = Z;
		19'b0010111010110010110: color_data = Z;
		19'b0010111010110010111: color_data = Z;
		19'b0010111010110011000: color_data = Z;
		19'b0010111010110011001: color_data = Z;
		19'b0010111010110011010: color_data = Z;
		19'b0010111010110011011: color_data = Z;
		19'b0010111010110011100: color_data = Z;
		19'b0010111010110011101: color_data = Z;
		19'b0010111010110011110: color_data = Z;
		19'b0010111010110011111: color_data = Z;
		19'b0010111010110100000: color_data = Z;
		19'b0010111010110100001: color_data = Z;
		19'b0010111010110100010: color_data = Z;
		19'b0010111010110100011: color_data = Z;
		19'b0010111010110100100: color_data = Z;
		19'b0010111010110100101: color_data = Z;
		19'b0010111010110100110: color_data = Z;
		19'b0010111010110100111: color_data = Z;
		19'b0010111010110101000: color_data = Z;
		19'b0010111010110101001: color_data = Z;
		19'b0010111010110101010: color_data = Z;
		19'b0010111010110101011: color_data = Z;
		19'b0010111010110101100: color_data = Z;
		19'b0010111010110101101: color_data = Z;
		19'b0010111010110101110: color_data = Z;
		19'b0010111010110101111: color_data = Z;
		19'b0010111010110110000: color_data = Z;
		19'b0010111010110110001: color_data = Z;
		19'b0010111010110110010: color_data = Z;
		19'b0010111010110110011: color_data = Z;
		19'b0010111010110110100: color_data = Z;
		19'b0010111010111000011: color_data = Z;
		19'b0010111010111000100: color_data = Z;
		19'b0010111010111000101: color_data = Z;
		19'b0010111010111000110: color_data = Z;
		19'b0010111010111000111: color_data = Z;
		19'b0010111010111001000: color_data = Z;
		19'b0010111010111001001: color_data = Z;
		19'b0010111010111001010: color_data = Z;
		19'b0010111010111001011: color_data = Z;
		19'b0010111010111001100: color_data = Z;
		19'b0010111010111001101: color_data = Z;
		19'b0010111010111001110: color_data = Z;
		19'b0010111010111001111: color_data = Z;
		19'b0010111100010111110: color_data = Z;
		19'b0010111100010111111: color_data = Z;
		19'b0010111100011000000: color_data = Z;
		19'b0010111100011000001: color_data = Z;
		19'b0010111100011000010: color_data = Z;
		19'b0010111100011000011: color_data = Z;
		19'b0010111100011000100: color_data = Z;
		19'b0010111100011000101: color_data = Z;
		19'b0010111100011000110: color_data = Z;
		19'b0010111100011000111: color_data = Z;
		19'b0010111100011001000: color_data = Z;
		19'b0010111100011001001: color_data = Z;
		19'b0010111100011001010: color_data = Z;
		19'b0010111100011001011: color_data = Z;
		19'b0010111100011001100: color_data = Z;
		19'b0010111100011001101: color_data = Z;
		19'b0010111100011001110: color_data = Z;
		19'b0010111100011001111: color_data = Z;
		19'b0010111100011010000: color_data = Z;
		19'b0010111100011010001: color_data = Z;
		19'b0010111100011010010: color_data = Z;
		19'b0010111100011010011: color_data = Z;
		19'b0010111100011010100: color_data = Z;
		19'b0010111100011010101: color_data = Z;
		19'b0010111100011010110: color_data = Z;
		19'b0010111100011010111: color_data = Z;
		19'b0010111100011011000: color_data = Z;
		19'b0010111100011011001: color_data = Z;
		19'b0010111100011011010: color_data = Z;
		19'b0010111100011011011: color_data = Z;
		19'b0010111100011011100: color_data = Z;
		19'b0010111100011011101: color_data = Z;
		19'b0010111100011011110: color_data = Z;
		19'b0010111100011011111: color_data = Z;
		19'b0010111100011100000: color_data = Z;
		19'b0010111100011100001: color_data = Z;
		19'b0010111100011100010: color_data = Z;
		19'b0010111100011100011: color_data = Z;
		19'b0010111100011100100: color_data = Z;
		19'b0010111100011100101: color_data = Z;
		19'b0010111100011100110: color_data = Z;
		19'b0010111100011100111: color_data = Z;
		19'b0010111100011101000: color_data = Z;
		19'b0010111100011101001: color_data = Z;
		19'b0010111100011101010: color_data = Z;
		19'b0010111100011101011: color_data = Z;
		19'b0010111100011101100: color_data = Z;
		19'b0010111100011101101: color_data = Z;
		19'b0010111100011101110: color_data = Z;
		19'b0010111100011101111: color_data = Z;
		19'b0010111100011110000: color_data = Z;
		19'b0010111100011110001: color_data = Z;
		19'b0010111100011110010: color_data = Z;
		19'b0010111100011110011: color_data = Z;
		19'b0010111100011110100: color_data = Z;
		19'b0010111100011110101: color_data = Z;
		19'b0010111100011110110: color_data = Z;
		19'b0010111100011110111: color_data = Z;
		19'b0010111100011111000: color_data = Z;
		19'b0010111100011111001: color_data = Z;
		19'b0010111100011111010: color_data = Z;
		19'b0010111100011111011: color_data = Z;
		19'b0010111100011111100: color_data = Z;
		19'b0010111100011111101: color_data = Z;
		19'b0010111100011111110: color_data = Z;
		19'b0010111100011111111: color_data = Z;
		19'b0010111100100000000: color_data = Z;
		19'b0010111100100000001: color_data = Z;
		19'b0010111100100000010: color_data = Z;
		19'b0010111100100000011: color_data = Z;
		19'b0010111100100000100: color_data = Z;
		19'b0010111100100000101: color_data = Z;
		19'b0010111100100000110: color_data = Z;
		19'b0010111100100000111: color_data = Z;
		19'b0010111100100001000: color_data = Z;
		19'b0010111100100001001: color_data = Z;
		19'b0010111100100001010: color_data = Z;
		19'b0010111100100001011: color_data = Z;
		19'b0010111100100001100: color_data = Z;
		19'b0010111100100001101: color_data = Z;
		19'b0010111100100001110: color_data = Z;
		19'b0010111100100001111: color_data = Z;
		19'b0010111100100010000: color_data = Z;
		19'b0010111100100010001: color_data = Z;
		19'b0010111100100010010: color_data = Z;
		19'b0010111100100010011: color_data = Z;
		19'b0010111100100010100: color_data = Z;
		19'b0010111100100010101: color_data = Z;
		19'b0010111100100010110: color_data = Z;
		19'b0010111100100010111: color_data = Z;
		19'b0010111100100011000: color_data = Z;
		19'b0010111100100011001: color_data = Z;
		19'b0010111100100011010: color_data = Z;
		19'b0010111100100011011: color_data = Z;
		19'b0010111100100011100: color_data = Z;
		19'b0010111100100011101: color_data = Z;
		19'b0010111100100011110: color_data = Z;
		19'b0010111100100011111: color_data = Z;
		19'b0010111100100100000: color_data = Z;
		19'b0010111100100100001: color_data = Z;
		19'b0010111100100100010: color_data = Z;
		19'b0010111100100100011: color_data = Z;
		19'b0010111100100100100: color_data = Z;
		19'b0010111100100100101: color_data = Z;
		19'b0010111100100100110: color_data = Z;
		19'b0010111100100100111: color_data = Z;
		19'b0010111100100101000: color_data = Z;
		19'b0010111100100101001: color_data = Z;
		19'b0010111100100101010: color_data = Z;
		19'b0010111100100101011: color_data = Z;
		19'b0010111100100101100: color_data = Z;
		19'b0010111100100101101: color_data = Z;
		19'b0010111100100101110: color_data = Z;
		19'b0010111100100101111: color_data = Z;
		19'b0010111100100110000: color_data = Z;
		19'b0010111100100110001: color_data = Z;
		19'b0010111100100110010: color_data = Z;
		19'b0010111100100110011: color_data = Z;
		19'b0010111100100110100: color_data = Z;
		19'b0010111100100110101: color_data = Z;
		19'b0010111100100110110: color_data = Z;
		19'b0010111100100110111: color_data = Z;
		19'b0010111100100111000: color_data = Z;
		19'b0010111100100111001: color_data = Z;
		19'b0010111100100111010: color_data = Z;
		19'b0010111100100111011: color_data = Z;
		19'b0010111100100111100: color_data = Z;
		19'b0010111100100111101: color_data = Z;
		19'b0010111100100111110: color_data = Z;
		19'b0010111100100111111: color_data = Z;
		19'b0010111100101000000: color_data = Z;
		19'b0010111100101000001: color_data = Z;
		19'b0010111100101000010: color_data = Z;
		19'b0010111100101000011: color_data = Z;
		19'b0010111100101000100: color_data = Z;
		19'b0010111100101000101: color_data = Z;
		19'b0010111100101000110: color_data = Z;
		19'b0010111100101000111: color_data = Z;
		19'b0010111100101001000: color_data = Z;
		19'b0010111100101001001: color_data = Z;
		19'b0010111100101001010: color_data = Z;
		19'b0010111100101001011: color_data = Z;
		19'b0010111100101001100: color_data = Z;
		19'b0010111100101001101: color_data = Z;
		19'b0010111100101001110: color_data = Z;
		19'b0010111100101001111: color_data = Z;
		19'b0010111100101010000: color_data = Z;
		19'b0010111100101010001: color_data = Z;
		19'b0010111100101010010: color_data = Z;
		19'b0010111100101010011: color_data = Z;
		19'b0010111100101010100: color_data = Z;
		19'b0010111100101010101: color_data = Z;
		19'b0010111100101010110: color_data = Z;
		19'b0010111100101010111: color_data = Z;
		19'b0010111100101011000: color_data = Z;
		19'b0010111100101011001: color_data = Z;
		19'b0010111100101011010: color_data = Z;
		19'b0010111100101011011: color_data = Z;
		19'b0010111100101011100: color_data = Z;
		19'b0010111100101011101: color_data = Z;
		19'b0010111100101011110: color_data = Z;
		19'b0010111100101011111: color_data = Z;
		19'b0010111100101100000: color_data = Z;
		19'b0010111100101100001: color_data = Z;
		19'b0010111100101100010: color_data = Z;
		19'b0010111100101100011: color_data = Z;
		19'b0010111100101100100: color_data = Z;
		19'b0010111100101100101: color_data = Z;
		19'b0010111100101100110: color_data = Z;
		19'b0010111100101100111: color_data = Z;
		19'b0010111100101101000: color_data = Z;
		19'b0010111100101101001: color_data = Z;
		19'b0010111100101101010: color_data = Z;
		19'b0010111100101101011: color_data = Z;
		19'b0010111100101101100: color_data = Z;
		19'b0010111100101101101: color_data = Z;
		19'b0010111100101101110: color_data = Z;
		19'b0010111100101101111: color_data = Z;
		19'b0010111100101110000: color_data = Z;
		19'b0010111100101110001: color_data = Z;
		19'b0010111100101110010: color_data = Z;
		19'b0010111100101110011: color_data = Z;
		19'b0010111100101110100: color_data = Z;
		19'b0010111100101110101: color_data = Z;
		19'b0010111100101110110: color_data = Z;
		19'b0010111100101110111: color_data = Z;
		19'b0010111100101111000: color_data = Z;
		19'b0010111100101111001: color_data = Z;
		19'b0010111100101111010: color_data = Z;
		19'b0010111100101111011: color_data = Z;
		19'b0010111100101111100: color_data = Z;
		19'b0010111100101111101: color_data = Z;
		19'b0010111100101111110: color_data = Z;
		19'b0010111100101111111: color_data = Z;
		19'b0010111100110000000: color_data = Z;
		19'b0010111100110000001: color_data = Z;
		19'b0010111100110000010: color_data = Z;
		19'b0010111100110000011: color_data = Z;
		19'b0010111100110000100: color_data = Z;
		19'b0010111100110000101: color_data = Z;
		19'b0010111100110000110: color_data = Z;
		19'b0010111100110000111: color_data = Z;
		19'b0010111100110001000: color_data = Z;
		19'b0010111100110001001: color_data = Z;
		19'b0010111100110001010: color_data = Z;
		19'b0010111100110001011: color_data = Z;
		19'b0010111100110001100: color_data = Z;
		19'b0010111100110001101: color_data = Z;
		19'b0010111100110001110: color_data = Z;
		19'b0010111100110001111: color_data = Z;
		19'b0010111100110010000: color_data = Z;
		19'b0010111100110010001: color_data = Z;
		19'b0010111100110010010: color_data = Z;
		19'b0010111100110010011: color_data = Z;
		19'b0010111100110010100: color_data = Z;
		19'b0010111100110010101: color_data = Z;
		19'b0010111100110010110: color_data = Z;
		19'b0010111100110010111: color_data = Z;
		19'b0010111100110011000: color_data = Z;
		19'b0010111100110011001: color_data = Z;
		19'b0010111100110011010: color_data = Z;
		19'b0010111100110011011: color_data = Z;
		19'b0010111100110011100: color_data = Z;
		19'b0010111100110011101: color_data = Z;
		19'b0010111100110011110: color_data = Z;
		19'b0010111100110011111: color_data = Z;
		19'b0010111100110100000: color_data = Z;
		19'b0010111100110100001: color_data = Z;
		19'b0010111100110100010: color_data = Z;
		19'b0010111100110100011: color_data = Z;
		19'b0010111100110100100: color_data = Z;
		19'b0010111100110100101: color_data = Z;
		19'b0010111100110100110: color_data = Z;
		19'b0010111100110100111: color_data = Z;
		19'b0010111100110101000: color_data = Z;
		19'b0010111100110101001: color_data = Z;
		19'b0010111100110101010: color_data = Z;
		19'b0010111100110101011: color_data = Z;
		19'b0010111100110101100: color_data = Z;
		19'b0010111100110101101: color_data = Z;
		19'b0010111100110101110: color_data = Z;
		19'b0010111100110101111: color_data = Z;
		19'b0010111100110110000: color_data = Z;
		19'b0010111100110110001: color_data = Z;
		19'b0010111100110110010: color_data = Z;
		19'b0010111100110110011: color_data = Z;
		19'b0010111100110110100: color_data = Z;
		19'b0010111100111000100: color_data = Z;
		19'b0010111100111000101: color_data = Z;
		19'b0010111100111000110: color_data = Z;
		19'b0010111100111000111: color_data = Z;
		19'b0010111100111001000: color_data = Z;
		19'b0010111100111001001: color_data = Z;
		19'b0010111100111001010: color_data = Z;
		19'b0010111100111001011: color_data = Z;
		19'b0010111100111001100: color_data = Z;
		19'b0010111100111001101: color_data = Z;
		19'b0010111100111001110: color_data = Z;
		19'b0010111100111001111: color_data = Z;
		19'b0010111110010111101: color_data = Z;
		19'b0010111110010111110: color_data = Z;
		19'b0010111110010111111: color_data = Z;
		19'b0010111110011000000: color_data = Z;
		19'b0010111110011000001: color_data = Z;
		19'b0010111110011000010: color_data = Z;
		19'b0010111110011000011: color_data = Z;
		19'b0010111110011000100: color_data = Z;
		19'b0010111110011000101: color_data = Z;
		19'b0010111110011000110: color_data = Z;
		19'b0010111110011000111: color_data = Z;
		19'b0010111110011001000: color_data = Z;
		19'b0010111110011001001: color_data = Z;
		19'b0010111110011001010: color_data = Z;
		19'b0010111110011001011: color_data = Z;
		19'b0010111110011001100: color_data = Z;
		19'b0010111110011001101: color_data = Z;
		19'b0010111110011001110: color_data = Z;
		19'b0010111110011001111: color_data = Z;
		19'b0010111110011010000: color_data = Z;
		19'b0010111110011010001: color_data = Z;
		19'b0010111110011010010: color_data = Z;
		19'b0010111110011010011: color_data = Z;
		19'b0010111110011010100: color_data = Z;
		19'b0010111110011010101: color_data = Z;
		19'b0010111110011010110: color_data = Z;
		19'b0010111110011010111: color_data = Z;
		19'b0010111110011011000: color_data = Z;
		19'b0010111110011011001: color_data = Z;
		19'b0010111110011011010: color_data = Z;
		19'b0010111110011011011: color_data = Z;
		19'b0010111110011011100: color_data = Z;
		19'b0010111110011011101: color_data = Z;
		19'b0010111110011011110: color_data = Z;
		19'b0010111110011011111: color_data = Z;
		19'b0010111110011100000: color_data = Z;
		19'b0010111110011100001: color_data = Z;
		19'b0010111110011100010: color_data = Z;
		19'b0010111110011100011: color_data = Z;
		19'b0010111110011100100: color_data = Z;
		19'b0010111110011100101: color_data = Z;
		19'b0010111110011100110: color_data = Z;
		19'b0010111110011100111: color_data = Z;
		19'b0010111110011101000: color_data = Z;
		19'b0010111110011101001: color_data = Z;
		19'b0010111110011101010: color_data = Z;
		19'b0010111110011101011: color_data = Z;
		19'b0010111110011101100: color_data = Z;
		19'b0010111110011101101: color_data = Z;
		19'b0010111110011101110: color_data = Z;
		19'b0010111110011101111: color_data = Z;
		19'b0010111110011110000: color_data = Z;
		19'b0010111110011110001: color_data = Z;
		19'b0010111110011110010: color_data = Z;
		19'b0010111110011110011: color_data = Z;
		19'b0010111110011110100: color_data = Z;
		19'b0010111110011110101: color_data = Z;
		19'b0010111110011110110: color_data = Z;
		19'b0010111110011110111: color_data = Z;
		19'b0010111110011111000: color_data = Z;
		19'b0010111110011111001: color_data = Z;
		19'b0010111110011111010: color_data = Z;
		19'b0010111110011111011: color_data = Z;
		19'b0010111110011111100: color_data = Z;
		19'b0010111110011111101: color_data = Z;
		19'b0010111110011111110: color_data = Z;
		19'b0010111110011111111: color_data = Z;
		19'b0010111110100000000: color_data = Z;
		19'b0010111110100000001: color_data = Z;
		19'b0010111110100000010: color_data = Z;
		19'b0010111110100000011: color_data = Z;
		19'b0010111110100000100: color_data = Z;
		19'b0010111110100000101: color_data = Z;
		19'b0010111110100000110: color_data = Z;
		19'b0010111110100000111: color_data = Z;
		19'b0010111110100001000: color_data = Z;
		19'b0010111110100001001: color_data = Z;
		19'b0010111110100001010: color_data = Z;
		19'b0010111110100001011: color_data = Z;
		19'b0010111110100001100: color_data = Z;
		19'b0010111110100001101: color_data = Z;
		19'b0010111110100001110: color_data = Z;
		19'b0010111110100001111: color_data = Z;
		19'b0010111110100010000: color_data = Z;
		19'b0010111110100010001: color_data = Z;
		19'b0010111110100010010: color_data = Z;
		19'b0010111110100010011: color_data = Z;
		19'b0010111110100010100: color_data = Z;
		19'b0010111110100010101: color_data = Z;
		19'b0010111110100010110: color_data = Z;
		19'b0010111110100010111: color_data = Z;
		19'b0010111110100011000: color_data = Z;
		19'b0010111110100011001: color_data = Z;
		19'b0010111110100011010: color_data = Z;
		19'b0010111110100011011: color_data = Z;
		19'b0010111110100011100: color_data = Z;
		19'b0010111110100011101: color_data = Z;
		19'b0010111110100011110: color_data = Z;
		19'b0010111110100011111: color_data = Z;
		19'b0010111110100100000: color_data = Z;
		19'b0010111110100100001: color_data = Z;
		19'b0010111110100100010: color_data = Z;
		19'b0010111110100100011: color_data = Z;
		19'b0010111110100100100: color_data = Z;
		19'b0010111110100100101: color_data = Z;
		19'b0010111110100100110: color_data = Z;
		19'b0010111110100100111: color_data = Z;
		19'b0010111110100101000: color_data = Z;
		19'b0010111110100101001: color_data = Z;
		19'b0010111110100101010: color_data = Z;
		19'b0010111110100101011: color_data = Z;
		19'b0010111110100101100: color_data = Z;
		19'b0010111110100101101: color_data = Z;
		19'b0010111110100101110: color_data = Z;
		19'b0010111110100101111: color_data = Z;
		19'b0010111110100110000: color_data = Z;
		19'b0010111110100110001: color_data = Z;
		19'b0010111110100110010: color_data = Z;
		19'b0010111110100110011: color_data = Z;
		19'b0010111110100110100: color_data = Z;
		19'b0010111110100110101: color_data = Z;
		19'b0010111110100110110: color_data = Z;
		19'b0010111110100110111: color_data = Z;
		19'b0010111110100111000: color_data = Z;
		19'b0010111110100111001: color_data = Z;
		19'b0010111110100111010: color_data = Z;
		19'b0010111110100111011: color_data = Z;
		19'b0010111110100111100: color_data = Z;
		19'b0010111110100111101: color_data = Z;
		19'b0010111110100111110: color_data = Z;
		19'b0010111110100111111: color_data = Z;
		19'b0010111110101000000: color_data = Z;
		19'b0010111110101000001: color_data = Z;
		19'b0010111110101000010: color_data = Z;
		19'b0010111110101000011: color_data = Z;
		19'b0010111110101000100: color_data = Z;
		19'b0010111110101000101: color_data = Z;
		19'b0010111110101000110: color_data = Z;
		19'b0010111110101000111: color_data = Z;
		19'b0010111110101001000: color_data = Z;
		19'b0010111110101001001: color_data = Z;
		19'b0010111110101001010: color_data = Z;
		19'b0010111110101001011: color_data = Z;
		19'b0010111110101001100: color_data = Z;
		19'b0010111110101001101: color_data = Z;
		19'b0010111110101001110: color_data = Z;
		19'b0010111110101001111: color_data = Z;
		19'b0010111110101010000: color_data = Z;
		19'b0010111110101010001: color_data = Z;
		19'b0010111110101010010: color_data = Z;
		19'b0010111110101010011: color_data = Z;
		19'b0010111110101010100: color_data = Z;
		19'b0010111110101010101: color_data = Z;
		19'b0010111110101010110: color_data = Z;
		19'b0010111110101010111: color_data = Z;
		19'b0010111110101011000: color_data = Z;
		19'b0010111110101011001: color_data = Z;
		19'b0010111110101011010: color_data = Z;
		19'b0010111110101011011: color_data = Z;
		19'b0010111110101011100: color_data = Z;
		19'b0010111110101011101: color_data = Z;
		19'b0010111110101011110: color_data = Z;
		19'b0010111110101011111: color_data = Z;
		19'b0010111110101100000: color_data = Z;
		19'b0010111110101100001: color_data = Z;
		19'b0010111110101100010: color_data = Z;
		19'b0010111110101100011: color_data = Z;
		19'b0010111110101100100: color_data = Z;
		19'b0010111110101100101: color_data = Z;
		19'b0010111110101100110: color_data = Z;
		19'b0010111110101100111: color_data = Z;
		19'b0010111110101101000: color_data = Z;
		19'b0010111110101101001: color_data = Z;
		19'b0010111110101101010: color_data = Z;
		19'b0010111110101101011: color_data = Z;
		19'b0010111110101101100: color_data = Z;
		19'b0010111110101101101: color_data = Z;
		19'b0010111110101101110: color_data = Z;
		19'b0010111110101101111: color_data = Z;
		19'b0010111110101110000: color_data = Z;
		19'b0010111110101110001: color_data = Z;
		19'b0010111110101110010: color_data = Z;
		19'b0010111110101110011: color_data = Z;
		19'b0010111110101110100: color_data = Z;
		19'b0010111110101110101: color_data = Z;
		19'b0010111110101110110: color_data = Z;
		19'b0010111110101110111: color_data = Z;
		19'b0010111110101111000: color_data = Z;
		19'b0010111110101111001: color_data = Z;
		19'b0010111110101111010: color_data = Z;
		19'b0010111110101111011: color_data = Z;
		19'b0010111110101111100: color_data = Z;
		19'b0010111110101111101: color_data = Z;
		19'b0010111110101111110: color_data = Z;
		19'b0010111110101111111: color_data = Z;
		19'b0010111110110000000: color_data = Z;
		19'b0010111110110000001: color_data = Z;
		19'b0010111110110000010: color_data = Z;
		19'b0010111110110000011: color_data = Z;
		19'b0010111110110000100: color_data = Z;
		19'b0010111110110000101: color_data = Z;
		19'b0010111110110000110: color_data = Z;
		19'b0010111110110000111: color_data = Z;
		19'b0010111110110001000: color_data = Z;
		19'b0010111110110001001: color_data = Z;
		19'b0010111110110001010: color_data = Z;
		19'b0010111110110001011: color_data = Z;
		19'b0010111110110001100: color_data = Z;
		19'b0010111110110001101: color_data = Z;
		19'b0010111110110001110: color_data = Z;
		19'b0010111110110001111: color_data = Z;
		19'b0010111110110010000: color_data = Z;
		19'b0010111110110010001: color_data = Z;
		19'b0010111110110010010: color_data = Z;
		19'b0010111110110010011: color_data = Z;
		19'b0010111110110010100: color_data = Z;
		19'b0010111110110010101: color_data = Z;
		19'b0010111110110010110: color_data = Z;
		19'b0010111110110010111: color_data = Z;
		19'b0010111110110011000: color_data = Z;
		19'b0010111110110011001: color_data = Z;
		19'b0010111110110011010: color_data = Z;
		19'b0010111110110011011: color_data = Z;
		19'b0010111110110011100: color_data = Z;
		19'b0010111110110011101: color_data = Z;
		19'b0010111110110011110: color_data = Z;
		19'b0010111110110011111: color_data = Z;
		19'b0010111110110100000: color_data = Z;
		19'b0010111110110100001: color_data = Z;
		19'b0010111110110100010: color_data = Z;
		19'b0010111110110100011: color_data = Z;
		19'b0010111110110100100: color_data = Z;
		19'b0010111110110100101: color_data = Z;
		19'b0010111110110100110: color_data = Z;
		19'b0010111110110100111: color_data = Z;
		19'b0010111110110101000: color_data = Z;
		19'b0010111110110101001: color_data = Z;
		19'b0010111110110101010: color_data = Z;
		19'b0010111110110101011: color_data = Z;
		19'b0010111110110101100: color_data = Z;
		19'b0010111110110101101: color_data = Z;
		19'b0010111110110101110: color_data = Z;
		19'b0010111110110101111: color_data = Z;
		19'b0010111110110110000: color_data = Z;
		19'b0010111110110110001: color_data = Z;
		19'b0010111110110110010: color_data = Z;
		19'b0010111110110110011: color_data = Z;
		19'b0010111110110110100: color_data = Z;
		19'b0010111110111000101: color_data = Z;
		19'b0010111110111000110: color_data = Z;
		19'b0010111110111000111: color_data = Z;
		19'b0010111110111001000: color_data = Z;
		19'b0010111110111001001: color_data = Z;
		19'b0010111110111001010: color_data = Z;
		19'b0010111110111001011: color_data = Z;
		19'b0010111110111001100: color_data = Z;
		19'b0010111110111001101: color_data = Z;
		19'b0010111110111001110: color_data = Z;
		19'b0010111110111001111: color_data = Z;
		19'b0010111110111010000: color_data = Z;
		19'b0011000000010111100: color_data = Z;
		19'b0011000000010111101: color_data = Z;
		19'b0011000000010111110: color_data = Z;
		19'b0011000000010111111: color_data = Z;
		19'b0011000000011000000: color_data = Z;
		19'b0011000000011000001: color_data = Z;
		19'b0011000000011000010: color_data = Z;
		19'b0011000000011000011: color_data = Z;
		19'b0011000000011000100: color_data = Z;
		19'b0011000000011000101: color_data = Z;
		19'b0011000000011000110: color_data = Z;
		19'b0011000000011000111: color_data = Z;
		19'b0011000000011001000: color_data = Z;
		19'b0011000000011001001: color_data = Z;
		19'b0011000000011001010: color_data = Z;
		19'b0011000000011001011: color_data = Z;
		19'b0011000000011001100: color_data = Z;
		19'b0011000000011001101: color_data = Z;
		19'b0011000000011001110: color_data = Z;
		19'b0011000000011001111: color_data = Z;
		19'b0011000000011010000: color_data = Z;
		19'b0011000000011010001: color_data = Z;
		19'b0011000000011010010: color_data = Z;
		19'b0011000000011010011: color_data = Z;
		19'b0011000000011010100: color_data = Z;
		19'b0011000000011010101: color_data = Z;
		19'b0011000000011010110: color_data = Z;
		19'b0011000000011010111: color_data = Z;
		19'b0011000000011011000: color_data = Z;
		19'b0011000000011011001: color_data = Z;
		19'b0011000000011011010: color_data = Z;
		19'b0011000000011011011: color_data = Z;
		19'b0011000000011011100: color_data = Z;
		19'b0011000000011011101: color_data = Z;
		19'b0011000000011011110: color_data = Z;
		19'b0011000000011011111: color_data = Z;
		19'b0011000000011100000: color_data = Z;
		19'b0011000000011100001: color_data = Z;
		19'b0011000000011100010: color_data = Z;
		19'b0011000000011100011: color_data = Z;
		19'b0011000000011100100: color_data = Z;
		19'b0011000000011100101: color_data = Z;
		19'b0011000000011100110: color_data = Z;
		19'b0011000000011100111: color_data = Z;
		19'b0011000000011101000: color_data = Z;
		19'b0011000000011101001: color_data = Z;
		19'b0011000000011101010: color_data = Z;
		19'b0011000000011101011: color_data = Z;
		19'b0011000000011101100: color_data = Z;
		19'b0011000000011101101: color_data = Z;
		19'b0011000000011101110: color_data = Z;
		19'b0011000000011101111: color_data = Z;
		19'b0011000000011110000: color_data = Z;
		19'b0011000000011110001: color_data = Z;
		19'b0011000000011110010: color_data = Z;
		19'b0011000000011110011: color_data = Z;
		19'b0011000000011110100: color_data = Z;
		19'b0011000000011110101: color_data = Z;
		19'b0011000000011110110: color_data = Z;
		19'b0011000000011110111: color_data = Z;
		19'b0011000000011111000: color_data = Z;
		19'b0011000000011111001: color_data = Z;
		19'b0011000000011111010: color_data = Z;
		19'b0011000000011111011: color_data = Z;
		19'b0011000000011111100: color_data = Z;
		19'b0011000000011111101: color_data = Z;
		19'b0011000000011111110: color_data = Z;
		19'b0011000000011111111: color_data = Z;
		19'b0011000000100000000: color_data = Z;
		19'b0011000000100000001: color_data = Z;
		19'b0011000000100000010: color_data = Z;
		19'b0011000000100000011: color_data = Z;
		19'b0011000000100000100: color_data = Z;
		19'b0011000000100000101: color_data = Z;
		19'b0011000000100000110: color_data = Z;
		19'b0011000000100000111: color_data = Z;
		19'b0011000000100001000: color_data = Z;
		19'b0011000000100001001: color_data = Z;
		19'b0011000000100001010: color_data = Z;
		19'b0011000000100001011: color_data = Z;
		19'b0011000000100001100: color_data = Z;
		19'b0011000000100001101: color_data = Z;
		19'b0011000000100001110: color_data = Z;
		19'b0011000000100001111: color_data = Z;
		19'b0011000000100010000: color_data = Z;
		19'b0011000000100010001: color_data = Z;
		19'b0011000000100010010: color_data = Z;
		19'b0011000000100010011: color_data = Z;
		19'b0011000000100010100: color_data = Z;
		19'b0011000000100010101: color_data = Z;
		19'b0011000000100010110: color_data = Z;
		19'b0011000000100010111: color_data = Z;
		19'b0011000000100011000: color_data = Z;
		19'b0011000000100011001: color_data = Z;
		19'b0011000000100011010: color_data = Z;
		19'b0011000000100011011: color_data = Z;
		19'b0011000000100011100: color_data = Z;
		19'b0011000000100011101: color_data = Z;
		19'b0011000000100011110: color_data = Z;
		19'b0011000000100011111: color_data = Z;
		19'b0011000000100100000: color_data = Z;
		19'b0011000000100100001: color_data = Z;
		19'b0011000000100100010: color_data = Z;
		19'b0011000000100100011: color_data = Z;
		19'b0011000000100100100: color_data = Z;
		19'b0011000000100100101: color_data = Z;
		19'b0011000000100100110: color_data = Z;
		19'b0011000000100100111: color_data = Z;
		19'b0011000000100101000: color_data = Z;
		19'b0011000000100101001: color_data = Z;
		19'b0011000000100101010: color_data = Z;
		19'b0011000000100101011: color_data = Z;
		19'b0011000000100101100: color_data = Z;
		19'b0011000000100101101: color_data = Z;
		19'b0011000000100101110: color_data = Z;
		19'b0011000000100101111: color_data = Z;
		19'b0011000000100110000: color_data = Z;
		19'b0011000000100110001: color_data = Z;
		19'b0011000000100110010: color_data = Z;
		19'b0011000000100110011: color_data = Z;
		19'b0011000000100110100: color_data = Z;
		19'b0011000000100110101: color_data = Z;
		19'b0011000000100110110: color_data = Z;
		19'b0011000000100110111: color_data = Z;
		19'b0011000000100111000: color_data = Z;
		19'b0011000000100111001: color_data = Z;
		19'b0011000000100111010: color_data = Z;
		19'b0011000000100111011: color_data = Z;
		19'b0011000000100111100: color_data = Z;
		19'b0011000000100111101: color_data = Z;
		19'b0011000000100111110: color_data = Z;
		19'b0011000000100111111: color_data = Z;
		19'b0011000000101000000: color_data = Z;
		19'b0011000000101000001: color_data = Z;
		19'b0011000000101000010: color_data = Z;
		19'b0011000000101000011: color_data = Z;
		19'b0011000000101000100: color_data = Z;
		19'b0011000000101000101: color_data = Z;
		19'b0011000000101000110: color_data = Z;
		19'b0011000000101000111: color_data = Z;
		19'b0011000000101001000: color_data = Z;
		19'b0011000000101001001: color_data = Z;
		19'b0011000000101001010: color_data = Z;
		19'b0011000000101001011: color_data = Z;
		19'b0011000000101001100: color_data = Z;
		19'b0011000000101001101: color_data = Z;
		19'b0011000000101001110: color_data = Z;
		19'b0011000000101001111: color_data = Z;
		19'b0011000000101010000: color_data = Z;
		19'b0011000000101010001: color_data = Z;
		19'b0011000000101010010: color_data = Z;
		19'b0011000000101010011: color_data = Z;
		19'b0011000000101010100: color_data = Z;
		19'b0011000000101010101: color_data = Z;
		19'b0011000000101010110: color_data = Z;
		19'b0011000000101010111: color_data = Z;
		19'b0011000000101011000: color_data = Z;
		19'b0011000000101011001: color_data = Z;
		19'b0011000000101011010: color_data = Z;
		19'b0011000000101011011: color_data = Z;
		19'b0011000000101011100: color_data = Z;
		19'b0011000000101011101: color_data = Z;
		19'b0011000000101011110: color_data = Z;
		19'b0011000000101011111: color_data = Z;
		19'b0011000000101100000: color_data = Z;
		19'b0011000000101100001: color_data = Z;
		19'b0011000000101100010: color_data = Z;
		19'b0011000000101100011: color_data = Z;
		19'b0011000000101100100: color_data = Z;
		19'b0011000000101100101: color_data = Z;
		19'b0011000000101100110: color_data = Z;
		19'b0011000000101100111: color_data = Z;
		19'b0011000000101101000: color_data = Z;
		19'b0011000000101101001: color_data = Z;
		19'b0011000000101101010: color_data = Z;
		19'b0011000000101101011: color_data = Z;
		19'b0011000000101101100: color_data = Z;
		19'b0011000000101101101: color_data = Z;
		19'b0011000000101101110: color_data = Z;
		19'b0011000000101101111: color_data = Z;
		19'b0011000000101110000: color_data = Z;
		19'b0011000000101110001: color_data = Z;
		19'b0011000000101110010: color_data = Z;
		19'b0011000000101110011: color_data = Z;
		19'b0011000000101110100: color_data = Z;
		19'b0011000000101110101: color_data = Z;
		19'b0011000000101110110: color_data = Z;
		19'b0011000000101110111: color_data = Z;
		19'b0011000000101111000: color_data = Z;
		19'b0011000000101111001: color_data = Z;
		19'b0011000000101111010: color_data = Z;
		19'b0011000000101111011: color_data = Z;
		19'b0011000000101111100: color_data = Z;
		19'b0011000000101111101: color_data = Z;
		19'b0011000000101111110: color_data = Z;
		19'b0011000000101111111: color_data = Z;
		19'b0011000000110000000: color_data = Z;
		19'b0011000000110000001: color_data = Z;
		19'b0011000000110000010: color_data = Z;
		19'b0011000000110000011: color_data = Z;
		19'b0011000000110000100: color_data = Z;
		19'b0011000000110000101: color_data = Z;
		19'b0011000000110000110: color_data = Z;
		19'b0011000000110000111: color_data = Z;
		19'b0011000000110001000: color_data = Z;
		19'b0011000000110001001: color_data = Z;
		19'b0011000000110001010: color_data = Z;
		19'b0011000000110001011: color_data = Z;
		19'b0011000000110001100: color_data = Z;
		19'b0011000000110001101: color_data = Z;
		19'b0011000000110001110: color_data = Z;
		19'b0011000000110001111: color_data = Z;
		19'b0011000000110010000: color_data = Z;
		19'b0011000000110010001: color_data = Z;
		19'b0011000000110010010: color_data = Z;
		19'b0011000000110010011: color_data = Z;
		19'b0011000000110010100: color_data = Z;
		19'b0011000000110010101: color_data = Z;
		19'b0011000000110010110: color_data = Z;
		19'b0011000000110010111: color_data = Z;
		19'b0011000000110011000: color_data = Z;
		19'b0011000000110011001: color_data = Z;
		19'b0011000000110011010: color_data = Z;
		19'b0011000000110011011: color_data = Z;
		19'b0011000000110011100: color_data = Z;
		19'b0011000000110011101: color_data = Z;
		19'b0011000000110011110: color_data = Z;
		19'b0011000000110011111: color_data = Z;
		19'b0011000000110100000: color_data = Z;
		19'b0011000000110100001: color_data = Z;
		19'b0011000000110100010: color_data = Z;
		19'b0011000000110100011: color_data = Z;
		19'b0011000000110100100: color_data = Z;
		19'b0011000000110100101: color_data = Z;
		19'b0011000000110100110: color_data = Z;
		19'b0011000000110100111: color_data = Z;
		19'b0011000000110101000: color_data = Z;
		19'b0011000000110101001: color_data = Z;
		19'b0011000000110101010: color_data = Z;
		19'b0011000000110101011: color_data = Z;
		19'b0011000000110101100: color_data = Z;
		19'b0011000000110101101: color_data = Z;
		19'b0011000000110101110: color_data = Z;
		19'b0011000000110101111: color_data = Z;
		19'b0011000000110110000: color_data = Z;
		19'b0011000000110110001: color_data = Z;
		19'b0011000000110110010: color_data = Z;
		19'b0011000000110110011: color_data = Z;
		19'b0011000000110110100: color_data = Z;
		19'b0011000000110110101: color_data = Z;
		19'b0011000000111000110: color_data = Z;
		19'b0011000000111000111: color_data = Z;
		19'b0011000000111001000: color_data = Z;
		19'b0011000000111001001: color_data = Z;
		19'b0011000000111001010: color_data = Z;
		19'b0011000000111001011: color_data = Z;
		19'b0011000000111001100: color_data = Z;
		19'b0011000000111001101: color_data = Z;
		19'b0011000000111001110: color_data = Z;
		19'b0011000000111001111: color_data = Z;
		19'b0011000010010111011: color_data = Z;
		19'b0011000010010111100: color_data = Z;
		19'b0011000010010111101: color_data = Z;
		19'b0011000010010111110: color_data = Z;
		19'b0011000010010111111: color_data = Z;
		19'b0011000010011000000: color_data = Z;
		19'b0011000010011000001: color_data = Z;
		19'b0011000010011000010: color_data = Z;
		19'b0011000010011000011: color_data = Z;
		19'b0011000010011000100: color_data = Z;
		19'b0011000010011000101: color_data = Z;
		19'b0011000010011000110: color_data = Z;
		19'b0011000010011000111: color_data = Z;
		19'b0011000010011001000: color_data = Z;
		19'b0011000010011001001: color_data = Z;
		19'b0011000010011001010: color_data = Z;
		19'b0011000010011001011: color_data = Z;
		19'b0011000010011001100: color_data = Z;
		19'b0011000010011001101: color_data = Z;
		19'b0011000010011001110: color_data = Z;
		19'b0011000010011001111: color_data = Z;
		19'b0011000010011010000: color_data = Z;
		19'b0011000010011010001: color_data = Z;
		19'b0011000010011010010: color_data = Z;
		19'b0011000010011010011: color_data = Z;
		19'b0011000010011010100: color_data = Z;
		19'b0011000010011010101: color_data = Z;
		19'b0011000010011010110: color_data = Z;
		19'b0011000010011010111: color_data = Z;
		19'b0011000010011011000: color_data = Z;
		19'b0011000010011011001: color_data = Z;
		19'b0011000010011011010: color_data = Z;
		19'b0011000010011011011: color_data = Z;
		19'b0011000010011011100: color_data = Z;
		19'b0011000010011011101: color_data = Z;
		19'b0011000010011011110: color_data = Z;
		19'b0011000010011011111: color_data = Z;
		19'b0011000010011100000: color_data = Z;
		19'b0011000010011100001: color_data = Z;
		19'b0011000010011100010: color_data = Z;
		19'b0011000010011100011: color_data = Z;
		19'b0011000010011100100: color_data = Z;
		19'b0011000010011100101: color_data = Z;
		19'b0011000010011100110: color_data = Z;
		19'b0011000010011100111: color_data = Z;
		19'b0011000010011101000: color_data = Z;
		19'b0011000010011101001: color_data = Z;
		19'b0011000010011101010: color_data = Z;
		19'b0011000010011101011: color_data = Z;
		19'b0011000010011101100: color_data = Z;
		19'b0011000010011101101: color_data = Z;
		19'b0011000010011101110: color_data = Z;
		19'b0011000010011101111: color_data = Z;
		19'b0011000010011110000: color_data = Z;
		19'b0011000010011110001: color_data = Z;
		19'b0011000010011110010: color_data = Z;
		19'b0011000010011110011: color_data = Z;
		19'b0011000010011110100: color_data = Z;
		19'b0011000010011110101: color_data = Z;
		19'b0011000010011110110: color_data = Z;
		19'b0011000010011110111: color_data = Z;
		19'b0011000010011111000: color_data = Z;
		19'b0011000010011111001: color_data = Z;
		19'b0011000010011111010: color_data = Z;
		19'b0011000010011111011: color_data = Z;
		19'b0011000010011111100: color_data = Z;
		19'b0011000010011111101: color_data = Z;
		19'b0011000010011111110: color_data = Z;
		19'b0011000010011111111: color_data = Z;
		19'b0011000010100000000: color_data = Z;
		19'b0011000010100000001: color_data = Z;
		19'b0011000010100000010: color_data = Z;
		19'b0011000010100000011: color_data = Z;
		19'b0011000010100000100: color_data = Z;
		19'b0011000010100000101: color_data = Z;
		19'b0011000010100000110: color_data = Z;
		19'b0011000010100000111: color_data = Z;
		19'b0011000010100001000: color_data = Z;
		19'b0011000010100001001: color_data = Z;
		19'b0011000010100001010: color_data = Z;
		19'b0011000010100001011: color_data = Z;
		19'b0011000010100001100: color_data = Z;
		19'b0011000010100001101: color_data = Z;
		19'b0011000010100001110: color_data = Z;
		19'b0011000010100001111: color_data = Z;
		19'b0011000010100010000: color_data = Z;
		19'b0011000010100010001: color_data = Z;
		19'b0011000010100010010: color_data = Z;
		19'b0011000010100010011: color_data = Z;
		19'b0011000010100010100: color_data = Z;
		19'b0011000010100010101: color_data = Z;
		19'b0011000010100010110: color_data = Z;
		19'b0011000010100010111: color_data = Z;
		19'b0011000010100011000: color_data = Z;
		19'b0011000010100011001: color_data = Z;
		19'b0011000010100011010: color_data = Z;
		19'b0011000010100011011: color_data = Z;
		19'b0011000010100011100: color_data = Z;
		19'b0011000010100011101: color_data = Z;
		19'b0011000010100011110: color_data = Z;
		19'b0011000010100011111: color_data = Z;
		19'b0011000010100100000: color_data = Z;
		19'b0011000010100100001: color_data = Z;
		19'b0011000010100100010: color_data = Z;
		19'b0011000010100100011: color_data = Z;
		19'b0011000010100100100: color_data = Z;
		19'b0011000010100100101: color_data = Z;
		19'b0011000010100100110: color_data = Z;
		19'b0011000010100100111: color_data = Z;
		19'b0011000010100101000: color_data = Z;
		19'b0011000010100101001: color_data = Z;
		19'b0011000010100101010: color_data = Z;
		19'b0011000010100101011: color_data = Z;
		19'b0011000010100101100: color_data = Z;
		19'b0011000010100101101: color_data = Z;
		19'b0011000010100101110: color_data = Z;
		19'b0011000010100101111: color_data = Z;
		19'b0011000010100110000: color_data = Z;
		19'b0011000010100110001: color_data = Z;
		19'b0011000010100110010: color_data = Z;
		19'b0011000010100110011: color_data = Z;
		19'b0011000010100110100: color_data = Z;
		19'b0011000010100110101: color_data = Z;
		19'b0011000010100110110: color_data = Z;
		19'b0011000010100110111: color_data = Z;
		19'b0011000010100111000: color_data = Z;
		19'b0011000010100111001: color_data = Z;
		19'b0011000010100111010: color_data = Z;
		19'b0011000010100111011: color_data = Z;
		19'b0011000010100111100: color_data = Z;
		19'b0011000010100111101: color_data = Z;
		19'b0011000010100111110: color_data = Z;
		19'b0011000010100111111: color_data = Z;
		19'b0011000010101000000: color_data = Z;
		19'b0011000010101000001: color_data = Z;
		19'b0011000010101000010: color_data = Z;
		19'b0011000010101000011: color_data = Z;
		19'b0011000010101000100: color_data = Z;
		19'b0011000010101000101: color_data = Z;
		19'b0011000010101000110: color_data = Z;
		19'b0011000010101000111: color_data = Z;
		19'b0011000010101001000: color_data = Z;
		19'b0011000010101001001: color_data = Z;
		19'b0011000010101001010: color_data = Z;
		19'b0011000010101001011: color_data = Z;
		19'b0011000010101001100: color_data = Z;
		19'b0011000010101001101: color_data = Z;
		19'b0011000010101001110: color_data = Z;
		19'b0011000010101001111: color_data = Z;
		19'b0011000010101010000: color_data = Z;
		19'b0011000010101010001: color_data = Z;
		19'b0011000010101010010: color_data = Z;
		19'b0011000010101010011: color_data = Z;
		19'b0011000010101010100: color_data = Z;
		19'b0011000010101010101: color_data = Z;
		19'b0011000010101010110: color_data = Z;
		19'b0011000010101010111: color_data = Z;
		19'b0011000010101011000: color_data = Z;
		19'b0011000010101011001: color_data = Z;
		19'b0011000010101011010: color_data = Z;
		19'b0011000010101011011: color_data = Z;
		19'b0011000010101011100: color_data = Z;
		19'b0011000010101011101: color_data = Z;
		19'b0011000010101011110: color_data = Z;
		19'b0011000010101011111: color_data = Z;
		19'b0011000010101100000: color_data = Z;
		19'b0011000010101100001: color_data = Z;
		19'b0011000010101100010: color_data = Z;
		19'b0011000010101100011: color_data = Z;
		19'b0011000010101100100: color_data = Z;
		19'b0011000010101100101: color_data = Z;
		19'b0011000010101100110: color_data = Z;
		19'b0011000010101100111: color_data = Z;
		19'b0011000010101101000: color_data = Z;
		19'b0011000010101101001: color_data = Z;
		19'b0011000010101101010: color_data = Z;
		19'b0011000010101101011: color_data = Z;
		19'b0011000010101101100: color_data = Z;
		19'b0011000010101101101: color_data = Z;
		19'b0011000010101101110: color_data = Z;
		19'b0011000010101101111: color_data = Z;
		19'b0011000010101110000: color_data = Z;
		19'b0011000010101110001: color_data = Z;
		19'b0011000010101110010: color_data = Z;
		19'b0011000010101110011: color_data = Z;
		19'b0011000010101110100: color_data = Z;
		19'b0011000010101110101: color_data = Z;
		19'b0011000010101110110: color_data = Z;
		19'b0011000010101110111: color_data = Z;
		19'b0011000010101111000: color_data = Z;
		19'b0011000010101111001: color_data = Z;
		19'b0011000010101111010: color_data = Z;
		19'b0011000010101111011: color_data = Z;
		19'b0011000010101111100: color_data = Z;
		19'b0011000010101111101: color_data = Z;
		19'b0011000010101111110: color_data = Z;
		19'b0011000010101111111: color_data = Z;
		19'b0011000010110000000: color_data = Z;
		19'b0011000010110000001: color_data = Z;
		19'b0011000010110000010: color_data = Z;
		19'b0011000010110000011: color_data = Z;
		19'b0011000010110000100: color_data = Z;
		19'b0011000010110000101: color_data = Z;
		19'b0011000010110000110: color_data = Z;
		19'b0011000010110000111: color_data = Z;
		19'b0011000010110001000: color_data = Z;
		19'b0011000010110001001: color_data = Z;
		19'b0011000010110001010: color_data = Z;
		19'b0011000010110001011: color_data = Z;
		19'b0011000010110001100: color_data = Z;
		19'b0011000010110001101: color_data = Z;
		19'b0011000010110001110: color_data = Z;
		19'b0011000010110001111: color_data = Z;
		19'b0011000010110010000: color_data = Z;
		19'b0011000010110010001: color_data = Z;
		19'b0011000010110010010: color_data = Z;
		19'b0011000010110010011: color_data = Z;
		19'b0011000010110010100: color_data = Z;
		19'b0011000010110010101: color_data = Z;
		19'b0011000010110010110: color_data = Z;
		19'b0011000010110010111: color_data = Z;
		19'b0011000010110011000: color_data = Z;
		19'b0011000010110011001: color_data = Z;
		19'b0011000010110011010: color_data = Z;
		19'b0011000010110011011: color_data = Z;
		19'b0011000010110011100: color_data = Z;
		19'b0011000010110011101: color_data = Z;
		19'b0011000010110011110: color_data = Z;
		19'b0011000010110011111: color_data = Z;
		19'b0011000010110100000: color_data = Z;
		19'b0011000010110100001: color_data = Z;
		19'b0011000010110100010: color_data = Z;
		19'b0011000010110100011: color_data = Z;
		19'b0011000010110100100: color_data = Z;
		19'b0011000010110100101: color_data = Z;
		19'b0011000010110100110: color_data = Z;
		19'b0011000010110100111: color_data = Z;
		19'b0011000010110101000: color_data = Z;
		19'b0011000010110101001: color_data = Z;
		19'b0011000010110101010: color_data = Z;
		19'b0011000010110101011: color_data = Z;
		19'b0011000010110101100: color_data = Z;
		19'b0011000010110101101: color_data = Z;
		19'b0011000010110101110: color_data = Z;
		19'b0011000010110101111: color_data = Z;
		19'b0011000010110110000: color_data = Z;
		19'b0011000010110110001: color_data = Z;
		19'b0011000010110110010: color_data = Z;
		19'b0011000010110110011: color_data = Z;
		19'b0011000010110110100: color_data = Z;
		19'b0011000010110110101: color_data = Z;
		19'b0011000010111000110: color_data = Z;
		19'b0011000010111000111: color_data = Z;
		19'b0011000010111001000: color_data = Z;
		19'b0011000010111001001: color_data = Z;
		19'b0011000010111001010: color_data = Z;
		19'b0011000010111001011: color_data = Z;
		19'b0011000010111001100: color_data = Z;
		19'b0011000010111001101: color_data = Z;
		19'b0011000010111001110: color_data = Z;
		19'b0011000010111001111: color_data = Z;
		19'b0011000100010111000: color_data = Z;
		19'b0011000100010111001: color_data = Z;
		19'b0011000100010111010: color_data = Z;
		19'b0011000100010111011: color_data = Z;
		19'b0011000100010111100: color_data = Z;
		19'b0011000100010111101: color_data = Z;
		19'b0011000100010111110: color_data = Z;
		19'b0011000100010111111: color_data = Z;
		19'b0011000100011000000: color_data = Z;
		19'b0011000100011000001: color_data = Z;
		19'b0011000100011000010: color_data = Z;
		19'b0011000100011000011: color_data = Z;
		19'b0011000100011000100: color_data = Z;
		19'b0011000100011000101: color_data = Z;
		19'b0011000100011000110: color_data = Z;
		19'b0011000100011000111: color_data = Z;
		19'b0011000100011001000: color_data = Z;
		19'b0011000100011001001: color_data = Z;
		19'b0011000100011001010: color_data = Z;
		19'b0011000100011001011: color_data = Z;
		19'b0011000100011001100: color_data = Z;
		19'b0011000100011001101: color_data = Z;
		19'b0011000100011001110: color_data = Z;
		19'b0011000100011001111: color_data = Z;
		19'b0011000100011010000: color_data = Z;
		19'b0011000100011010001: color_data = Z;
		19'b0011000100011010010: color_data = Z;
		19'b0011000100011010011: color_data = Z;
		19'b0011000100011010100: color_data = Z;
		19'b0011000100011010101: color_data = Z;
		19'b0011000100011010110: color_data = Z;
		19'b0011000100011010111: color_data = Z;
		19'b0011000100011011000: color_data = Z;
		19'b0011000100011011001: color_data = Z;
		19'b0011000100011011010: color_data = Z;
		19'b0011000100011011011: color_data = Z;
		19'b0011000100011011100: color_data = Z;
		19'b0011000100011011101: color_data = Z;
		19'b0011000100011011110: color_data = Z;
		19'b0011000100011011111: color_data = Z;
		19'b0011000100011100000: color_data = Z;
		19'b0011000100011100001: color_data = Z;
		19'b0011000100011100010: color_data = Z;
		19'b0011000100011100011: color_data = Z;
		19'b0011000100011100100: color_data = Z;
		19'b0011000100011100101: color_data = Z;
		19'b0011000100011100110: color_data = Z;
		19'b0011000100011100111: color_data = Z;
		19'b0011000100011101000: color_data = Z;
		19'b0011000100011101001: color_data = Z;
		19'b0011000100011101010: color_data = Z;
		19'b0011000100011101011: color_data = Z;
		19'b0011000100011101100: color_data = Z;
		19'b0011000100011101101: color_data = Z;
		19'b0011000100011101110: color_data = Z;
		19'b0011000100011101111: color_data = Z;
		19'b0011000100011110000: color_data = Z;
		19'b0011000100011110001: color_data = Z;
		19'b0011000100011110010: color_data = Z;
		19'b0011000100011110011: color_data = Z;
		19'b0011000100011110100: color_data = Z;
		19'b0011000100011110101: color_data = Z;
		19'b0011000100011110110: color_data = Z;
		19'b0011000100011110111: color_data = Z;
		19'b0011000100011111000: color_data = Z;
		19'b0011000100011111001: color_data = Z;
		19'b0011000100011111010: color_data = Z;
		19'b0011000100011111011: color_data = Z;
		19'b0011000100011111100: color_data = Z;
		19'b0011000100011111101: color_data = Z;
		19'b0011000100011111110: color_data = Z;
		19'b0011000100011111111: color_data = Z;
		19'b0011000100100000000: color_data = Z;
		19'b0011000100100000001: color_data = Z;
		19'b0011000100100000010: color_data = Z;
		19'b0011000100100000011: color_data = Z;
		19'b0011000100100000100: color_data = Z;
		19'b0011000100100000101: color_data = Z;
		19'b0011000100100000110: color_data = Z;
		19'b0011000100100000111: color_data = Z;
		19'b0011000100100001000: color_data = Z;
		19'b0011000100100001001: color_data = Z;
		19'b0011000100100001010: color_data = Z;
		19'b0011000100100001011: color_data = Z;
		19'b0011000100100001100: color_data = Z;
		19'b0011000100100001101: color_data = Z;
		19'b0011000100100001110: color_data = Z;
		19'b0011000100100001111: color_data = Z;
		19'b0011000100100010000: color_data = Z;
		19'b0011000100100010001: color_data = Z;
		19'b0011000100100010010: color_data = Z;
		19'b0011000100100010011: color_data = Z;
		19'b0011000100100010100: color_data = Z;
		19'b0011000100100010101: color_data = Z;
		19'b0011000100100010110: color_data = Z;
		19'b0011000100100010111: color_data = Z;
		19'b0011000100100011000: color_data = Z;
		19'b0011000100100011001: color_data = Z;
		19'b0011000100100011010: color_data = Z;
		19'b0011000100100011011: color_data = Z;
		19'b0011000100100011100: color_data = Z;
		19'b0011000100100011101: color_data = Z;
		19'b0011000100100011110: color_data = Z;
		19'b0011000100100011111: color_data = Z;
		19'b0011000100100100000: color_data = Z;
		19'b0011000100100100001: color_data = Z;
		19'b0011000100100100010: color_data = Z;
		19'b0011000100100100011: color_data = Z;
		19'b0011000100100100100: color_data = Z;
		19'b0011000100100100101: color_data = Z;
		19'b0011000100100100110: color_data = Z;
		19'b0011000100100100111: color_data = Z;
		19'b0011000100100101000: color_data = Z;
		19'b0011000100100101001: color_data = Z;
		19'b0011000100100101010: color_data = Z;
		19'b0011000100100101011: color_data = Z;
		19'b0011000100100101100: color_data = Z;
		19'b0011000100100101101: color_data = Z;
		19'b0011000100100101110: color_data = Z;
		19'b0011000100100101111: color_data = Z;
		19'b0011000100100110000: color_data = Z;
		19'b0011000100100110001: color_data = Z;
		19'b0011000100100110010: color_data = Z;
		19'b0011000100100110011: color_data = Z;
		19'b0011000100100110100: color_data = Z;
		19'b0011000100100110101: color_data = Z;
		19'b0011000100100110110: color_data = Z;
		19'b0011000100100110111: color_data = Z;
		19'b0011000100100111000: color_data = Z;
		19'b0011000100100111001: color_data = Z;
		19'b0011000100100111010: color_data = Z;
		19'b0011000100100111011: color_data = Z;
		19'b0011000100100111100: color_data = Z;
		19'b0011000100100111101: color_data = Z;
		19'b0011000100100111110: color_data = Z;
		19'b0011000100100111111: color_data = Z;
		19'b0011000100101000000: color_data = Z;
		19'b0011000100101000001: color_data = Z;
		19'b0011000100101000010: color_data = Z;
		19'b0011000100101000011: color_data = Z;
		19'b0011000100101000100: color_data = Z;
		19'b0011000100101000101: color_data = Z;
		19'b0011000100101000110: color_data = Z;
		19'b0011000100101000111: color_data = Z;
		19'b0011000100101001000: color_data = Z;
		19'b0011000100101001001: color_data = Z;
		19'b0011000100101001010: color_data = Z;
		19'b0011000100101001011: color_data = Z;
		19'b0011000100101001100: color_data = Z;
		19'b0011000100101001101: color_data = Z;
		19'b0011000100101001110: color_data = Z;
		19'b0011000100101001111: color_data = Z;
		19'b0011000100101010000: color_data = Z;
		19'b0011000100101010001: color_data = Z;
		19'b0011000100101010010: color_data = Z;
		19'b0011000100101010011: color_data = Z;
		19'b0011000100101010100: color_data = Z;
		19'b0011000100101010101: color_data = Z;
		19'b0011000100101010110: color_data = Z;
		19'b0011000100101010111: color_data = Z;
		19'b0011000100101011000: color_data = Z;
		19'b0011000100101011001: color_data = Z;
		19'b0011000100101011010: color_data = Z;
		19'b0011000100101011011: color_data = Z;
		19'b0011000100101011100: color_data = Z;
		19'b0011000100101011101: color_data = Z;
		19'b0011000100101011110: color_data = Z;
		19'b0011000100101011111: color_data = Z;
		19'b0011000100101100000: color_data = Z;
		19'b0011000100101100001: color_data = Z;
		19'b0011000100101100010: color_data = Z;
		19'b0011000100101100011: color_data = Z;
		19'b0011000100101100100: color_data = Z;
		19'b0011000100101100101: color_data = Z;
		19'b0011000100101100110: color_data = Z;
		19'b0011000100101100111: color_data = Z;
		19'b0011000100101101000: color_data = Z;
		19'b0011000100101101001: color_data = Z;
		19'b0011000100101101010: color_data = Z;
		19'b0011000100101101011: color_data = Z;
		19'b0011000100101101100: color_data = Z;
		19'b0011000100101101101: color_data = Z;
		19'b0011000100101101110: color_data = Z;
		19'b0011000100101101111: color_data = Z;
		19'b0011000100101110000: color_data = Z;
		19'b0011000100101110001: color_data = Z;
		19'b0011000100101110010: color_data = Z;
		19'b0011000100101110011: color_data = Z;
		19'b0011000100101110100: color_data = Z;
		19'b0011000100101110101: color_data = Z;
		19'b0011000100101110110: color_data = Z;
		19'b0011000100101110111: color_data = Z;
		19'b0011000100101111000: color_data = Z;
		19'b0011000100101111001: color_data = Z;
		19'b0011000100101111010: color_data = Z;
		19'b0011000100101111011: color_data = Z;
		19'b0011000100101111100: color_data = Z;
		19'b0011000100101111101: color_data = Z;
		19'b0011000100101111110: color_data = Z;
		19'b0011000100101111111: color_data = Z;
		19'b0011000100110000000: color_data = Z;
		19'b0011000100110000001: color_data = Z;
		19'b0011000100110000010: color_data = Z;
		19'b0011000100110000011: color_data = Z;
		19'b0011000100110000100: color_data = Z;
		19'b0011000100110000101: color_data = Z;
		19'b0011000100110000110: color_data = Z;
		19'b0011000100110000111: color_data = Z;
		19'b0011000100110001000: color_data = Z;
		19'b0011000100110001001: color_data = Z;
		19'b0011000100110001010: color_data = Z;
		19'b0011000100110001011: color_data = Z;
		19'b0011000100110001100: color_data = Z;
		19'b0011000100110001101: color_data = Z;
		19'b0011000100110001110: color_data = Z;
		19'b0011000100110001111: color_data = Z;
		19'b0011000100110010000: color_data = Z;
		19'b0011000100110010001: color_data = Z;
		19'b0011000100110010010: color_data = Z;
		19'b0011000100110010011: color_data = Z;
		19'b0011000100110010100: color_data = Z;
		19'b0011000100110010101: color_data = Z;
		19'b0011000100110010110: color_data = Z;
		19'b0011000100110010111: color_data = Z;
		19'b0011000100110011000: color_data = Z;
		19'b0011000100110011001: color_data = Z;
		19'b0011000100110011010: color_data = Z;
		19'b0011000100110011011: color_data = Z;
		19'b0011000100110011100: color_data = Z;
		19'b0011000100110011101: color_data = Z;
		19'b0011000100110011110: color_data = Z;
		19'b0011000100110011111: color_data = Z;
		19'b0011000100110100000: color_data = Z;
		19'b0011000100110100001: color_data = Z;
		19'b0011000100110100010: color_data = Z;
		19'b0011000100110100011: color_data = Z;
		19'b0011000100110100100: color_data = Z;
		19'b0011000100110100101: color_data = Z;
		19'b0011000100110100110: color_data = Z;
		19'b0011000100110100111: color_data = Z;
		19'b0011000100110101000: color_data = Z;
		19'b0011000100110101001: color_data = Z;
		19'b0011000100110101010: color_data = Z;
		19'b0011000100110101011: color_data = Z;
		19'b0011000100110101100: color_data = Z;
		19'b0011000100110101101: color_data = Z;
		19'b0011000100110101110: color_data = Z;
		19'b0011000100110101111: color_data = Z;
		19'b0011000100110110000: color_data = Z;
		19'b0011000100110110001: color_data = Z;
		19'b0011000100110110010: color_data = Z;
		19'b0011000100110110011: color_data = Z;
		19'b0011000100110110100: color_data = Z;
		19'b0011000100110110101: color_data = Z;
		19'b0011000100111000111: color_data = Z;
		19'b0011000100111001000: color_data = Z;
		19'b0011000100111001001: color_data = Z;
		19'b0011000100111001010: color_data = Z;
		19'b0011000100111001011: color_data = Z;
		19'b0011000100111001100: color_data = Z;
		19'b0011000100111001101: color_data = Z;
		19'b0011000110010110110: color_data = Z;
		19'b0011000110010110111: color_data = Z;
		19'b0011000110010111000: color_data = Z;
		19'b0011000110010111001: color_data = Z;
		19'b0011000110010111010: color_data = Z;
		19'b0011000110010111011: color_data = Z;
		19'b0011000110010111100: color_data = Z;
		19'b0011000110010111101: color_data = Z;
		19'b0011000110010111110: color_data = Z;
		19'b0011000110010111111: color_data = Z;
		19'b0011000110011000000: color_data = Z;
		19'b0011000110011000001: color_data = Z;
		19'b0011000110011000010: color_data = Z;
		19'b0011000110011000011: color_data = Z;
		19'b0011000110011000100: color_data = Z;
		19'b0011000110011000101: color_data = Z;
		19'b0011000110011000110: color_data = Z;
		19'b0011000110011000111: color_data = Z;
		19'b0011000110011001000: color_data = Z;
		19'b0011000110011001001: color_data = Z;
		19'b0011000110011001010: color_data = Z;
		19'b0011000110011001011: color_data = Z;
		19'b0011000110011001100: color_data = Z;
		19'b0011000110011001101: color_data = Z;
		19'b0011000110011001110: color_data = Z;
		19'b0011000110011001111: color_data = Z;
		19'b0011000110011010000: color_data = Z;
		19'b0011000110011010001: color_data = Z;
		19'b0011000110011010010: color_data = Z;
		19'b0011000110011010011: color_data = Z;
		19'b0011000110011010100: color_data = Z;
		19'b0011000110011010101: color_data = Z;
		19'b0011000110011010110: color_data = Z;
		19'b0011000110011010111: color_data = Z;
		19'b0011000110011011000: color_data = Z;
		19'b0011000110011011001: color_data = Z;
		19'b0011000110011011010: color_data = Z;
		19'b0011000110011011011: color_data = Z;
		19'b0011000110011011100: color_data = Z;
		19'b0011000110011011101: color_data = Z;
		19'b0011000110011011110: color_data = Z;
		19'b0011000110011011111: color_data = Z;
		19'b0011000110011100000: color_data = Z;
		19'b0011000110011100001: color_data = Z;
		19'b0011000110011100010: color_data = Z;
		19'b0011000110011100011: color_data = Z;
		19'b0011000110011100100: color_data = Z;
		19'b0011000110011100101: color_data = Z;
		19'b0011000110011100110: color_data = Z;
		19'b0011000110011100111: color_data = Z;
		19'b0011000110011101000: color_data = Z;
		19'b0011000110011101001: color_data = Z;
		19'b0011000110011101010: color_data = Z;
		19'b0011000110011101011: color_data = Z;
		19'b0011000110011101100: color_data = Z;
		19'b0011000110011101101: color_data = Z;
		19'b0011000110011101110: color_data = Z;
		19'b0011000110011101111: color_data = Z;
		19'b0011000110011110000: color_data = Z;
		19'b0011000110011110001: color_data = Z;
		19'b0011000110011110010: color_data = Z;
		19'b0011000110011110011: color_data = Z;
		19'b0011000110011110100: color_data = Z;
		19'b0011000110011110101: color_data = Z;
		19'b0011000110011110110: color_data = Z;
		19'b0011000110011110111: color_data = Z;
		19'b0011000110011111000: color_data = Z;
		19'b0011000110011111001: color_data = Z;
		19'b0011000110011111010: color_data = Z;
		19'b0011000110011111011: color_data = Z;
		19'b0011000110011111100: color_data = Z;
		19'b0011000110011111101: color_data = Z;
		19'b0011000110011111110: color_data = Z;
		19'b0011000110011111111: color_data = Z;
		19'b0011000110100000000: color_data = Z;
		19'b0011000110100000001: color_data = Z;
		19'b0011000110100000010: color_data = Z;
		19'b0011000110100000011: color_data = Z;
		19'b0011000110100000100: color_data = Z;
		19'b0011000110100000101: color_data = Z;
		19'b0011000110100000110: color_data = Z;
		19'b0011000110100000111: color_data = Z;
		19'b0011000110100001000: color_data = Z;
		19'b0011000110100001001: color_data = Z;
		19'b0011000110100001010: color_data = Z;
		19'b0011000110100001011: color_data = Z;
		19'b0011000110100001100: color_data = Z;
		19'b0011000110100001101: color_data = Z;
		19'b0011000110100001110: color_data = Z;
		19'b0011000110100001111: color_data = Z;
		19'b0011000110100010000: color_data = Z;
		19'b0011000110100010001: color_data = Z;
		19'b0011000110100010010: color_data = Z;
		19'b0011000110100010011: color_data = Z;
		19'b0011000110100010100: color_data = Z;
		19'b0011000110100010101: color_data = Z;
		19'b0011000110100010110: color_data = Z;
		19'b0011000110100010111: color_data = Z;
		19'b0011000110100011000: color_data = Z;
		19'b0011000110100011001: color_data = Z;
		19'b0011000110100011010: color_data = Z;
		19'b0011000110100011011: color_data = Z;
		19'b0011000110100011100: color_data = Z;
		19'b0011000110100011101: color_data = Z;
		19'b0011000110100011110: color_data = Z;
		19'b0011000110100011111: color_data = Z;
		19'b0011000110100100000: color_data = Z;
		19'b0011000110100100001: color_data = Z;
		19'b0011000110100100010: color_data = Z;
		19'b0011000110100100011: color_data = Z;
		19'b0011000110100100100: color_data = Z;
		19'b0011000110100100101: color_data = Z;
		19'b0011000110100100110: color_data = Z;
		19'b0011000110100100111: color_data = Z;
		19'b0011000110100101000: color_data = Z;
		19'b0011000110100101001: color_data = Z;
		19'b0011000110100101010: color_data = Z;
		19'b0011000110100101011: color_data = Z;
		19'b0011000110100101100: color_data = Z;
		19'b0011000110100101101: color_data = Z;
		19'b0011000110100101110: color_data = Z;
		19'b0011000110100101111: color_data = Z;
		19'b0011000110100110000: color_data = Z;
		19'b0011000110100110001: color_data = Z;
		19'b0011000110100110010: color_data = Z;
		19'b0011000110100110011: color_data = Z;
		19'b0011000110100110100: color_data = Z;
		19'b0011000110100110101: color_data = Z;
		19'b0011000110100110110: color_data = Z;
		19'b0011000110100110111: color_data = Z;
		19'b0011000110100111000: color_data = Z;
		19'b0011000110100111001: color_data = Z;
		19'b0011000110100111010: color_data = Z;
		19'b0011000110100111011: color_data = Z;
		19'b0011000110100111100: color_data = Z;
		19'b0011000110100111101: color_data = Z;
		19'b0011000110100111110: color_data = Z;
		19'b0011000110100111111: color_data = Z;
		19'b0011000110101000000: color_data = Z;
		19'b0011000110101000001: color_data = Z;
		19'b0011000110101000010: color_data = Z;
		19'b0011000110101000011: color_data = Z;
		19'b0011000110101000100: color_data = Z;
		19'b0011000110101000101: color_data = Z;
		19'b0011000110101000110: color_data = Z;
		19'b0011000110101000111: color_data = Z;
		19'b0011000110101001000: color_data = Z;
		19'b0011000110101001001: color_data = Z;
		19'b0011000110101001010: color_data = Z;
		19'b0011000110101001011: color_data = Z;
		19'b0011000110101001100: color_data = Z;
		19'b0011000110101001101: color_data = Z;
		19'b0011000110101001110: color_data = Z;
		19'b0011000110101001111: color_data = Z;
		19'b0011000110101010000: color_data = Z;
		19'b0011000110101010001: color_data = Z;
		19'b0011000110101010010: color_data = Z;
		19'b0011000110101010011: color_data = Z;
		19'b0011000110101010100: color_data = Z;
		19'b0011000110101010101: color_data = Z;
		19'b0011000110101010110: color_data = Z;
		19'b0011000110101010111: color_data = Z;
		19'b0011000110101011000: color_data = Z;
		19'b0011000110101011001: color_data = Z;
		19'b0011000110101011010: color_data = Z;
		19'b0011000110101011011: color_data = Z;
		19'b0011000110101011100: color_data = Z;
		19'b0011000110101011101: color_data = Z;
		19'b0011000110101011110: color_data = Z;
		19'b0011000110101011111: color_data = Z;
		19'b0011000110101100000: color_data = Z;
		19'b0011000110101100001: color_data = Z;
		19'b0011000110101100010: color_data = Z;
		19'b0011000110101100011: color_data = Z;
		19'b0011000110101100100: color_data = Z;
		19'b0011000110101100101: color_data = Z;
		19'b0011000110101100110: color_data = Z;
		19'b0011000110101100111: color_data = Z;
		19'b0011000110101101000: color_data = Z;
		19'b0011000110101101001: color_data = Z;
		19'b0011000110101101010: color_data = Z;
		19'b0011000110101101011: color_data = Z;
		19'b0011000110101101100: color_data = Z;
		19'b0011000110101101101: color_data = Z;
		19'b0011000110101101110: color_data = Z;
		19'b0011000110101101111: color_data = Z;
		19'b0011000110101110000: color_data = Z;
		19'b0011000110101110001: color_data = Z;
		19'b0011000110101110010: color_data = Z;
		19'b0011000110101110011: color_data = Z;
		19'b0011000110101110100: color_data = Z;
		19'b0011000110101110101: color_data = Z;
		19'b0011000110101110110: color_data = Z;
		19'b0011000110101110111: color_data = Z;
		19'b0011000110101111000: color_data = Z;
		19'b0011000110101111001: color_data = Z;
		19'b0011000110101111010: color_data = Z;
		19'b0011000110101111011: color_data = Z;
		19'b0011000110101111100: color_data = Z;
		19'b0011000110101111101: color_data = Z;
		19'b0011000110101111110: color_data = Z;
		19'b0011000110101111111: color_data = Z;
		19'b0011000110110000000: color_data = Z;
		19'b0011000110110000001: color_data = Z;
		19'b0011000110110000010: color_data = Z;
		19'b0011000110110000011: color_data = Z;
		19'b0011000110110000100: color_data = Z;
		19'b0011000110110000101: color_data = Z;
		19'b0011000110110000110: color_data = Z;
		19'b0011000110110000111: color_data = Z;
		19'b0011000110110001000: color_data = Z;
		19'b0011000110110001001: color_data = Z;
		19'b0011000110110001010: color_data = Z;
		19'b0011000110110001011: color_data = Z;
		19'b0011000110110001100: color_data = Z;
		19'b0011000110110001101: color_data = Z;
		19'b0011000110110001110: color_data = Z;
		19'b0011000110110001111: color_data = Z;
		19'b0011000110110010000: color_data = Z;
		19'b0011000110110010001: color_data = Z;
		19'b0011000110110010010: color_data = Z;
		19'b0011000110110010011: color_data = Z;
		19'b0011000110110010100: color_data = Z;
		19'b0011000110110010101: color_data = Z;
		19'b0011000110110010110: color_data = Z;
		19'b0011000110110010111: color_data = Z;
		19'b0011000110110011000: color_data = Z;
		19'b0011000110110011001: color_data = Z;
		19'b0011000110110011010: color_data = Z;
		19'b0011000110110011011: color_data = Z;
		19'b0011000110110011100: color_data = Z;
		19'b0011000110110011101: color_data = Z;
		19'b0011000110110011110: color_data = Z;
		19'b0011000110110011111: color_data = Z;
		19'b0011000110110100000: color_data = Z;
		19'b0011000110110100001: color_data = Z;
		19'b0011000110110100010: color_data = Z;
		19'b0011000110110100011: color_data = Z;
		19'b0011000110110100100: color_data = Z;
		19'b0011000110110100101: color_data = Z;
		19'b0011000110110100110: color_data = Z;
		19'b0011000110110100111: color_data = Z;
		19'b0011000110110101000: color_data = Z;
		19'b0011000110110101001: color_data = Z;
		19'b0011000110110101010: color_data = Z;
		19'b0011000110110101011: color_data = Z;
		19'b0011000110110101100: color_data = Z;
		19'b0011000110110101101: color_data = Z;
		19'b0011000110110101110: color_data = Z;
		19'b0011000110110101111: color_data = Z;
		19'b0011000110110110000: color_data = Z;
		19'b0011000110110110001: color_data = Z;
		19'b0011000110110110010: color_data = Z;
		19'b0011000110110110011: color_data = Z;
		19'b0011000110110110100: color_data = Z;
		19'b0011000110110110101: color_data = Z;
		19'b0011000110111001000: color_data = Z;
		19'b0011000110111001001: color_data = Z;
		19'b0011000110111001010: color_data = Z;
		19'b0011000110111001011: color_data = Z;
		19'b0011000110111001100: color_data = Z;
		19'b0011001000010110101: color_data = Z;
		19'b0011001000010110110: color_data = Z;
		19'b0011001000010110111: color_data = Z;
		19'b0011001000010111000: color_data = Z;
		19'b0011001000010111001: color_data = Z;
		19'b0011001000010111010: color_data = Z;
		19'b0011001000010111011: color_data = Z;
		19'b0011001000010111100: color_data = Z;
		19'b0011001000010111101: color_data = Z;
		19'b0011001000010111110: color_data = Z;
		19'b0011001000010111111: color_data = Z;
		19'b0011001000011000000: color_data = Z;
		19'b0011001000011000001: color_data = Z;
		19'b0011001000011000010: color_data = Z;
		19'b0011001000011000011: color_data = Z;
		19'b0011001000011000100: color_data = Z;
		19'b0011001000011000101: color_data = Z;
		19'b0011001000011000110: color_data = Z;
		19'b0011001000011000111: color_data = Z;
		19'b0011001000011001000: color_data = Z;
		19'b0011001000011001001: color_data = Z;
		19'b0011001000011001010: color_data = Z;
		19'b0011001000011001011: color_data = Z;
		19'b0011001000011001100: color_data = Z;
		19'b0011001000011001101: color_data = Z;
		19'b0011001000011001110: color_data = Z;
		19'b0011001000011001111: color_data = Z;
		19'b0011001000011010000: color_data = Z;
		19'b0011001000011010001: color_data = Z;
		19'b0011001000011010010: color_data = Z;
		19'b0011001000011010011: color_data = Z;
		19'b0011001000011010100: color_data = Z;
		19'b0011001000011010101: color_data = Z;
		19'b0011001000011010110: color_data = Z;
		19'b0011001000011010111: color_data = Z;
		19'b0011001000011011000: color_data = Z;
		19'b0011001000011011001: color_data = Z;
		19'b0011001000011011010: color_data = Z;
		19'b0011001000011011011: color_data = Z;
		19'b0011001000011011100: color_data = Z;
		19'b0011001000011011101: color_data = Z;
		19'b0011001000011011110: color_data = Z;
		19'b0011001000011011111: color_data = Z;
		19'b0011001000011100000: color_data = Z;
		19'b0011001000011100001: color_data = Z;
		19'b0011001000011100010: color_data = Z;
		19'b0011001000011100011: color_data = Z;
		19'b0011001000011100100: color_data = Z;
		19'b0011001000011100101: color_data = Z;
		19'b0011001000011100110: color_data = Z;
		19'b0011001000011100111: color_data = Z;
		19'b0011001000011101000: color_data = Z;
		19'b0011001000011101001: color_data = Z;
		19'b0011001000011101010: color_data = Z;
		19'b0011001000011101011: color_data = Z;
		19'b0011001000011101100: color_data = Z;
		19'b0011001000011101101: color_data = Z;
		19'b0011001000011101110: color_data = Z;
		19'b0011001000011101111: color_data = Z;
		19'b0011001000011110000: color_data = Z;
		19'b0011001000011110001: color_data = Z;
		19'b0011001000011110010: color_data = Z;
		19'b0011001000011110011: color_data = Z;
		19'b0011001000011110100: color_data = Z;
		19'b0011001000011110101: color_data = Z;
		19'b0011001000011110110: color_data = Z;
		19'b0011001000011110111: color_data = Z;
		19'b0011001000011111000: color_data = Z;
		19'b0011001000011111001: color_data = Z;
		19'b0011001000011111010: color_data = Z;
		19'b0011001000011111011: color_data = Z;
		19'b0011001000011111100: color_data = Z;
		19'b0011001000011111101: color_data = Z;
		19'b0011001000011111110: color_data = Z;
		19'b0011001000011111111: color_data = Z;
		19'b0011001000100000000: color_data = Z;
		19'b0011001000100000001: color_data = Z;
		19'b0011001000100000010: color_data = Z;
		19'b0011001000100000011: color_data = Z;
		19'b0011001000100000100: color_data = Z;
		19'b0011001000100000101: color_data = Z;
		19'b0011001000100000110: color_data = Z;
		19'b0011001000100000111: color_data = Z;
		19'b0011001000100001000: color_data = Z;
		19'b0011001000100001001: color_data = Z;
		19'b0011001000100001010: color_data = Z;
		19'b0011001000100001011: color_data = Z;
		19'b0011001000100001100: color_data = Z;
		19'b0011001000100001101: color_data = Z;
		19'b0011001000100001110: color_data = Z;
		19'b0011001000100001111: color_data = Z;
		19'b0011001000100010000: color_data = Z;
		19'b0011001000100010001: color_data = Z;
		19'b0011001000100010010: color_data = Z;
		19'b0011001000100010011: color_data = Z;
		19'b0011001000100010100: color_data = Z;
		19'b0011001000100010101: color_data = Z;
		19'b0011001000100010110: color_data = Z;
		19'b0011001000100010111: color_data = Z;
		19'b0011001000100011000: color_data = Z;
		19'b0011001000100011001: color_data = Z;
		19'b0011001000100011010: color_data = Z;
		19'b0011001000100011011: color_data = Z;
		19'b0011001000100011100: color_data = Z;
		19'b0011001000100011101: color_data = Z;
		19'b0011001000100011110: color_data = Z;
		19'b0011001000100011111: color_data = Z;
		19'b0011001000100100000: color_data = Z;
		19'b0011001000100100001: color_data = Z;
		19'b0011001000100100010: color_data = Z;
		19'b0011001000100100011: color_data = Z;
		19'b0011001000100100100: color_data = Z;
		19'b0011001000100100101: color_data = Z;
		19'b0011001000100100110: color_data = Z;
		19'b0011001000100100111: color_data = Z;
		19'b0011001000100101000: color_data = Z;
		19'b0011001000100101001: color_data = Z;
		19'b0011001000100101010: color_data = Z;
		19'b0011001000100101011: color_data = Z;
		19'b0011001000100101100: color_data = Z;
		19'b0011001000100101101: color_data = Z;
		19'b0011001000100101110: color_data = Z;
		19'b0011001000100101111: color_data = Z;
		19'b0011001000100110000: color_data = Z;
		19'b0011001000100110001: color_data = Z;
		19'b0011001000100110010: color_data = Z;
		19'b0011001000100110011: color_data = Z;
		19'b0011001000100110100: color_data = Z;
		19'b0011001000100110101: color_data = Z;
		19'b0011001000100110110: color_data = Z;
		19'b0011001000100110111: color_data = Z;
		19'b0011001000100111000: color_data = Z;
		19'b0011001000100111001: color_data = Z;
		19'b0011001000100111010: color_data = Z;
		19'b0011001000100111011: color_data = Z;
		19'b0011001000100111100: color_data = Z;
		19'b0011001000100111101: color_data = Z;
		19'b0011001000100111110: color_data = Z;
		19'b0011001000100111111: color_data = Z;
		19'b0011001000101000000: color_data = Z;
		19'b0011001000101000001: color_data = Z;
		19'b0011001000101000010: color_data = Z;
		19'b0011001000101000011: color_data = Z;
		19'b0011001000101000100: color_data = Z;
		19'b0011001000101000101: color_data = Z;
		19'b0011001000101000110: color_data = Z;
		19'b0011001000101000111: color_data = Z;
		19'b0011001000101001000: color_data = Z;
		19'b0011001000101001001: color_data = Z;
		19'b0011001000101001010: color_data = Z;
		19'b0011001000101001011: color_data = Z;
		19'b0011001000101001100: color_data = Z;
		19'b0011001000101001101: color_data = Z;
		19'b0011001000101001110: color_data = Z;
		19'b0011001000101001111: color_data = Z;
		19'b0011001000101010000: color_data = Z;
		19'b0011001000101010001: color_data = Z;
		19'b0011001000101010010: color_data = Z;
		19'b0011001000101010011: color_data = Z;
		19'b0011001000101010100: color_data = Z;
		19'b0011001000101010101: color_data = Z;
		19'b0011001000101010110: color_data = Z;
		19'b0011001000101010111: color_data = Z;
		19'b0011001000101011000: color_data = Z;
		19'b0011001000101011001: color_data = Z;
		19'b0011001000101011010: color_data = Z;
		19'b0011001000101011011: color_data = Z;
		19'b0011001000101011100: color_data = Z;
		19'b0011001000101011101: color_data = Z;
		19'b0011001000101011110: color_data = Z;
		19'b0011001000101011111: color_data = Z;
		19'b0011001000101100000: color_data = Z;
		19'b0011001000101100001: color_data = Z;
		19'b0011001000101100010: color_data = Z;
		19'b0011001000101100011: color_data = Z;
		19'b0011001000101100100: color_data = Z;
		19'b0011001000101100101: color_data = Z;
		19'b0011001000101100110: color_data = Z;
		19'b0011001000101100111: color_data = Z;
		19'b0011001000101101000: color_data = Z;
		19'b0011001000101101001: color_data = Z;
		19'b0011001000101101010: color_data = Z;
		19'b0011001000101101011: color_data = Z;
		19'b0011001000101101100: color_data = Z;
		19'b0011001000101101101: color_data = Z;
		19'b0011001000101101110: color_data = Z;
		19'b0011001000101101111: color_data = Z;
		19'b0011001000101110000: color_data = Z;
		19'b0011001000101110001: color_data = Z;
		19'b0011001000101110010: color_data = Z;
		19'b0011001000101110011: color_data = Z;
		19'b0011001000101110100: color_data = Z;
		19'b0011001000101110101: color_data = Z;
		19'b0011001000101110110: color_data = Z;
		19'b0011001000101110111: color_data = Z;
		19'b0011001000101111000: color_data = Z;
		19'b0011001000101111001: color_data = Z;
		19'b0011001000101111010: color_data = Z;
		19'b0011001000101111011: color_data = Z;
		19'b0011001000101111100: color_data = Z;
		19'b0011001000101111101: color_data = Z;
		19'b0011001000101111110: color_data = Z;
		19'b0011001000101111111: color_data = Z;
		19'b0011001000110000000: color_data = Z;
		19'b0011001000110000001: color_data = Z;
		19'b0011001000110000010: color_data = Z;
		19'b0011001000110000011: color_data = Z;
		19'b0011001000110000100: color_data = Z;
		19'b0011001000110000101: color_data = Z;
		19'b0011001000110000110: color_data = Z;
		19'b0011001000110000111: color_data = Z;
		19'b0011001000110001000: color_data = Z;
		19'b0011001000110001001: color_data = Z;
		19'b0011001000110001010: color_data = Z;
		19'b0011001000110001011: color_data = Z;
		19'b0011001000110001100: color_data = Z;
		19'b0011001000110001101: color_data = Z;
		19'b0011001000110001110: color_data = Z;
		19'b0011001000110001111: color_data = Z;
		19'b0011001000110010000: color_data = Z;
		19'b0011001000110010001: color_data = Z;
		19'b0011001000110010010: color_data = Z;
		19'b0011001000110010011: color_data = Z;
		19'b0011001000110010100: color_data = Z;
		19'b0011001000110010101: color_data = Z;
		19'b0011001000110010110: color_data = Z;
		19'b0011001000110010111: color_data = Z;
		19'b0011001000110011000: color_data = Z;
		19'b0011001000110011001: color_data = Z;
		19'b0011001000110011010: color_data = Z;
		19'b0011001000110011011: color_data = Z;
		19'b0011001000110011100: color_data = Z;
		19'b0011001000110011101: color_data = Z;
		19'b0011001000110011110: color_data = Z;
		19'b0011001000110011111: color_data = Z;
		19'b0011001000110100000: color_data = Z;
		19'b0011001000110100001: color_data = Z;
		19'b0011001000110100010: color_data = Z;
		19'b0011001000110100011: color_data = Z;
		19'b0011001000110100100: color_data = Z;
		19'b0011001000110100101: color_data = Z;
		19'b0011001000110100110: color_data = Z;
		19'b0011001000110100111: color_data = Z;
		19'b0011001000110101000: color_data = Z;
		19'b0011001000110101001: color_data = Z;
		19'b0011001000110101010: color_data = Z;
		19'b0011001000110101011: color_data = Z;
		19'b0011001000110101100: color_data = Z;
		19'b0011001000110101101: color_data = Z;
		19'b0011001000110101110: color_data = Z;
		19'b0011001000110101111: color_data = Z;
		19'b0011001000110110000: color_data = Z;
		19'b0011001000110110001: color_data = Z;
		19'b0011001000110110010: color_data = Z;
		19'b0011001000110110011: color_data = Z;
		19'b0011001000110110100: color_data = Z;
		19'b0011001000110110101: color_data = Z;
		19'b0011001000111001010: color_data = Z;
		19'b0011001000111001111: color_data = Z;
		19'b0011001010010110100: color_data = Z;
		19'b0011001010010110101: color_data = Z;
		19'b0011001010010110110: color_data = Z;
		19'b0011001010010110111: color_data = Z;
		19'b0011001010010111000: color_data = Z;
		19'b0011001010010111001: color_data = Z;
		19'b0011001010010111010: color_data = Z;
		19'b0011001010010111011: color_data = Z;
		19'b0011001010010111100: color_data = Z;
		19'b0011001010010111101: color_data = Z;
		19'b0011001010010111110: color_data = Z;
		19'b0011001010010111111: color_data = Z;
		19'b0011001010011000000: color_data = Z;
		19'b0011001010011000001: color_data = Z;
		19'b0011001010011000010: color_data = Z;
		19'b0011001010011000011: color_data = Z;
		19'b0011001010011000100: color_data = Z;
		19'b0011001010011000101: color_data = Z;
		19'b0011001010011000110: color_data = Z;
		19'b0011001010011000111: color_data = Z;
		19'b0011001010011001000: color_data = Z;
		19'b0011001010011001001: color_data = Z;
		19'b0011001010011001010: color_data = Z;
		19'b0011001010011001011: color_data = Z;
		19'b0011001010011001100: color_data = Z;
		19'b0011001010011001101: color_data = Z;
		19'b0011001010011001110: color_data = Z;
		19'b0011001010011001111: color_data = Z;
		19'b0011001010011010000: color_data = Z;
		19'b0011001010011010001: color_data = Z;
		19'b0011001010011010010: color_data = Z;
		19'b0011001010011010011: color_data = Z;
		19'b0011001010011010100: color_data = Z;
		19'b0011001010011010101: color_data = Z;
		19'b0011001010011010110: color_data = Z;
		19'b0011001010011010111: color_data = Z;
		19'b0011001010011011000: color_data = Z;
		19'b0011001010011011001: color_data = Z;
		19'b0011001010011011010: color_data = Z;
		19'b0011001010011011011: color_data = Z;
		19'b0011001010011011100: color_data = Z;
		19'b0011001010011011101: color_data = Z;
		19'b0011001010011011110: color_data = Z;
		19'b0011001010011011111: color_data = Z;
		19'b0011001010011100000: color_data = Z;
		19'b0011001010011100001: color_data = Z;
		19'b0011001010011100010: color_data = Z;
		19'b0011001010011100011: color_data = Z;
		19'b0011001010011100100: color_data = Z;
		19'b0011001010011100101: color_data = Z;
		19'b0011001010011100110: color_data = Z;
		19'b0011001010011100111: color_data = Z;
		19'b0011001010011101000: color_data = Z;
		19'b0011001010011101001: color_data = Z;
		19'b0011001010011101010: color_data = Z;
		19'b0011001010011101011: color_data = Z;
		19'b0011001010011101100: color_data = Z;
		19'b0011001010011101101: color_data = Z;
		19'b0011001010011101110: color_data = Z;
		19'b0011001010011101111: color_data = Z;
		19'b0011001010011110000: color_data = Z;
		19'b0011001010011110001: color_data = Z;
		19'b0011001010011110010: color_data = Z;
		19'b0011001010011110011: color_data = Z;
		19'b0011001010011110100: color_data = Z;
		19'b0011001010011110101: color_data = Z;
		19'b0011001010011110110: color_data = Z;
		19'b0011001010011110111: color_data = Z;
		19'b0011001010011111000: color_data = Z;
		19'b0011001010011111001: color_data = Z;
		19'b0011001010011111010: color_data = Z;
		19'b0011001010011111011: color_data = Z;
		19'b0011001010011111100: color_data = Z;
		19'b0011001010011111101: color_data = Z;
		19'b0011001010011111110: color_data = Z;
		19'b0011001010011111111: color_data = Z;
		19'b0011001010100000000: color_data = Z;
		19'b0011001010100000001: color_data = Z;
		19'b0011001010100000010: color_data = Z;
		19'b0011001010100000011: color_data = Z;
		19'b0011001010100000100: color_data = Z;
		19'b0011001010100000101: color_data = Z;
		19'b0011001010100000110: color_data = Z;
		19'b0011001010100000111: color_data = Z;
		19'b0011001010100001000: color_data = Z;
		19'b0011001010100001001: color_data = Z;
		19'b0011001010100001010: color_data = Z;
		19'b0011001010100001011: color_data = Z;
		19'b0011001010100001100: color_data = Z;
		19'b0011001010100001101: color_data = Z;
		19'b0011001010100001110: color_data = Z;
		19'b0011001010100001111: color_data = Z;
		19'b0011001010100010000: color_data = Z;
		19'b0011001010100010001: color_data = Z;
		19'b0011001010100010010: color_data = Z;
		19'b0011001010100010011: color_data = Z;
		19'b0011001010100010100: color_data = Z;
		19'b0011001010100010101: color_data = Z;
		19'b0011001010100010110: color_data = Z;
		19'b0011001010100010111: color_data = Z;
		19'b0011001010100011000: color_data = Z;
		19'b0011001010100011001: color_data = Z;
		19'b0011001010100011010: color_data = Z;
		19'b0011001010100011011: color_data = Z;
		19'b0011001010100011100: color_data = Z;
		19'b0011001010100011101: color_data = Z;
		19'b0011001010100011110: color_data = Z;
		19'b0011001010100011111: color_data = Z;
		19'b0011001010100100000: color_data = Z;
		19'b0011001010100100001: color_data = Z;
		19'b0011001010100100010: color_data = Z;
		19'b0011001010100100011: color_data = Z;
		19'b0011001010100100100: color_data = Z;
		19'b0011001010100100101: color_data = Z;
		19'b0011001010100100110: color_data = Z;
		19'b0011001010100100111: color_data = Z;
		19'b0011001010100101000: color_data = Z;
		19'b0011001010100101001: color_data = Z;
		19'b0011001010100101010: color_data = Z;
		19'b0011001010100101011: color_data = Z;
		19'b0011001010100101100: color_data = Z;
		19'b0011001010100101101: color_data = Z;
		19'b0011001010100101110: color_data = Z;
		19'b0011001010100101111: color_data = Z;
		19'b0011001010100110000: color_data = Z;
		19'b0011001010100110001: color_data = Z;
		19'b0011001010100110010: color_data = Z;
		19'b0011001010100110011: color_data = Z;
		19'b0011001010100110100: color_data = Z;
		19'b0011001010100110101: color_data = Z;
		19'b0011001010100110110: color_data = Z;
		19'b0011001010100110111: color_data = Z;
		19'b0011001010100111000: color_data = Z;
		19'b0011001010100111001: color_data = Z;
		19'b0011001010100111010: color_data = Z;
		19'b0011001010100111011: color_data = Z;
		19'b0011001010100111100: color_data = Z;
		19'b0011001010100111101: color_data = Z;
		19'b0011001010100111110: color_data = Z;
		19'b0011001010100111111: color_data = Z;
		19'b0011001010101000000: color_data = Z;
		19'b0011001010101000001: color_data = Z;
		19'b0011001010101000010: color_data = Z;
		19'b0011001010101000011: color_data = Z;
		19'b0011001010101000100: color_data = Z;
		19'b0011001010101000101: color_data = Z;
		19'b0011001010101000110: color_data = Z;
		19'b0011001010101000111: color_data = Z;
		19'b0011001010101001000: color_data = Z;
		19'b0011001010101001001: color_data = Z;
		19'b0011001010101001010: color_data = Z;
		19'b0011001010101001011: color_data = Z;
		19'b0011001010101001100: color_data = Z;
		19'b0011001010101001101: color_data = Z;
		19'b0011001010101001110: color_data = Z;
		19'b0011001010101001111: color_data = Z;
		19'b0011001010101010000: color_data = Z;
		19'b0011001010101010001: color_data = Z;
		19'b0011001010101010010: color_data = Z;
		19'b0011001010101010011: color_data = Z;
		19'b0011001010101010100: color_data = Z;
		19'b0011001010101010101: color_data = Z;
		19'b0011001010101010110: color_data = Z;
		19'b0011001010101010111: color_data = Z;
		19'b0011001010101011000: color_data = Z;
		19'b0011001010101011001: color_data = Z;
		19'b0011001010101011010: color_data = Z;
		19'b0011001010101011011: color_data = Z;
		19'b0011001010101011100: color_data = Z;
		19'b0011001010101011101: color_data = Z;
		19'b0011001010101011110: color_data = Z;
		19'b0011001010101011111: color_data = Z;
		19'b0011001010101100000: color_data = Z;
		19'b0011001010101100001: color_data = Z;
		19'b0011001010101100010: color_data = Z;
		19'b0011001010101100011: color_data = Z;
		19'b0011001010101100100: color_data = Z;
		19'b0011001010101100101: color_data = Z;
		19'b0011001010101100110: color_data = Z;
		19'b0011001010101100111: color_data = Z;
		19'b0011001010101101000: color_data = Z;
		19'b0011001010101101001: color_data = Z;
		19'b0011001010101101010: color_data = Z;
		19'b0011001010101101011: color_data = Z;
		19'b0011001010101101100: color_data = Z;
		19'b0011001010101101101: color_data = Z;
		19'b0011001010101101110: color_data = Z;
		19'b0011001010101101111: color_data = Z;
		19'b0011001010101110000: color_data = Z;
		19'b0011001010101110001: color_data = Z;
		19'b0011001010101110010: color_data = Z;
		19'b0011001010101110011: color_data = Z;
		19'b0011001010101110100: color_data = Z;
		19'b0011001010101110101: color_data = Z;
		19'b0011001010101110110: color_data = Z;
		19'b0011001010101110111: color_data = Z;
		19'b0011001010101111000: color_data = Z;
		19'b0011001010101111001: color_data = Z;
		19'b0011001010101111010: color_data = Z;
		19'b0011001010101111011: color_data = Z;
		19'b0011001010101111100: color_data = Z;
		19'b0011001010101111101: color_data = Z;
		19'b0011001010101111110: color_data = Z;
		19'b0011001010101111111: color_data = Z;
		19'b0011001010110000000: color_data = Z;
		19'b0011001010110000001: color_data = Z;
		19'b0011001010110000010: color_data = Z;
		19'b0011001010110000011: color_data = Z;
		19'b0011001010110000100: color_data = Z;
		19'b0011001010110000101: color_data = Z;
		19'b0011001010110000110: color_data = Z;
		19'b0011001010110000111: color_data = Z;
		19'b0011001010110001000: color_data = Z;
		19'b0011001010110001001: color_data = Z;
		19'b0011001010110001010: color_data = Z;
		19'b0011001010110001011: color_data = Z;
		19'b0011001010110001100: color_data = Z;
		19'b0011001010110001101: color_data = Z;
		19'b0011001010110001110: color_data = Z;
		19'b0011001010110001111: color_data = Z;
		19'b0011001010110010000: color_data = Z;
		19'b0011001010110010001: color_data = Z;
		19'b0011001010110010010: color_data = Z;
		19'b0011001010110010011: color_data = Z;
		19'b0011001010110010100: color_data = Z;
		19'b0011001010110010101: color_data = Z;
		19'b0011001010110010110: color_data = Z;
		19'b0011001010110010111: color_data = Z;
		19'b0011001010110011000: color_data = Z;
		19'b0011001010110011001: color_data = Z;
		19'b0011001010110011010: color_data = Z;
		19'b0011001010110011011: color_data = Z;
		19'b0011001010110011100: color_data = Z;
		19'b0011001010110011101: color_data = Z;
		19'b0011001010110011110: color_data = Z;
		19'b0011001010110011111: color_data = Z;
		19'b0011001010110100000: color_data = Z;
		19'b0011001010110100001: color_data = Z;
		19'b0011001010110100010: color_data = Z;
		19'b0011001010110100011: color_data = Z;
		19'b0011001010110100100: color_data = Z;
		19'b0011001010110100101: color_data = Z;
		19'b0011001010110100110: color_data = Z;
		19'b0011001010110100111: color_data = Z;
		19'b0011001010110101000: color_data = Z;
		19'b0011001010110101111: color_data = Z;
		19'b0011001010110110000: color_data = Z;
		19'b0011001010110110001: color_data = Z;
		19'b0011001010110110010: color_data = Z;
		19'b0011001010110110011: color_data = Z;
		19'b0011001010110110100: color_data = Z;
		19'b0011001010110110101: color_data = Z;
		19'b0011001010110110110: color_data = Z;
		19'b0011001010111001010: color_data = Z;
		19'b0011001100010110011: color_data = Z;
		19'b0011001100010110100: color_data = Z;
		19'b0011001100010110101: color_data = Z;
		19'b0011001100010110110: color_data = Z;
		19'b0011001100010110111: color_data = Z;
		19'b0011001100010111000: color_data = Z;
		19'b0011001100010111001: color_data = Z;
		19'b0011001100010111010: color_data = Z;
		19'b0011001100010111011: color_data = Z;
		19'b0011001100010111100: color_data = Z;
		19'b0011001100010111101: color_data = Z;
		19'b0011001100010111110: color_data = Z;
		19'b0011001100010111111: color_data = Z;
		19'b0011001100011000000: color_data = Z;
		19'b0011001100011000001: color_data = Z;
		19'b0011001100011000010: color_data = Z;
		19'b0011001100011000011: color_data = Z;
		19'b0011001100011000100: color_data = Z;
		19'b0011001100011000101: color_data = Z;
		19'b0011001100011000110: color_data = Z;
		19'b0011001100011000111: color_data = Z;
		19'b0011001100011001000: color_data = Z;
		19'b0011001100011001001: color_data = Z;
		19'b0011001100011001010: color_data = Z;
		19'b0011001100011001011: color_data = Z;
		19'b0011001100011001100: color_data = Z;
		19'b0011001100011001101: color_data = Z;
		19'b0011001100011001110: color_data = Z;
		19'b0011001100011001111: color_data = Z;
		19'b0011001100011010000: color_data = Z;
		19'b0011001100011010001: color_data = Z;
		19'b0011001100011010010: color_data = Z;
		19'b0011001100011010011: color_data = Z;
		19'b0011001100011010100: color_data = Z;
		19'b0011001100011010101: color_data = Z;
		19'b0011001100011010110: color_data = Z;
		19'b0011001100011010111: color_data = Z;
		19'b0011001100011011000: color_data = Z;
		19'b0011001100011011001: color_data = Z;
		19'b0011001100011011010: color_data = Z;
		19'b0011001100011011011: color_data = Z;
		19'b0011001100011011100: color_data = Z;
		19'b0011001100011011101: color_data = Z;
		19'b0011001100011011110: color_data = Z;
		19'b0011001100011011111: color_data = Z;
		19'b0011001100011100000: color_data = Z;
		19'b0011001100011100001: color_data = Z;
		19'b0011001100011100010: color_data = Z;
		19'b0011001100011100011: color_data = Z;
		19'b0011001100011100100: color_data = Z;
		19'b0011001100011100101: color_data = Z;
		19'b0011001100011100110: color_data = Z;
		19'b0011001100011100111: color_data = Z;
		19'b0011001100011101000: color_data = Z;
		19'b0011001100011101001: color_data = Z;
		19'b0011001100011101010: color_data = Z;
		19'b0011001100011101011: color_data = Z;
		19'b0011001100011101100: color_data = Z;
		19'b0011001100011101101: color_data = Z;
		19'b0011001100011101110: color_data = Z;
		19'b0011001100011101111: color_data = Z;
		19'b0011001100011110000: color_data = Z;
		19'b0011001100011110001: color_data = Z;
		19'b0011001100011110010: color_data = Z;
		19'b0011001100011110011: color_data = Z;
		19'b0011001100011110100: color_data = Z;
		19'b0011001100011110101: color_data = Z;
		19'b0011001100011110110: color_data = Z;
		19'b0011001100011110111: color_data = Z;
		19'b0011001100011111000: color_data = Z;
		19'b0011001100011111001: color_data = Z;
		19'b0011001100011111010: color_data = Z;
		19'b0011001100011111011: color_data = Z;
		19'b0011001100011111100: color_data = Z;
		19'b0011001100011111101: color_data = Z;
		19'b0011001100011111110: color_data = Z;
		19'b0011001100011111111: color_data = Z;
		19'b0011001100100000000: color_data = Z;
		19'b0011001100100000001: color_data = Z;
		19'b0011001100100000010: color_data = Z;
		19'b0011001100100000011: color_data = Z;
		19'b0011001100100000100: color_data = Z;
		19'b0011001100100000101: color_data = Z;
		19'b0011001100100000110: color_data = Z;
		19'b0011001100100000111: color_data = Z;
		19'b0011001100100001000: color_data = Z;
		19'b0011001100100001001: color_data = Z;
		19'b0011001100100001010: color_data = Z;
		19'b0011001100100001011: color_data = Z;
		19'b0011001100100001100: color_data = Z;
		19'b0011001100100001101: color_data = Z;
		19'b0011001100100001110: color_data = Z;
		19'b0011001100100001111: color_data = Z;
		19'b0011001100100010000: color_data = Z;
		19'b0011001100100010001: color_data = Z;
		19'b0011001100100010010: color_data = Z;
		19'b0011001100100010011: color_data = Z;
		19'b0011001100100010100: color_data = Z;
		19'b0011001100100010101: color_data = Z;
		19'b0011001100100010110: color_data = Z;
		19'b0011001100100010111: color_data = Z;
		19'b0011001100100011000: color_data = Z;
		19'b0011001100100011001: color_data = Z;
		19'b0011001100100011010: color_data = Z;
		19'b0011001100100011011: color_data = Z;
		19'b0011001100100011100: color_data = Z;
		19'b0011001100100011101: color_data = Z;
		19'b0011001100100011110: color_data = Z;
		19'b0011001100100011111: color_data = Z;
		19'b0011001100100100000: color_data = Z;
		19'b0011001100100100001: color_data = Z;
		19'b0011001100100100010: color_data = Z;
		19'b0011001100100100011: color_data = Z;
		19'b0011001100100100100: color_data = Z;
		19'b0011001100100100101: color_data = Z;
		19'b0011001100100100110: color_data = Z;
		19'b0011001100100100111: color_data = Z;
		19'b0011001100100101000: color_data = Z;
		19'b0011001100100101001: color_data = Z;
		19'b0011001100100101010: color_data = Z;
		19'b0011001100100101011: color_data = Z;
		19'b0011001100100101100: color_data = Z;
		19'b0011001100100101101: color_data = Z;
		19'b0011001100100101110: color_data = Z;
		19'b0011001100100101111: color_data = Z;
		19'b0011001100100110000: color_data = Z;
		19'b0011001100100110001: color_data = Z;
		19'b0011001100100110010: color_data = Z;
		19'b0011001100100110011: color_data = Z;
		19'b0011001100100110100: color_data = Z;
		19'b0011001100100110101: color_data = Z;
		19'b0011001100100110110: color_data = Z;
		19'b0011001100100110111: color_data = Z;
		19'b0011001100100111000: color_data = Z;
		19'b0011001100100111001: color_data = Z;
		19'b0011001100100111010: color_data = Z;
		19'b0011001100100111011: color_data = Z;
		19'b0011001100100111100: color_data = Z;
		19'b0011001100100111101: color_data = Z;
		19'b0011001100100111110: color_data = Z;
		19'b0011001100100111111: color_data = Z;
		19'b0011001100101000000: color_data = Z;
		19'b0011001100101000001: color_data = Z;
		19'b0011001100101000010: color_data = Z;
		19'b0011001100101000011: color_data = Z;
		19'b0011001100101000100: color_data = Z;
		19'b0011001100101000101: color_data = Z;
		19'b0011001100101000110: color_data = Z;
		19'b0011001100101000111: color_data = Z;
		19'b0011001100101001000: color_data = Z;
		19'b0011001100101001001: color_data = Z;
		19'b0011001100101001010: color_data = Z;
		19'b0011001100101001011: color_data = Z;
		19'b0011001100101001100: color_data = Z;
		19'b0011001100101001101: color_data = Z;
		19'b0011001100101001110: color_data = Z;
		19'b0011001100101001111: color_data = Z;
		19'b0011001100101010000: color_data = Z;
		19'b0011001100101010001: color_data = Z;
		19'b0011001100101010010: color_data = Z;
		19'b0011001100101010011: color_data = Z;
		19'b0011001100101010100: color_data = Z;
		19'b0011001100101010101: color_data = Z;
		19'b0011001100101010110: color_data = Z;
		19'b0011001100101010111: color_data = Z;
		19'b0011001100101011000: color_data = Z;
		19'b0011001100101011001: color_data = Z;
		19'b0011001100101011010: color_data = Z;
		19'b0011001100101011011: color_data = Z;
		19'b0011001100101011100: color_data = Z;
		19'b0011001100101011101: color_data = Z;
		19'b0011001100101011110: color_data = Z;
		19'b0011001100101011111: color_data = Z;
		19'b0011001100101100000: color_data = Z;
		19'b0011001100101100001: color_data = Z;
		19'b0011001100101100010: color_data = Z;
		19'b0011001100101100011: color_data = Z;
		19'b0011001100101100100: color_data = Z;
		19'b0011001100101100101: color_data = Z;
		19'b0011001100101100110: color_data = Z;
		19'b0011001100101100111: color_data = Z;
		19'b0011001100101101000: color_data = Z;
		19'b0011001100101101001: color_data = Z;
		19'b0011001100101101010: color_data = Z;
		19'b0011001100101101011: color_data = Z;
		19'b0011001100101101100: color_data = Z;
		19'b0011001100101101101: color_data = Z;
		19'b0011001100101101110: color_data = Z;
		19'b0011001100101101111: color_data = Z;
		19'b0011001100101110000: color_data = Z;
		19'b0011001100101110001: color_data = Z;
		19'b0011001100101110010: color_data = Z;
		19'b0011001100101110011: color_data = Z;
		19'b0011001100101110100: color_data = Z;
		19'b0011001100101110101: color_data = Z;
		19'b0011001100101110110: color_data = Z;
		19'b0011001100101110111: color_data = Z;
		19'b0011001100101111000: color_data = Z;
		19'b0011001100101111001: color_data = Z;
		19'b0011001100101111010: color_data = Z;
		19'b0011001100101111011: color_data = Z;
		19'b0011001100101111100: color_data = Z;
		19'b0011001100101111101: color_data = Z;
		19'b0011001100101111110: color_data = Z;
		19'b0011001100101111111: color_data = Z;
		19'b0011001100110000000: color_data = Z;
		19'b0011001100110000001: color_data = Z;
		19'b0011001100110000010: color_data = Z;
		19'b0011001100110000011: color_data = Z;
		19'b0011001100110000100: color_data = Z;
		19'b0011001100110000101: color_data = Z;
		19'b0011001100110000110: color_data = Z;
		19'b0011001100110000111: color_data = Z;
		19'b0011001100110001000: color_data = Z;
		19'b0011001100110001001: color_data = Z;
		19'b0011001100110001010: color_data = Z;
		19'b0011001100110001011: color_data = Z;
		19'b0011001100110001100: color_data = Z;
		19'b0011001100110001101: color_data = Z;
		19'b0011001100110001110: color_data = Z;
		19'b0011001100110001111: color_data = Z;
		19'b0011001100110010000: color_data = Z;
		19'b0011001100110010001: color_data = Z;
		19'b0011001100110010010: color_data = Z;
		19'b0011001100110010011: color_data = Z;
		19'b0011001100110010100: color_data = Z;
		19'b0011001100110010101: color_data = Z;
		19'b0011001100110010110: color_data = Z;
		19'b0011001100110010111: color_data = Z;
		19'b0011001100110011000: color_data = Z;
		19'b0011001100110011001: color_data = Z;
		19'b0011001100110011010: color_data = Z;
		19'b0011001100110011011: color_data = Z;
		19'b0011001100110011100: color_data = Z;
		19'b0011001100110011101: color_data = Z;
		19'b0011001100110011110: color_data = Z;
		19'b0011001100110011111: color_data = Z;
		19'b0011001100110100000: color_data = Z;
		19'b0011001100110100001: color_data = Z;
		19'b0011001100110100010: color_data = Z;
		19'b0011001100110100011: color_data = Z;
		19'b0011001100110110000: color_data = Z;
		19'b0011001100110110001: color_data = Z;
		19'b0011001100110110010: color_data = Z;
		19'b0011001100110110011: color_data = Z;
		19'b0011001100110110100: color_data = Z;
		19'b0011001100110110101: color_data = Z;
		19'b0011001100110110110: color_data = Z;
		19'b0011001100110110111: color_data = Z;
		19'b0011001110010110010: color_data = Z;
		19'b0011001110010110011: color_data = Z;
		19'b0011001110010110100: color_data = Z;
		19'b0011001110010110101: color_data = Z;
		19'b0011001110010110110: color_data = Z;
		19'b0011001110010110111: color_data = Z;
		19'b0011001110010111000: color_data = Z;
		19'b0011001110010111001: color_data = Z;
		19'b0011001110010111010: color_data = Z;
		19'b0011001110010111011: color_data = Z;
		19'b0011001110010111100: color_data = Z;
		19'b0011001110010111101: color_data = Z;
		19'b0011001110010111110: color_data = Z;
		19'b0011001110010111111: color_data = Z;
		19'b0011001110011000000: color_data = Z;
		19'b0011001110011000001: color_data = Z;
		19'b0011001110011000010: color_data = Z;
		19'b0011001110011000011: color_data = Z;
		19'b0011001110011000100: color_data = Z;
		19'b0011001110011000101: color_data = Z;
		19'b0011001110011000110: color_data = Z;
		19'b0011001110011000111: color_data = Z;
		19'b0011001110011001000: color_data = Z;
		19'b0011001110011001001: color_data = Z;
		19'b0011001110011001010: color_data = Z;
		19'b0011001110011001011: color_data = Z;
		19'b0011001110011001100: color_data = Z;
		19'b0011001110011001101: color_data = Z;
		19'b0011001110011001110: color_data = Z;
		19'b0011001110011001111: color_data = Z;
		19'b0011001110011010000: color_data = Z;
		19'b0011001110011010001: color_data = Z;
		19'b0011001110011010010: color_data = Z;
		19'b0011001110011010011: color_data = Z;
		19'b0011001110011010100: color_data = Z;
		19'b0011001110011010101: color_data = Z;
		19'b0011001110011010110: color_data = Z;
		19'b0011001110011010111: color_data = Z;
		19'b0011001110011011000: color_data = Z;
		19'b0011001110011011001: color_data = Z;
		19'b0011001110011011010: color_data = Z;
		19'b0011001110011011011: color_data = Z;
		19'b0011001110011011100: color_data = Z;
		19'b0011001110011011101: color_data = Z;
		19'b0011001110011011110: color_data = Z;
		19'b0011001110011011111: color_data = Z;
		19'b0011001110011100000: color_data = Z;
		19'b0011001110011100001: color_data = Z;
		19'b0011001110011100010: color_data = Z;
		19'b0011001110011100011: color_data = Z;
		19'b0011001110011100100: color_data = Z;
		19'b0011001110011100101: color_data = Z;
		19'b0011001110011100110: color_data = Z;
		19'b0011001110011100111: color_data = Z;
		19'b0011001110011101000: color_data = Z;
		19'b0011001110011101001: color_data = Z;
		19'b0011001110011101010: color_data = Z;
		19'b0011001110011101011: color_data = Z;
		19'b0011001110011101100: color_data = Z;
		19'b0011001110011101101: color_data = Z;
		19'b0011001110011101110: color_data = Z;
		19'b0011001110011101111: color_data = Z;
		19'b0011001110011110000: color_data = Z;
		19'b0011001110011110001: color_data = Z;
		19'b0011001110011110010: color_data = Z;
		19'b0011001110011110011: color_data = Z;
		19'b0011001110011110100: color_data = Z;
		19'b0011001110011110101: color_data = Z;
		19'b0011001110011110110: color_data = Z;
		19'b0011001110011110111: color_data = Z;
		19'b0011001110011111000: color_data = Z;
		19'b0011001110011111001: color_data = Z;
		19'b0011001110011111010: color_data = Z;
		19'b0011001110011111011: color_data = Z;
		19'b0011001110011111100: color_data = Z;
		19'b0011001110011111101: color_data = Z;
		19'b0011001110011111110: color_data = Z;
		19'b0011001110011111111: color_data = Z;
		19'b0011001110100000000: color_data = Z;
		19'b0011001110100000001: color_data = Z;
		19'b0011001110100000010: color_data = Z;
		19'b0011001110100000011: color_data = Z;
		19'b0011001110100000100: color_data = Z;
		19'b0011001110100000101: color_data = Z;
		19'b0011001110100000110: color_data = Z;
		19'b0011001110100000111: color_data = Z;
		19'b0011001110100001000: color_data = Z;
		19'b0011001110100001001: color_data = Z;
		19'b0011001110100001010: color_data = Z;
		19'b0011001110100001011: color_data = Z;
		19'b0011001110100001100: color_data = Z;
		19'b0011001110100001101: color_data = Z;
		19'b0011001110100001110: color_data = Z;
		19'b0011001110100001111: color_data = Z;
		19'b0011001110100010000: color_data = Z;
		19'b0011001110100010001: color_data = Z;
		19'b0011001110100010010: color_data = Z;
		19'b0011001110100010011: color_data = Z;
		19'b0011001110100010100: color_data = Z;
		19'b0011001110100010101: color_data = Z;
		19'b0011001110100010110: color_data = Z;
		19'b0011001110100010111: color_data = Z;
		19'b0011001110100011000: color_data = Z;
		19'b0011001110100011001: color_data = Z;
		19'b0011001110100011010: color_data = Z;
		19'b0011001110100011011: color_data = Z;
		19'b0011001110100011100: color_data = Z;
		19'b0011001110100011101: color_data = Z;
		19'b0011001110100011110: color_data = Z;
		19'b0011001110100011111: color_data = Z;
		19'b0011001110100100000: color_data = Z;
		19'b0011001110100100001: color_data = Z;
		19'b0011001110100100010: color_data = Z;
		19'b0011001110100100011: color_data = Z;
		19'b0011001110100100100: color_data = Z;
		19'b0011001110100100101: color_data = Z;
		19'b0011001110100100110: color_data = Z;
		19'b0011001110100100111: color_data = Z;
		19'b0011001110100101000: color_data = Z;
		19'b0011001110100101001: color_data = Z;
		19'b0011001110100101010: color_data = Z;
		19'b0011001110100101011: color_data = Z;
		19'b0011001110100101100: color_data = Z;
		19'b0011001110100101101: color_data = Z;
		19'b0011001110100101110: color_data = Z;
		19'b0011001110100101111: color_data = Z;
		19'b0011001110100110000: color_data = Z;
		19'b0011001110100110001: color_data = Z;
		19'b0011001110100110010: color_data = Z;
		19'b0011001110100110011: color_data = Z;
		19'b0011001110100110100: color_data = Z;
		19'b0011001110100110101: color_data = Z;
		19'b0011001110100110110: color_data = Z;
		19'b0011001110100110111: color_data = Z;
		19'b0011001110100111000: color_data = Z;
		19'b0011001110100111001: color_data = Z;
		19'b0011001110100111010: color_data = Z;
		19'b0011001110100111011: color_data = Z;
		19'b0011001110100111100: color_data = Z;
		19'b0011001110100111101: color_data = Z;
		19'b0011001110100111110: color_data = Z;
		19'b0011001110100111111: color_data = Z;
		19'b0011001110101000000: color_data = Z;
		19'b0011001110101000001: color_data = Z;
		19'b0011001110101000010: color_data = Z;
		19'b0011001110101000011: color_data = Z;
		19'b0011001110101000100: color_data = Z;
		19'b0011001110101000101: color_data = Z;
		19'b0011001110101000110: color_data = Z;
		19'b0011001110101000111: color_data = Z;
		19'b0011001110101001000: color_data = Z;
		19'b0011001110101001001: color_data = Z;
		19'b0011001110101001010: color_data = Z;
		19'b0011001110101001011: color_data = Z;
		19'b0011001110101001100: color_data = Z;
		19'b0011001110101001101: color_data = Z;
		19'b0011001110101001110: color_data = Z;
		19'b0011001110101001111: color_data = Z;
		19'b0011001110101010000: color_data = Z;
		19'b0011001110101010001: color_data = Z;
		19'b0011001110101010010: color_data = Z;
		19'b0011001110101010011: color_data = Z;
		19'b0011001110101010100: color_data = Z;
		19'b0011001110101010101: color_data = Z;
		19'b0011001110101010110: color_data = Z;
		19'b0011001110101010111: color_data = Z;
		19'b0011001110101011000: color_data = Z;
		19'b0011001110101011001: color_data = Z;
		19'b0011001110101011010: color_data = Z;
		19'b0011001110101011011: color_data = Z;
		19'b0011001110101011100: color_data = Z;
		19'b0011001110101011101: color_data = Z;
		19'b0011001110101011110: color_data = Z;
		19'b0011001110101011111: color_data = Z;
		19'b0011001110101100000: color_data = Z;
		19'b0011001110101100001: color_data = Z;
		19'b0011001110101100010: color_data = Z;
		19'b0011001110101100011: color_data = Z;
		19'b0011001110101100100: color_data = Z;
		19'b0011001110101100101: color_data = Z;
		19'b0011001110101100110: color_data = Z;
		19'b0011001110101100111: color_data = Z;
		19'b0011001110101101000: color_data = Z;
		19'b0011001110101101001: color_data = Z;
		19'b0011001110101101010: color_data = Z;
		19'b0011001110101101011: color_data = Z;
		19'b0011001110101101100: color_data = Z;
		19'b0011001110101101101: color_data = Z;
		19'b0011001110101101110: color_data = Z;
		19'b0011001110101101111: color_data = Z;
		19'b0011001110101110000: color_data = Z;
		19'b0011001110101110001: color_data = Z;
		19'b0011001110101110010: color_data = Z;
		19'b0011001110101110011: color_data = Z;
		19'b0011001110101110100: color_data = Z;
		19'b0011001110101110101: color_data = Z;
		19'b0011001110101110110: color_data = Z;
		19'b0011001110101110111: color_data = Z;
		19'b0011001110101111000: color_data = Z;
		19'b0011001110101111001: color_data = Z;
		19'b0011001110101111010: color_data = Z;
		19'b0011001110101111011: color_data = Z;
		19'b0011001110101111100: color_data = Z;
		19'b0011001110101111101: color_data = Z;
		19'b0011001110101111110: color_data = Z;
		19'b0011001110101111111: color_data = Z;
		19'b0011001110110000000: color_data = Z;
		19'b0011001110110000001: color_data = Z;
		19'b0011001110110000010: color_data = Z;
		19'b0011001110110000011: color_data = Z;
		19'b0011001110110000100: color_data = Z;
		19'b0011001110110000101: color_data = Z;
		19'b0011001110110000110: color_data = Z;
		19'b0011001110110000111: color_data = Z;
		19'b0011001110110001000: color_data = Z;
		19'b0011001110110001001: color_data = Z;
		19'b0011001110110001010: color_data = Z;
		19'b0011001110110001011: color_data = Z;
		19'b0011001110110001100: color_data = Z;
		19'b0011001110110001101: color_data = Z;
		19'b0011001110110001110: color_data = Z;
		19'b0011001110110001111: color_data = Z;
		19'b0011001110110010000: color_data = Z;
		19'b0011001110110010001: color_data = Z;
		19'b0011001110110010010: color_data = Z;
		19'b0011001110110010011: color_data = Z;
		19'b0011001110110010100: color_data = Z;
		19'b0011001110110010101: color_data = Z;
		19'b0011001110110010110: color_data = Z;
		19'b0011001110110010111: color_data = Z;
		19'b0011001110110011000: color_data = Z;
		19'b0011001110110011001: color_data = Z;
		19'b0011001110110011010: color_data = Z;
		19'b0011001110110011011: color_data = Z;
		19'b0011001110110011100: color_data = Z;
		19'b0011001110110011101: color_data = Z;
		19'b0011001110110011110: color_data = Z;
		19'b0011001110110101111: color_data = Z;
		19'b0011001110110110000: color_data = Z;
		19'b0011001110110110001: color_data = Z;
		19'b0011001110110110010: color_data = Z;
		19'b0011001110110110011: color_data = Z;
		19'b0011001110110110100: color_data = Z;
		19'b0011001110110110101: color_data = Z;
		19'b0011001110110110110: color_data = Z;
		19'b0011001110110110111: color_data = Z;
		19'b0011001110110111000: color_data = Z;
		19'b0011010000010110001: color_data = Z;
		19'b0011010000010110010: color_data = Z;
		19'b0011010000010110011: color_data = Z;
		19'b0011010000010110100: color_data = Z;
		19'b0011010000010110101: color_data = Z;
		19'b0011010000010110110: color_data = Z;
		19'b0011010000010110111: color_data = Z;
		19'b0011010000010111000: color_data = Z;
		19'b0011010000010111001: color_data = Z;
		19'b0011010000010111010: color_data = Z;
		19'b0011010000010111011: color_data = Z;
		19'b0011010000010111100: color_data = Z;
		19'b0011010000010111101: color_data = Z;
		19'b0011010000010111110: color_data = Z;
		19'b0011010000010111111: color_data = Z;
		19'b0011010000011000000: color_data = Z;
		19'b0011010000011000001: color_data = Z;
		19'b0011010000011000010: color_data = Z;
		19'b0011010000011000011: color_data = Z;
		19'b0011010000011000100: color_data = Z;
		19'b0011010000011000101: color_data = Z;
		19'b0011010000011000110: color_data = Z;
		19'b0011010000011000111: color_data = Z;
		19'b0011010000011001000: color_data = Z;
		19'b0011010000011001001: color_data = Z;
		19'b0011010000011001010: color_data = Z;
		19'b0011010000011001011: color_data = Z;
		19'b0011010000011001100: color_data = Z;
		19'b0011010000011001101: color_data = Z;
		19'b0011010000011001110: color_data = Z;
		19'b0011010000011001111: color_data = Z;
		19'b0011010000011010000: color_data = Z;
		19'b0011010000011010001: color_data = Z;
		19'b0011010000011010010: color_data = Z;
		19'b0011010000011010011: color_data = Z;
		19'b0011010000011010100: color_data = Z;
		19'b0011010000011010101: color_data = Z;
		19'b0011010000011010110: color_data = Z;
		19'b0011010000011010111: color_data = Z;
		19'b0011010000011011000: color_data = Z;
		19'b0011010000011011001: color_data = Z;
		19'b0011010000011011010: color_data = Z;
		19'b0011010000011011011: color_data = Z;
		19'b0011010000011011100: color_data = Z;
		19'b0011010000011011101: color_data = Z;
		19'b0011010000011011110: color_data = Z;
		19'b0011010000011011111: color_data = Z;
		19'b0011010000011100000: color_data = Z;
		19'b0011010000011100001: color_data = Z;
		19'b0011010000011100010: color_data = Z;
		19'b0011010000011100011: color_data = Z;
		19'b0011010000011100100: color_data = Z;
		19'b0011010000011100101: color_data = Z;
		19'b0011010000011100110: color_data = Z;
		19'b0011010000011100111: color_data = Z;
		19'b0011010000011101000: color_data = Z;
		19'b0011010000011101001: color_data = Z;
		19'b0011010000011101010: color_data = Z;
		19'b0011010000011101011: color_data = Z;
		19'b0011010000011101100: color_data = Z;
		19'b0011010000011101101: color_data = Z;
		19'b0011010000011101110: color_data = Z;
		19'b0011010000011101111: color_data = Z;
		19'b0011010000011110000: color_data = Z;
		19'b0011010000011110001: color_data = Z;
		19'b0011010000011110010: color_data = Z;
		19'b0011010000011110011: color_data = Z;
		19'b0011010000011110100: color_data = Z;
		19'b0011010000011110101: color_data = Z;
		19'b0011010000011110110: color_data = Z;
		19'b0011010000011110111: color_data = Z;
		19'b0011010000011111000: color_data = Z;
		19'b0011010000011111001: color_data = Z;
		19'b0011010000011111010: color_data = Z;
		19'b0011010000011111011: color_data = Z;
		19'b0011010000011111100: color_data = Z;
		19'b0011010000011111101: color_data = Z;
		19'b0011010000011111110: color_data = Z;
		19'b0011010000011111111: color_data = Z;
		19'b0011010000100000000: color_data = Z;
		19'b0011010000100000001: color_data = Z;
		19'b0011010000100000010: color_data = Z;
		19'b0011010000100000011: color_data = Z;
		19'b0011010000100000100: color_data = Z;
		19'b0011010000100000101: color_data = Z;
		19'b0011010000100000110: color_data = Z;
		19'b0011010000100000111: color_data = Z;
		19'b0011010000100001000: color_data = Z;
		19'b0011010000100001001: color_data = Z;
		19'b0011010000100001010: color_data = Z;
		19'b0011010000100001011: color_data = Z;
		19'b0011010000100001100: color_data = Z;
		19'b0011010000100001101: color_data = Z;
		19'b0011010000100001110: color_data = Z;
		19'b0011010000100001111: color_data = Z;
		19'b0011010000100010000: color_data = Z;
		19'b0011010000100010001: color_data = Z;
		19'b0011010000100010010: color_data = Z;
		19'b0011010000100010011: color_data = Z;
		19'b0011010000100010100: color_data = Z;
		19'b0011010000100010101: color_data = Z;
		19'b0011010000100010110: color_data = Z;
		19'b0011010000100010111: color_data = Z;
		19'b0011010000100011000: color_data = Z;
		19'b0011010000100011001: color_data = Z;
		19'b0011010000100011010: color_data = Z;
		19'b0011010000100011011: color_data = Z;
		19'b0011010000100011100: color_data = Z;
		19'b0011010000100011101: color_data = Z;
		19'b0011010000100011110: color_data = Z;
		19'b0011010000100011111: color_data = Z;
		19'b0011010000100100000: color_data = Z;
		19'b0011010000100100001: color_data = Z;
		19'b0011010000100100010: color_data = Z;
		19'b0011010000100100011: color_data = Z;
		19'b0011010000100100100: color_data = Z;
		19'b0011010000100100101: color_data = Z;
		19'b0011010000100100110: color_data = Z;
		19'b0011010000100100111: color_data = Z;
		19'b0011010000100101000: color_data = Z;
		19'b0011010000100101001: color_data = Z;
		19'b0011010000100101010: color_data = Z;
		19'b0011010000100101011: color_data = Z;
		19'b0011010000100101100: color_data = Z;
		19'b0011010000100101101: color_data = Z;
		19'b0011010000100101110: color_data = Z;
		19'b0011010000100101111: color_data = Z;
		19'b0011010000100110000: color_data = Z;
		19'b0011010000100110001: color_data = Z;
		19'b0011010000100110010: color_data = Z;
		19'b0011010000100110011: color_data = Z;
		19'b0011010000100110100: color_data = Z;
		19'b0011010000100110101: color_data = Z;
		19'b0011010000100110110: color_data = Z;
		19'b0011010000100110111: color_data = Z;
		19'b0011010000100111000: color_data = Z;
		19'b0011010000100111001: color_data = Z;
		19'b0011010000100111010: color_data = Z;
		19'b0011010000100111011: color_data = Z;
		19'b0011010000100111100: color_data = Z;
		19'b0011010000100111101: color_data = Z;
		19'b0011010000100111110: color_data = Z;
		19'b0011010000100111111: color_data = Z;
		19'b0011010000101000000: color_data = Z;
		19'b0011010000101000001: color_data = Z;
		19'b0011010000101000010: color_data = Z;
		19'b0011010000101000011: color_data = Z;
		19'b0011010000101000100: color_data = Z;
		19'b0011010000101000101: color_data = Z;
		19'b0011010000101000110: color_data = Z;
		19'b0011010000101000111: color_data = Z;
		19'b0011010000101001000: color_data = Z;
		19'b0011010000101001001: color_data = Z;
		19'b0011010000101001010: color_data = Z;
		19'b0011010000101001011: color_data = Z;
		19'b0011010000101001100: color_data = Z;
		19'b0011010000101001101: color_data = Z;
		19'b0011010000101001110: color_data = Z;
		19'b0011010000101001111: color_data = Z;
		19'b0011010000101010000: color_data = Z;
		19'b0011010000101010001: color_data = Z;
		19'b0011010000101010010: color_data = Z;
		19'b0011010000101010011: color_data = Z;
		19'b0011010000101010100: color_data = Z;
		19'b0011010000101010101: color_data = Z;
		19'b0011010000101010110: color_data = Z;
		19'b0011010000101010111: color_data = Z;
		19'b0011010000101011000: color_data = Z;
		19'b0011010000101011001: color_data = Z;
		19'b0011010000101011010: color_data = Z;
		19'b0011010000101011011: color_data = Z;
		19'b0011010000101011100: color_data = Z;
		19'b0011010000101011101: color_data = Z;
		19'b0011010000101011110: color_data = Z;
		19'b0011010000101011111: color_data = Z;
		19'b0011010000101100000: color_data = Z;
		19'b0011010000101100001: color_data = Z;
		19'b0011010000101100010: color_data = Z;
		19'b0011010000101100011: color_data = Z;
		19'b0011010000101100100: color_data = Z;
		19'b0011010000101100101: color_data = Z;
		19'b0011010000101100110: color_data = Z;
		19'b0011010000101100111: color_data = Z;
		19'b0011010000101101000: color_data = Z;
		19'b0011010000101101001: color_data = Z;
		19'b0011010000101101010: color_data = Z;
		19'b0011010000101101011: color_data = Z;
		19'b0011010000101101100: color_data = Z;
		19'b0011010000101101101: color_data = Z;
		19'b0011010000101101110: color_data = Z;
		19'b0011010000101101111: color_data = Z;
		19'b0011010000101110000: color_data = Z;
		19'b0011010000101110001: color_data = Z;
		19'b0011010000101110010: color_data = Z;
		19'b0011010000101110011: color_data = Z;
		19'b0011010000101110100: color_data = Z;
		19'b0011010000101110101: color_data = Z;
		19'b0011010000101110110: color_data = Z;
		19'b0011010000101110111: color_data = Z;
		19'b0011010000101111000: color_data = Z;
		19'b0011010000101111001: color_data = Z;
		19'b0011010000101111010: color_data = Z;
		19'b0011010000101111011: color_data = Z;
		19'b0011010000101111100: color_data = Z;
		19'b0011010000101111101: color_data = Z;
		19'b0011010000101111110: color_data = Z;
		19'b0011010000101111111: color_data = Z;
		19'b0011010000110000000: color_data = Z;
		19'b0011010000110000001: color_data = Z;
		19'b0011010000110000010: color_data = Z;
		19'b0011010000110000011: color_data = Z;
		19'b0011010000110000100: color_data = Z;
		19'b0011010000110000101: color_data = Z;
		19'b0011010000110000110: color_data = Z;
		19'b0011010000110000111: color_data = Z;
		19'b0011010000110001000: color_data = Z;
		19'b0011010000110001001: color_data = Z;
		19'b0011010000110001010: color_data = Z;
		19'b0011010000110001011: color_data = Z;
		19'b0011010000110001100: color_data = Z;
		19'b0011010000110001101: color_data = Z;
		19'b0011010000110001110: color_data = Z;
		19'b0011010000110001111: color_data = Z;
		19'b0011010000110010000: color_data = Z;
		19'b0011010000110010001: color_data = Z;
		19'b0011010000110010010: color_data = Z;
		19'b0011010000110010011: color_data = Z;
		19'b0011010000110010100: color_data = Z;
		19'b0011010000110010101: color_data = Z;
		19'b0011010000110010110: color_data = Z;
		19'b0011010000110010111: color_data = Z;
		19'b0011010000110011000: color_data = Z;
		19'b0011010000110011001: color_data = Z;
		19'b0011010000110011010: color_data = Z;
		19'b0011010000110011011: color_data = Z;
		19'b0011010000110011100: color_data = Z;
		19'b0011010000110110011: color_data = Z;
		19'b0011010000110110100: color_data = Z;
		19'b0011010000110110101: color_data = Z;
		19'b0011010000110110110: color_data = Z;
		19'b0011010000110110111: color_data = Z;
		19'b0011010000110111000: color_data = Z;
		19'b0011010000111010011: color_data = Z;
		19'b0011010000111011000: color_data = Z;
		19'b0011010010010110001: color_data = Z;
		19'b0011010010010110010: color_data = Z;
		19'b0011010010010110011: color_data = Z;
		19'b0011010010010110100: color_data = Z;
		19'b0011010010010110101: color_data = Z;
		19'b0011010010010110110: color_data = Z;
		19'b0011010010010110111: color_data = Z;
		19'b0011010010010111000: color_data = Z;
		19'b0011010010010111001: color_data = Z;
		19'b0011010010010111010: color_data = Z;
		19'b0011010010010111011: color_data = Z;
		19'b0011010010010111100: color_data = Z;
		19'b0011010010010111101: color_data = Z;
		19'b0011010010010111110: color_data = Z;
		19'b0011010010010111111: color_data = Z;
		19'b0011010010011000000: color_data = Z;
		19'b0011010010011000001: color_data = Z;
		19'b0011010010011000010: color_data = Z;
		19'b0011010010011000011: color_data = Z;
		19'b0011010010011000100: color_data = Z;
		19'b0011010010011000101: color_data = Z;
		19'b0011010010011000110: color_data = Z;
		19'b0011010010011000111: color_data = Z;
		19'b0011010010011001000: color_data = Z;
		19'b0011010010011001001: color_data = Z;
		19'b0011010010011001010: color_data = Z;
		19'b0011010010011001011: color_data = Z;
		19'b0011010010011001100: color_data = Z;
		19'b0011010010011001101: color_data = Z;
		19'b0011010010011001110: color_data = Z;
		19'b0011010010011001111: color_data = Z;
		19'b0011010010011010000: color_data = Z;
		19'b0011010010011010001: color_data = Z;
		19'b0011010010011010010: color_data = Z;
		19'b0011010010011010011: color_data = Z;
		19'b0011010010011010100: color_data = Z;
		19'b0011010010011010101: color_data = Z;
		19'b0011010010011010110: color_data = Z;
		19'b0011010010011010111: color_data = Z;
		19'b0011010010011011000: color_data = Z;
		19'b0011010010011011001: color_data = Z;
		19'b0011010010011011010: color_data = Z;
		19'b0011010010011011011: color_data = Z;
		19'b0011010010011011100: color_data = Z;
		19'b0011010010011011101: color_data = Z;
		19'b0011010010011011110: color_data = Z;
		19'b0011010010011011111: color_data = Z;
		19'b0011010010011100000: color_data = Z;
		19'b0011010010011100001: color_data = Z;
		19'b0011010010011100010: color_data = Z;
		19'b0011010010011100011: color_data = Z;
		19'b0011010010011100100: color_data = Z;
		19'b0011010010011100101: color_data = Z;
		19'b0011010010011100110: color_data = Z;
		19'b0011010010011100111: color_data = Z;
		19'b0011010010011101000: color_data = Z;
		19'b0011010010011101001: color_data = Z;
		19'b0011010010011101010: color_data = Z;
		19'b0011010010011101011: color_data = Z;
		19'b0011010010011101100: color_data = Z;
		19'b0011010010011101101: color_data = Z;
		19'b0011010010011101110: color_data = Z;
		19'b0011010010011101111: color_data = Z;
		19'b0011010010011110000: color_data = Z;
		19'b0011010010011110001: color_data = Z;
		19'b0011010010011110010: color_data = Z;
		19'b0011010010011110011: color_data = Z;
		19'b0011010010011110100: color_data = Z;
		19'b0011010010011110101: color_data = Z;
		19'b0011010010011110110: color_data = Z;
		19'b0011010010011110111: color_data = Z;
		19'b0011010010011111000: color_data = Z;
		19'b0011010010011111001: color_data = Z;
		19'b0011010010011111010: color_data = Z;
		19'b0011010010011111011: color_data = Z;
		19'b0011010010011111100: color_data = Z;
		19'b0011010010011111101: color_data = Z;
		19'b0011010010011111110: color_data = Z;
		19'b0011010010011111111: color_data = Z;
		19'b0011010010100000000: color_data = Z;
		19'b0011010010100000001: color_data = Z;
		19'b0011010010100000010: color_data = Z;
		19'b0011010010100000011: color_data = Z;
		19'b0011010010100000100: color_data = Z;
		19'b0011010010100000101: color_data = Z;
		19'b0011010010100000110: color_data = Z;
		19'b0011010010100000111: color_data = Z;
		19'b0011010010100001000: color_data = Z;
		19'b0011010010100001001: color_data = Z;
		19'b0011010010100001010: color_data = Z;
		19'b0011010010100001011: color_data = Z;
		19'b0011010010100001100: color_data = Z;
		19'b0011010010100001101: color_data = Z;
		19'b0011010010100001110: color_data = Z;
		19'b0011010010100001111: color_data = Z;
		19'b0011010010100010000: color_data = Z;
		19'b0011010010100010001: color_data = Z;
		19'b0011010010100010010: color_data = Z;
		19'b0011010010100010011: color_data = Z;
		19'b0011010010100010100: color_data = Z;
		19'b0011010010100010101: color_data = Z;
		19'b0011010010100010110: color_data = Z;
		19'b0011010010100010111: color_data = Z;
		19'b0011010010100011000: color_data = Z;
		19'b0011010010100011001: color_data = Z;
		19'b0011010010100011010: color_data = Z;
		19'b0011010010100011011: color_data = Z;
		19'b0011010010100011100: color_data = Z;
		19'b0011010010100011101: color_data = Z;
		19'b0011010010100011110: color_data = Z;
		19'b0011010010100011111: color_data = Z;
		19'b0011010010100100000: color_data = Z;
		19'b0011010010100100001: color_data = Z;
		19'b0011010010100100010: color_data = Z;
		19'b0011010010100100011: color_data = Z;
		19'b0011010010100100100: color_data = Z;
		19'b0011010010100100101: color_data = Z;
		19'b0011010010100100110: color_data = Z;
		19'b0011010010100100111: color_data = Z;
		19'b0011010010100101000: color_data = Z;
		19'b0011010010100101001: color_data = Z;
		19'b0011010010100101010: color_data = Z;
		19'b0011010010100101011: color_data = Z;
		19'b0011010010100101100: color_data = Z;
		19'b0011010010100101101: color_data = Z;
		19'b0011010010100101110: color_data = Z;
		19'b0011010010100101111: color_data = Z;
		19'b0011010010100110000: color_data = Z;
		19'b0011010010100110001: color_data = Z;
		19'b0011010010100110010: color_data = Z;
		19'b0011010010100110011: color_data = Z;
		19'b0011010010100110100: color_data = Z;
		19'b0011010010100110101: color_data = Z;
		19'b0011010010100110110: color_data = Z;
		19'b0011010010100110111: color_data = Z;
		19'b0011010010100111000: color_data = Z;
		19'b0011010010100111001: color_data = Z;
		19'b0011010010100111010: color_data = Z;
		19'b0011010010100111011: color_data = Z;
		19'b0011010010100111100: color_data = Z;
		19'b0011010010100111101: color_data = Z;
		19'b0011010010100111110: color_data = Z;
		19'b0011010010100111111: color_data = Z;
		19'b0011010010101000000: color_data = Z;
		19'b0011010010101000001: color_data = Z;
		19'b0011010010101000010: color_data = Z;
		19'b0011010010101000011: color_data = Z;
		19'b0011010010101000100: color_data = Z;
		19'b0011010010101000101: color_data = Z;
		19'b0011010010101000110: color_data = Z;
		19'b0011010010101000111: color_data = Z;
		19'b0011010010101001000: color_data = Z;
		19'b0011010010101001001: color_data = Z;
		19'b0011010010101001010: color_data = Z;
		19'b0011010010101001011: color_data = Z;
		19'b0011010010101001100: color_data = Z;
		19'b0011010010101001101: color_data = Z;
		19'b0011010010101001110: color_data = Z;
		19'b0011010010101001111: color_data = Z;
		19'b0011010010101010000: color_data = Z;
		19'b0011010010101010001: color_data = Z;
		19'b0011010010101010010: color_data = Z;
		19'b0011010010101010011: color_data = Z;
		19'b0011010010101010100: color_data = Z;
		19'b0011010010101010101: color_data = Z;
		19'b0011010010101010110: color_data = Z;
		19'b0011010010101010111: color_data = Z;
		19'b0011010010101011000: color_data = Z;
		19'b0011010010101011001: color_data = Z;
		19'b0011010010101011010: color_data = Z;
		19'b0011010010101011011: color_data = Z;
		19'b0011010010101011100: color_data = Z;
		19'b0011010010101011101: color_data = Z;
		19'b0011010010101011110: color_data = Z;
		19'b0011010010101011111: color_data = Z;
		19'b0011010010101100000: color_data = Z;
		19'b0011010010101100001: color_data = Z;
		19'b0011010010101100010: color_data = Z;
		19'b0011010010101100011: color_data = Z;
		19'b0011010010101100100: color_data = Z;
		19'b0011010010101100101: color_data = Z;
		19'b0011010010101100110: color_data = Z;
		19'b0011010010101100111: color_data = Z;
		19'b0011010010101101000: color_data = Z;
		19'b0011010010101101001: color_data = Z;
		19'b0011010010101101010: color_data = Z;
		19'b0011010010101101011: color_data = Z;
		19'b0011010010101101100: color_data = Z;
		19'b0011010010101101101: color_data = Z;
		19'b0011010010101101110: color_data = Z;
		19'b0011010010101101111: color_data = Z;
		19'b0011010010101110000: color_data = Z;
		19'b0011010010101110001: color_data = Z;
		19'b0011010010101110010: color_data = Z;
		19'b0011010010101110011: color_data = Z;
		19'b0011010010101110100: color_data = Z;
		19'b0011010010101110101: color_data = Z;
		19'b0011010010101110110: color_data = Z;
		19'b0011010010101110111: color_data = Z;
		19'b0011010010101111000: color_data = Z;
		19'b0011010010101111001: color_data = Z;
		19'b0011010010101111010: color_data = Z;
		19'b0011010010101111011: color_data = Z;
		19'b0011010010101111100: color_data = Z;
		19'b0011010010101111101: color_data = Z;
		19'b0011010010101111110: color_data = Z;
		19'b0011010010101111111: color_data = Z;
		19'b0011010010110000000: color_data = Z;
		19'b0011010010110000001: color_data = Z;
		19'b0011010010110000010: color_data = Z;
		19'b0011010010110000011: color_data = Z;
		19'b0011010010110000100: color_data = Z;
		19'b0011010010110000101: color_data = Z;
		19'b0011010010110000110: color_data = Z;
		19'b0011010010110000111: color_data = Z;
		19'b0011010010110001000: color_data = Z;
		19'b0011010010110001001: color_data = Z;
		19'b0011010010110001010: color_data = Z;
		19'b0011010010110001011: color_data = Z;
		19'b0011010010110001100: color_data = Z;
		19'b0011010010110001101: color_data = Z;
		19'b0011010010110001110: color_data = Z;
		19'b0011010010110001111: color_data = Z;
		19'b0011010010110010000: color_data = Z;
		19'b0011010010110010001: color_data = Z;
		19'b0011010010110010010: color_data = Z;
		19'b0011010010110010011: color_data = Z;
		19'b0011010010110010100: color_data = Z;
		19'b0011010010110010101: color_data = Z;
		19'b0011010010110010110: color_data = Z;
		19'b0011010010110010111: color_data = Z;
		19'b0011010010110011000: color_data = Z;
		19'b0011010010110011001: color_data = Z;
		19'b0011010010110011100: color_data = Z;
		19'b0011010010110011101: color_data = Z;
		19'b0011010010110110101: color_data = Z;
		19'b0011010010110110110: color_data = Z;
		19'b0011010010110110111: color_data = Z;
		19'b0011010010110111000: color_data = Z;
		19'b0011010010110111001: color_data = Z;
		19'b0011010010111010011: color_data = Z;
		19'b0011010100010110000: color_data = Z;
		19'b0011010100010110001: color_data = Z;
		19'b0011010100010110010: color_data = Z;
		19'b0011010100010110011: color_data = Z;
		19'b0011010100010110100: color_data = Z;
		19'b0011010100010110101: color_data = Z;
		19'b0011010100010110110: color_data = Z;
		19'b0011010100010110111: color_data = Z;
		19'b0011010100010111000: color_data = Z;
		19'b0011010100010111001: color_data = Z;
		19'b0011010100010111010: color_data = Z;
		19'b0011010100010111011: color_data = Z;
		19'b0011010100010111100: color_data = Z;
		19'b0011010100010111101: color_data = Z;
		19'b0011010100010111110: color_data = Z;
		19'b0011010100010111111: color_data = Z;
		19'b0011010100011000000: color_data = Z;
		19'b0011010100011000001: color_data = Z;
		19'b0011010100011000010: color_data = Z;
		19'b0011010100011000011: color_data = Z;
		19'b0011010100011000100: color_data = Z;
		19'b0011010100011000101: color_data = Z;
		19'b0011010100011000110: color_data = Z;
		19'b0011010100011000111: color_data = Z;
		19'b0011010100011001000: color_data = Z;
		19'b0011010100011001001: color_data = Z;
		19'b0011010100011001010: color_data = Z;
		19'b0011010100011001011: color_data = Z;
		19'b0011010100011001100: color_data = Z;
		19'b0011010100011001101: color_data = Z;
		19'b0011010100011001110: color_data = Z;
		19'b0011010100011001111: color_data = Z;
		19'b0011010100011010000: color_data = Z;
		19'b0011010100011010001: color_data = Z;
		19'b0011010100011010010: color_data = Z;
		19'b0011010100011010011: color_data = Z;
		19'b0011010100011010100: color_data = Z;
		19'b0011010100011010101: color_data = Z;
		19'b0011010100011010110: color_data = Z;
		19'b0011010100011010111: color_data = Z;
		19'b0011010100011011000: color_data = Z;
		19'b0011010100011011001: color_data = Z;
		19'b0011010100011011010: color_data = Z;
		19'b0011010100011011011: color_data = Z;
		19'b0011010100011011100: color_data = Z;
		19'b0011010100011011101: color_data = Z;
		19'b0011010100011011110: color_data = Z;
		19'b0011010100011011111: color_data = Z;
		19'b0011010100011100000: color_data = Z;
		19'b0011010100011100001: color_data = Z;
		19'b0011010100011100010: color_data = Z;
		19'b0011010100011100011: color_data = Z;
		19'b0011010100011100100: color_data = Z;
		19'b0011010100011100101: color_data = Z;
		19'b0011010100011100110: color_data = Z;
		19'b0011010100011100111: color_data = Z;
		19'b0011010100011101000: color_data = Z;
		19'b0011010100011101001: color_data = Z;
		19'b0011010100011101010: color_data = Z;
		19'b0011010100011101011: color_data = Z;
		19'b0011010100011101100: color_data = Z;
		19'b0011010100011101101: color_data = Z;
		19'b0011010100011101110: color_data = Z;
		19'b0011010100011101111: color_data = Z;
		19'b0011010100011110000: color_data = Z;
		19'b0011010100011110001: color_data = Z;
		19'b0011010100011110010: color_data = Z;
		19'b0011010100011110011: color_data = Z;
		19'b0011010100011110100: color_data = Z;
		19'b0011010100011110101: color_data = Z;
		19'b0011010100011110110: color_data = Z;
		19'b0011010100011110111: color_data = Z;
		19'b0011010100011111000: color_data = Z;
		19'b0011010100011111001: color_data = Z;
		19'b0011010100011111010: color_data = Z;
		19'b0011010100011111011: color_data = Z;
		19'b0011010100011111100: color_data = Z;
		19'b0011010100011111101: color_data = Z;
		19'b0011010100011111110: color_data = Z;
		19'b0011010100011111111: color_data = Z;
		19'b0011010100100000000: color_data = Z;
		19'b0011010100100000001: color_data = Z;
		19'b0011010100100000010: color_data = Z;
		19'b0011010100100000011: color_data = Z;
		19'b0011010100100000100: color_data = Z;
		19'b0011010100100000101: color_data = Z;
		19'b0011010100100000110: color_data = Z;
		19'b0011010100100000111: color_data = Z;
		19'b0011010100100001000: color_data = Z;
		19'b0011010100100001001: color_data = Z;
		19'b0011010100100001010: color_data = Z;
		19'b0011010100100001011: color_data = Z;
		19'b0011010100100001100: color_data = Z;
		19'b0011010100100001101: color_data = Z;
		19'b0011010100100001110: color_data = Z;
		19'b0011010100100001111: color_data = Z;
		19'b0011010100100010000: color_data = Z;
		19'b0011010100100010001: color_data = Z;
		19'b0011010100100010010: color_data = Z;
		19'b0011010100100010011: color_data = Z;
		19'b0011010100100010100: color_data = Z;
		19'b0011010100100010101: color_data = Z;
		19'b0011010100100010110: color_data = Z;
		19'b0011010100100010111: color_data = Z;
		19'b0011010100100011000: color_data = Z;
		19'b0011010100100011001: color_data = Z;
		19'b0011010100100011010: color_data = Z;
		19'b0011010100100011011: color_data = Z;
		19'b0011010100100011100: color_data = Z;
		19'b0011010100100011101: color_data = Z;
		19'b0011010100100011110: color_data = Z;
		19'b0011010100100011111: color_data = Z;
		19'b0011010100100100000: color_data = Z;
		19'b0011010100100100001: color_data = Z;
		19'b0011010100100100010: color_data = Z;
		19'b0011010100100100011: color_data = Z;
		19'b0011010100100100100: color_data = Z;
		19'b0011010100100100101: color_data = Z;
		19'b0011010100100100110: color_data = Z;
		19'b0011010100100100111: color_data = Z;
		19'b0011010100100101000: color_data = Z;
		19'b0011010100100101001: color_data = Z;
		19'b0011010100100101010: color_data = Z;
		19'b0011010100100101011: color_data = Z;
		19'b0011010100100101100: color_data = Z;
		19'b0011010100100101101: color_data = Z;
		19'b0011010100100101110: color_data = Z;
		19'b0011010100100101111: color_data = Z;
		19'b0011010100100110000: color_data = Z;
		19'b0011010100100110001: color_data = Z;
		19'b0011010100100110010: color_data = Z;
		19'b0011010100100110011: color_data = Z;
		19'b0011010100100110100: color_data = Z;
		19'b0011010100100110101: color_data = Z;
		19'b0011010100100110110: color_data = Z;
		19'b0011010100100110111: color_data = Z;
		19'b0011010100100111000: color_data = Z;
		19'b0011010100100111001: color_data = Z;
		19'b0011010100100111010: color_data = Z;
		19'b0011010100100111011: color_data = Z;
		19'b0011010100100111100: color_data = Z;
		19'b0011010100100111101: color_data = Z;
		19'b0011010100100111110: color_data = Z;
		19'b0011010100100111111: color_data = Z;
		19'b0011010100101000000: color_data = Z;
		19'b0011010100101000001: color_data = Z;
		19'b0011010100101000010: color_data = Z;
		19'b0011010100101000011: color_data = Z;
		19'b0011010100101000100: color_data = Z;
		19'b0011010100101000101: color_data = Z;
		19'b0011010100101000110: color_data = Z;
		19'b0011010100101000111: color_data = Z;
		19'b0011010100101001000: color_data = Z;
		19'b0011010100101001001: color_data = Z;
		19'b0011010100101001010: color_data = Z;
		19'b0011010100101001011: color_data = Z;
		19'b0011010100101001100: color_data = Z;
		19'b0011010100101001101: color_data = Z;
		19'b0011010100101001110: color_data = Z;
		19'b0011010100101001111: color_data = Z;
		19'b0011010100101010000: color_data = Z;
		19'b0011010100101010001: color_data = Z;
		19'b0011010100101010010: color_data = Z;
		19'b0011010100101010011: color_data = Z;
		19'b0011010100101010100: color_data = Z;
		19'b0011010100101010101: color_data = Z;
		19'b0011010100101010110: color_data = Z;
		19'b0011010100101010111: color_data = Z;
		19'b0011010100101011000: color_data = Z;
		19'b0011010100101011001: color_data = Z;
		19'b0011010100101011010: color_data = Z;
		19'b0011010100101011011: color_data = Z;
		19'b0011010100101011100: color_data = Z;
		19'b0011010100101011101: color_data = Z;
		19'b0011010100101011110: color_data = Z;
		19'b0011010100101011111: color_data = Z;
		19'b0011010100101100000: color_data = Z;
		19'b0011010100101100001: color_data = Z;
		19'b0011010100101100010: color_data = Z;
		19'b0011010100101100011: color_data = Z;
		19'b0011010100101100100: color_data = Z;
		19'b0011010100101100101: color_data = Z;
		19'b0011010100101100110: color_data = Z;
		19'b0011010100101100111: color_data = Z;
		19'b0011010100101101000: color_data = Z;
		19'b0011010100101101001: color_data = Z;
		19'b0011010100101101010: color_data = Z;
		19'b0011010100101101011: color_data = Z;
		19'b0011010100101101100: color_data = Z;
		19'b0011010100101101101: color_data = Z;
		19'b0011010100101101110: color_data = Z;
		19'b0011010100101101111: color_data = Z;
		19'b0011010100101110000: color_data = Z;
		19'b0011010100101110001: color_data = Z;
		19'b0011010100101110010: color_data = Z;
		19'b0011010100101110011: color_data = Z;
		19'b0011010100101110100: color_data = Z;
		19'b0011010100101110101: color_data = Z;
		19'b0011010100101110110: color_data = Z;
		19'b0011010100101110111: color_data = Z;
		19'b0011010100101111000: color_data = Z;
		19'b0011010100101111001: color_data = Z;
		19'b0011010100101111010: color_data = Z;
		19'b0011010100101111011: color_data = Z;
		19'b0011010100101111100: color_data = Z;
		19'b0011010100101111101: color_data = Z;
		19'b0011010100101111110: color_data = Z;
		19'b0011010100101111111: color_data = Z;
		19'b0011010100110000000: color_data = Z;
		19'b0011010100110000001: color_data = Z;
		19'b0011010100110000010: color_data = Z;
		19'b0011010100110000011: color_data = Z;
		19'b0011010100110000100: color_data = Z;
		19'b0011010100110000101: color_data = Z;
		19'b0011010100110000110: color_data = Z;
		19'b0011010100110000111: color_data = Z;
		19'b0011010100110001000: color_data = Z;
		19'b0011010100110001001: color_data = Z;
		19'b0011010100110001010: color_data = Z;
		19'b0011010100110001011: color_data = Z;
		19'b0011010100110001100: color_data = Z;
		19'b0011010100110001101: color_data = Z;
		19'b0011010100110001110: color_data = Z;
		19'b0011010100110001111: color_data = Z;
		19'b0011010100110010000: color_data = Z;
		19'b0011010100110010001: color_data = Z;
		19'b0011010100110010010: color_data = Z;
		19'b0011010100110010011: color_data = Z;
		19'b0011010100110010100: color_data = Z;
		19'b0011010100110010101: color_data = Z;
		19'b0011010100110010110: color_data = Z;
		19'b0011010100110010111: color_data = Z;
		19'b0011010100110011000: color_data = Z;
		19'b0011010100110110110: color_data = Z;
		19'b0011010100110110111: color_data = Z;
		19'b0011010100110111000: color_data = Z;
		19'b0011010100110111001: color_data = Z;
		19'b0011010100111001100: color_data = Z;
		19'b0011010110010101111: color_data = Z;
		19'b0011010110010110000: color_data = Z;
		19'b0011010110010110001: color_data = Z;
		19'b0011010110010110010: color_data = Z;
		19'b0011010110010110011: color_data = Z;
		19'b0011010110010110100: color_data = Z;
		19'b0011010110010110101: color_data = Z;
		19'b0011010110010110110: color_data = Z;
		19'b0011010110010110111: color_data = Z;
		19'b0011010110010111000: color_data = Z;
		19'b0011010110010111001: color_data = Z;
		19'b0011010110010111010: color_data = Z;
		19'b0011010110010111011: color_data = Z;
		19'b0011010110010111100: color_data = Z;
		19'b0011010110010111101: color_data = Z;
		19'b0011010110010111110: color_data = Z;
		19'b0011010110010111111: color_data = Z;
		19'b0011010110011000000: color_data = Z;
		19'b0011010110011000001: color_data = Z;
		19'b0011010110011000010: color_data = Z;
		19'b0011010110011000011: color_data = Z;
		19'b0011010110011000100: color_data = Z;
		19'b0011010110011000101: color_data = Z;
		19'b0011010110011000110: color_data = Z;
		19'b0011010110011000111: color_data = Z;
		19'b0011010110011001000: color_data = Z;
		19'b0011010110011001001: color_data = Z;
		19'b0011010110011001010: color_data = Z;
		19'b0011010110011001011: color_data = Z;
		19'b0011010110011001100: color_data = Z;
		19'b0011010110011001101: color_data = Z;
		19'b0011010110011001110: color_data = Z;
		19'b0011010110011001111: color_data = Z;
		19'b0011010110011010000: color_data = Z;
		19'b0011010110011010001: color_data = Z;
		19'b0011010110011010010: color_data = Z;
		19'b0011010110011010011: color_data = Z;
		19'b0011010110011010100: color_data = Z;
		19'b0011010110011010101: color_data = Z;
		19'b0011010110011010110: color_data = Z;
		19'b0011010110011010111: color_data = Z;
		19'b0011010110011011000: color_data = Z;
		19'b0011010110011011001: color_data = Z;
		19'b0011010110011011010: color_data = Z;
		19'b0011010110011011011: color_data = Z;
		19'b0011010110011011100: color_data = Z;
		19'b0011010110011011101: color_data = Z;
		19'b0011010110011011110: color_data = Z;
		19'b0011010110011011111: color_data = Z;
		19'b0011010110011100000: color_data = Z;
		19'b0011010110011100001: color_data = Z;
		19'b0011010110011100010: color_data = Z;
		19'b0011010110011100011: color_data = Z;
		19'b0011010110011100100: color_data = Z;
		19'b0011010110011100101: color_data = Z;
		19'b0011010110011100110: color_data = Z;
		19'b0011010110011100111: color_data = Z;
		19'b0011010110011101000: color_data = Z;
		19'b0011010110011101001: color_data = Z;
		19'b0011010110011101010: color_data = Z;
		19'b0011010110011101011: color_data = Z;
		19'b0011010110011101100: color_data = Z;
		19'b0011010110011101101: color_data = Z;
		19'b0011010110011101110: color_data = Z;
		19'b0011010110011101111: color_data = Z;
		19'b0011010110011110000: color_data = Z;
		19'b0011010110011110001: color_data = Z;
		19'b0011010110011110010: color_data = Z;
		19'b0011010110011110011: color_data = Z;
		19'b0011010110011110100: color_data = Z;
		19'b0011010110011110101: color_data = Z;
		19'b0011010110011110110: color_data = Z;
		19'b0011010110011110111: color_data = Z;
		19'b0011010110011111000: color_data = Z;
		19'b0011010110011111001: color_data = Z;
		19'b0011010110011111010: color_data = Z;
		19'b0011010110011111011: color_data = Z;
		19'b0011010110011111100: color_data = Z;
		19'b0011010110011111101: color_data = Z;
		19'b0011010110011111110: color_data = Z;
		19'b0011010110011111111: color_data = Z;
		19'b0011010110100000000: color_data = Z;
		19'b0011010110100000001: color_data = Z;
		19'b0011010110100000010: color_data = Z;
		19'b0011010110100000011: color_data = Z;
		19'b0011010110100000100: color_data = Z;
		19'b0011010110100000101: color_data = Z;
		19'b0011010110100000110: color_data = Z;
		19'b0011010110100000111: color_data = Z;
		19'b0011010110100001000: color_data = Z;
		19'b0011010110100001001: color_data = Z;
		19'b0011010110100001010: color_data = Z;
		19'b0011010110100001011: color_data = Z;
		19'b0011010110100001100: color_data = Z;
		19'b0011010110100001101: color_data = Z;
		19'b0011010110100001110: color_data = Z;
		19'b0011010110100001111: color_data = Z;
		19'b0011010110100010000: color_data = Z;
		19'b0011010110100010001: color_data = Z;
		19'b0011010110100010010: color_data = Z;
		19'b0011010110100010011: color_data = Z;
		19'b0011010110100010100: color_data = Z;
		19'b0011010110100010101: color_data = Z;
		19'b0011010110100010110: color_data = Z;
		19'b0011010110100010111: color_data = Z;
		19'b0011010110100011000: color_data = Z;
		19'b0011010110100011001: color_data = Z;
		19'b0011010110100011010: color_data = Z;
		19'b0011010110100011011: color_data = Z;
		19'b0011010110100011100: color_data = Z;
		19'b0011010110100011101: color_data = Z;
		19'b0011010110100011110: color_data = Z;
		19'b0011010110100011111: color_data = Z;
		19'b0011010110100100000: color_data = Z;
		19'b0011010110100100001: color_data = Z;
		19'b0011010110100100010: color_data = Z;
		19'b0011010110100100011: color_data = Z;
		19'b0011010110100100100: color_data = Z;
		19'b0011010110100100101: color_data = Z;
		19'b0011010110100100110: color_data = Z;
		19'b0011010110100100111: color_data = Z;
		19'b0011010110100101000: color_data = Z;
		19'b0011010110100101001: color_data = Z;
		19'b0011010110100101010: color_data = Z;
		19'b0011010110100101011: color_data = Z;
		19'b0011010110100101100: color_data = Z;
		19'b0011010110100101101: color_data = Z;
		19'b0011010110100101110: color_data = Z;
		19'b0011010110100101111: color_data = Z;
		19'b0011010110100110000: color_data = Z;
		19'b0011010110100110001: color_data = Z;
		19'b0011010110100110010: color_data = Z;
		19'b0011010110100110011: color_data = Z;
		19'b0011010110100110100: color_data = Z;
		19'b0011010110100110101: color_data = Z;
		19'b0011010110100110110: color_data = Z;
		19'b0011010110100110111: color_data = Z;
		19'b0011010110100111000: color_data = Z;
		19'b0011010110100111001: color_data = Z;
		19'b0011010110100111010: color_data = Z;
		19'b0011010110100111011: color_data = Z;
		19'b0011010110100111100: color_data = Z;
		19'b0011010110100111101: color_data = Z;
		19'b0011010110100111110: color_data = Z;
		19'b0011010110100111111: color_data = Z;
		19'b0011010110101000000: color_data = Z;
		19'b0011010110101000001: color_data = Z;
		19'b0011010110101000010: color_data = Z;
		19'b0011010110101000011: color_data = Z;
		19'b0011010110101000100: color_data = Z;
		19'b0011010110101000101: color_data = Z;
		19'b0011010110101000110: color_data = Z;
		19'b0011010110101000111: color_data = Z;
		19'b0011010110101001000: color_data = Z;
		19'b0011010110101001001: color_data = Z;
		19'b0011010110101001010: color_data = Z;
		19'b0011010110101001011: color_data = Z;
		19'b0011010110101001100: color_data = Z;
		19'b0011010110101001101: color_data = Z;
		19'b0011010110101001110: color_data = Z;
		19'b0011010110101001111: color_data = Z;
		19'b0011010110101010000: color_data = Z;
		19'b0011010110101010001: color_data = Z;
		19'b0011010110101010010: color_data = Z;
		19'b0011010110101010011: color_data = Z;
		19'b0011010110101010100: color_data = Z;
		19'b0011010110101010101: color_data = Z;
		19'b0011010110101010110: color_data = Z;
		19'b0011010110101010111: color_data = Z;
		19'b0011010110101011000: color_data = Z;
		19'b0011010110101011001: color_data = Z;
		19'b0011010110101011010: color_data = Z;
		19'b0011010110101011011: color_data = Z;
		19'b0011010110101011100: color_data = Z;
		19'b0011010110101011101: color_data = Z;
		19'b0011010110101011110: color_data = Z;
		19'b0011010110101011111: color_data = Z;
		19'b0011010110101100000: color_data = Z;
		19'b0011010110101100001: color_data = Z;
		19'b0011010110101100010: color_data = Z;
		19'b0011010110101100011: color_data = Z;
		19'b0011010110101100100: color_data = Z;
		19'b0011010110101100101: color_data = Z;
		19'b0011010110101100110: color_data = Z;
		19'b0011010110101100111: color_data = Z;
		19'b0011010110101101000: color_data = Z;
		19'b0011010110101101001: color_data = Z;
		19'b0011010110101101010: color_data = Z;
		19'b0011010110101101011: color_data = Z;
		19'b0011010110101101100: color_data = Z;
		19'b0011010110101101101: color_data = Z;
		19'b0011010110101101110: color_data = Z;
		19'b0011010110101101111: color_data = Z;
		19'b0011010110101110000: color_data = Z;
		19'b0011010110101110001: color_data = Z;
		19'b0011010110101110010: color_data = Z;
		19'b0011010110101110011: color_data = Z;
		19'b0011010110101110100: color_data = Z;
		19'b0011010110101110101: color_data = Z;
		19'b0011010110101110110: color_data = Z;
		19'b0011010110101110111: color_data = Z;
		19'b0011010110101111000: color_data = Z;
		19'b0011010110101111001: color_data = Z;
		19'b0011010110101111010: color_data = Z;
		19'b0011010110101111011: color_data = Z;
		19'b0011010110101111100: color_data = Z;
		19'b0011010110101111101: color_data = Z;
		19'b0011010110101111110: color_data = Z;
		19'b0011010110101111111: color_data = Z;
		19'b0011010110110000000: color_data = Z;
		19'b0011010110110000001: color_data = Z;
		19'b0011010110110000010: color_data = Z;
		19'b0011010110110000011: color_data = Z;
		19'b0011010110110000100: color_data = Z;
		19'b0011010110110000101: color_data = Z;
		19'b0011010110110000110: color_data = Z;
		19'b0011010110110000111: color_data = Z;
		19'b0011010110110001000: color_data = Z;
		19'b0011010110110001001: color_data = Z;
		19'b0011010110110001010: color_data = Z;
		19'b0011010110110001011: color_data = Z;
		19'b0011010110110001100: color_data = Z;
		19'b0011010110110001101: color_data = Z;
		19'b0011010110110001110: color_data = Z;
		19'b0011010110110001111: color_data = Z;
		19'b0011010110110010000: color_data = Z;
		19'b0011010110110010001: color_data = Z;
		19'b0011010110110010010: color_data = Z;
		19'b0011010110110010011: color_data = Z;
		19'b0011010110110010100: color_data = Z;
		19'b0011010110110010101: color_data = Z;
		19'b0011010110110010110: color_data = Z;
		19'b0011010110110010111: color_data = Z;
		19'b0011010110110111000: color_data = Z;
		19'b0011010110110111001: color_data = Z;
		19'b0011010110110111010: color_data = Z;
		19'b0011010110111001100: color_data = Z;
		19'b0011010110111001101: color_data = Z;
		19'b0011011000010101111: color_data = Z;
		19'b0011011000010110000: color_data = Z;
		19'b0011011000010110001: color_data = Z;
		19'b0011011000010110010: color_data = Z;
		19'b0011011000010110011: color_data = Z;
		19'b0011011000010110100: color_data = Z;
		19'b0011011000010110101: color_data = Z;
		19'b0011011000010110110: color_data = Z;
		19'b0011011000010110111: color_data = Z;
		19'b0011011000010111000: color_data = Z;
		19'b0011011000010111001: color_data = Z;
		19'b0011011000010111010: color_data = Z;
		19'b0011011000010111011: color_data = Z;
		19'b0011011000010111100: color_data = Z;
		19'b0011011000010111101: color_data = Z;
		19'b0011011000010111110: color_data = Z;
		19'b0011011000010111111: color_data = Z;
		19'b0011011000011000000: color_data = Z;
		19'b0011011000011000001: color_data = Z;
		19'b0011011000011000010: color_data = Z;
		19'b0011011000011000011: color_data = Z;
		19'b0011011000011000100: color_data = Z;
		19'b0011011000011000101: color_data = Z;
		19'b0011011000011000110: color_data = Z;
		19'b0011011000011000111: color_data = Z;
		19'b0011011000011001000: color_data = Z;
		19'b0011011000011001001: color_data = Z;
		19'b0011011000011001010: color_data = Z;
		19'b0011011000011001011: color_data = Z;
		19'b0011011000011001100: color_data = Z;
		19'b0011011000011001101: color_data = Z;
		19'b0011011000011001110: color_data = Z;
		19'b0011011000011001111: color_data = Z;
		19'b0011011000011010000: color_data = Z;
		19'b0011011000011010001: color_data = Z;
		19'b0011011000011010010: color_data = Z;
		19'b0011011000011010011: color_data = Z;
		19'b0011011000011010100: color_data = Z;
		19'b0011011000011010101: color_data = Z;
		19'b0011011000011010110: color_data = Z;
		19'b0011011000011010111: color_data = Z;
		19'b0011011000011011000: color_data = Z;
		19'b0011011000011011001: color_data = Z;
		19'b0011011000011011010: color_data = Z;
		19'b0011011000011011011: color_data = Z;
		19'b0011011000011011100: color_data = Z;
		19'b0011011000011011101: color_data = Z;
		19'b0011011000011011110: color_data = Z;
		19'b0011011000011011111: color_data = Z;
		19'b0011011000011100000: color_data = Z;
		19'b0011011000011100001: color_data = Z;
		19'b0011011000011100010: color_data = Z;
		19'b0011011000011100011: color_data = Z;
		19'b0011011000011100100: color_data = Z;
		19'b0011011000011100101: color_data = Z;
		19'b0011011000011100110: color_data = Z;
		19'b0011011000011100111: color_data = Z;
		19'b0011011000011101000: color_data = Z;
		19'b0011011000011101001: color_data = Z;
		19'b0011011000011101010: color_data = Z;
		19'b0011011000011101011: color_data = Z;
		19'b0011011000011101100: color_data = Z;
		19'b0011011000011101101: color_data = Z;
		19'b0011011000011101110: color_data = Z;
		19'b0011011000011101111: color_data = Z;
		19'b0011011000011110000: color_data = Z;
		19'b0011011000011110001: color_data = Z;
		19'b0011011000011110010: color_data = Z;
		19'b0011011000011110011: color_data = Z;
		19'b0011011000011110100: color_data = Z;
		19'b0011011000011110101: color_data = Z;
		19'b0011011000011110110: color_data = Z;
		19'b0011011000011110111: color_data = Z;
		19'b0011011000011111000: color_data = Z;
		19'b0011011000011111001: color_data = Z;
		19'b0011011000011111010: color_data = Z;
		19'b0011011000011111011: color_data = Z;
		19'b0011011000011111100: color_data = Z;
		19'b0011011000011111101: color_data = Z;
		19'b0011011000011111110: color_data = Z;
		19'b0011011000011111111: color_data = Z;
		19'b0011011000100000000: color_data = Z;
		19'b0011011000100000001: color_data = Z;
		19'b0011011000100000010: color_data = Z;
		19'b0011011000100000011: color_data = Z;
		19'b0011011000100000100: color_data = Z;
		19'b0011011000100000101: color_data = Z;
		19'b0011011000100000110: color_data = Z;
		19'b0011011000100000111: color_data = Z;
		19'b0011011000100001000: color_data = Z;
		19'b0011011000100001001: color_data = Z;
		19'b0011011000100001010: color_data = Z;
		19'b0011011000100001011: color_data = Z;
		19'b0011011000100001100: color_data = Z;
		19'b0011011000100001101: color_data = Z;
		19'b0011011000100001110: color_data = Z;
		19'b0011011000100001111: color_data = Z;
		19'b0011011000100010000: color_data = Z;
		19'b0011011000100010001: color_data = Z;
		19'b0011011000100010010: color_data = Z;
		19'b0011011000100010011: color_data = Z;
		19'b0011011000100010100: color_data = Z;
		19'b0011011000100010101: color_data = Z;
		19'b0011011000100010110: color_data = Z;
		19'b0011011000100010111: color_data = Z;
		19'b0011011000100011000: color_data = Z;
		19'b0011011000100011001: color_data = Z;
		19'b0011011000100011010: color_data = Z;
		19'b0011011000100011011: color_data = Z;
		19'b0011011000100011100: color_data = Z;
		19'b0011011000100011101: color_data = Z;
		19'b0011011000100011110: color_data = Z;
		19'b0011011000100011111: color_data = Z;
		19'b0011011000100100000: color_data = Z;
		19'b0011011000100100001: color_data = Z;
		19'b0011011000100100010: color_data = Z;
		19'b0011011000100100011: color_data = Z;
		19'b0011011000100100100: color_data = Z;
		19'b0011011000100100101: color_data = Z;
		19'b0011011000100100110: color_data = Z;
		19'b0011011000100100111: color_data = Z;
		19'b0011011000100101000: color_data = Z;
		19'b0011011000100101001: color_data = Z;
		19'b0011011000100101010: color_data = Z;
		19'b0011011000100101011: color_data = Z;
		19'b0011011000100101100: color_data = Z;
		19'b0011011000100101101: color_data = Z;
		19'b0011011000100101110: color_data = Z;
		19'b0011011000100101111: color_data = Z;
		19'b0011011000100110000: color_data = Z;
		19'b0011011000100110001: color_data = Z;
		19'b0011011000100110010: color_data = Z;
		19'b0011011000100110011: color_data = Z;
		19'b0011011000100110100: color_data = Z;
		19'b0011011000100110101: color_data = Z;
		19'b0011011000100110110: color_data = Z;
		19'b0011011000100110111: color_data = Z;
		19'b0011011000100111000: color_data = Z;
		19'b0011011000100111001: color_data = Z;
		19'b0011011000100111010: color_data = Z;
		19'b0011011000100111011: color_data = Z;
		19'b0011011000100111100: color_data = Z;
		19'b0011011000100111101: color_data = Z;
		19'b0011011000100111110: color_data = Z;
		19'b0011011000100111111: color_data = Z;
		19'b0011011000101000000: color_data = Z;
		19'b0011011000101000001: color_data = Z;
		19'b0011011000101000010: color_data = Z;
		19'b0011011000101000011: color_data = Z;
		19'b0011011000101000100: color_data = Z;
		19'b0011011000101000101: color_data = Z;
		19'b0011011000101000110: color_data = Z;
		19'b0011011000101000111: color_data = Z;
		19'b0011011000101001000: color_data = Z;
		19'b0011011000101001001: color_data = Z;
		19'b0011011000101001010: color_data = Z;
		19'b0011011000101001011: color_data = Z;
		19'b0011011000101001100: color_data = Z;
		19'b0011011000101001101: color_data = Z;
		19'b0011011000101001110: color_data = Z;
		19'b0011011000101001111: color_data = Z;
		19'b0011011000101010000: color_data = Z;
		19'b0011011000101010001: color_data = Z;
		19'b0011011000101010010: color_data = Z;
		19'b0011011000101010011: color_data = Z;
		19'b0011011000101010100: color_data = Z;
		19'b0011011000101010101: color_data = Z;
		19'b0011011000101010110: color_data = Z;
		19'b0011011000101010111: color_data = Z;
		19'b0011011000101011000: color_data = Z;
		19'b0011011000101011001: color_data = Z;
		19'b0011011000101011010: color_data = Z;
		19'b0011011000101011011: color_data = Z;
		19'b0011011000101011100: color_data = Z;
		19'b0011011000101011101: color_data = Z;
		19'b0011011000101011110: color_data = Z;
		19'b0011011000101011111: color_data = Z;
		19'b0011011000101100000: color_data = Z;
		19'b0011011000101100001: color_data = Z;
		19'b0011011000101100010: color_data = Z;
		19'b0011011000101100011: color_data = Z;
		19'b0011011000101100100: color_data = Z;
		19'b0011011000101100101: color_data = Z;
		19'b0011011000101100110: color_data = Z;
		19'b0011011000101100111: color_data = Z;
		19'b0011011000101101000: color_data = Z;
		19'b0011011000101101001: color_data = Z;
		19'b0011011000101101010: color_data = Z;
		19'b0011011000101101011: color_data = Z;
		19'b0011011000101101100: color_data = Z;
		19'b0011011000101101101: color_data = Z;
		19'b0011011000101101110: color_data = Z;
		19'b0011011000101101111: color_data = Z;
		19'b0011011000101110000: color_data = Z;
		19'b0011011000101110001: color_data = Z;
		19'b0011011000101110010: color_data = Z;
		19'b0011011000101110011: color_data = Z;
		19'b0011011000101110100: color_data = Z;
		19'b0011011000101110101: color_data = Z;
		19'b0011011000101110110: color_data = Z;
		19'b0011011000101110111: color_data = Z;
		19'b0011011000101111000: color_data = Z;
		19'b0011011000101111001: color_data = Z;
		19'b0011011000101111010: color_data = Z;
		19'b0011011000101111011: color_data = Z;
		19'b0011011000101111100: color_data = Z;
		19'b0011011000101111101: color_data = Z;
		19'b0011011000101111110: color_data = Z;
		19'b0011011000101111111: color_data = Z;
		19'b0011011000110000000: color_data = Z;
		19'b0011011000110000001: color_data = Z;
		19'b0011011000110000010: color_data = Z;
		19'b0011011000110000011: color_data = Z;
		19'b0011011000110000100: color_data = Z;
		19'b0011011000110000101: color_data = Z;
		19'b0011011000110000110: color_data = Z;
		19'b0011011000110000111: color_data = Z;
		19'b0011011000110001000: color_data = Z;
		19'b0011011000110001001: color_data = Z;
		19'b0011011000110001010: color_data = Z;
		19'b0011011000110001011: color_data = Z;
		19'b0011011000110001100: color_data = Z;
		19'b0011011000110001101: color_data = Z;
		19'b0011011000110001110: color_data = Z;
		19'b0011011000110001111: color_data = Z;
		19'b0011011000110010000: color_data = Z;
		19'b0011011000110010001: color_data = Z;
		19'b0011011000110010010: color_data = Z;
		19'b0011011000110010011: color_data = Z;
		19'b0011011000110010100: color_data = Z;
		19'b0011011000110010101: color_data = Z;
		19'b0011011000110010110: color_data = Z;
		19'b0011011000110111000: color_data = Z;
		19'b0011011000110111001: color_data = Z;
		19'b0011011000110111010: color_data = Z;
		19'b0011011000110111011: color_data = Z;
		19'b0011011000111011011: color_data = Z;
		19'b0011011010010101110: color_data = Z;
		19'b0011011010010101111: color_data = Z;
		19'b0011011010010110000: color_data = Z;
		19'b0011011010010110001: color_data = Z;
		19'b0011011010010110010: color_data = Z;
		19'b0011011010010110011: color_data = Z;
		19'b0011011010010110100: color_data = Z;
		19'b0011011010010110101: color_data = Z;
		19'b0011011010010110110: color_data = Z;
		19'b0011011010010110111: color_data = Z;
		19'b0011011010010111000: color_data = Z;
		19'b0011011010010111001: color_data = Z;
		19'b0011011010010111010: color_data = Z;
		19'b0011011010010111011: color_data = Z;
		19'b0011011010010111100: color_data = Z;
		19'b0011011010010111101: color_data = Z;
		19'b0011011010010111110: color_data = Z;
		19'b0011011010010111111: color_data = Z;
		19'b0011011010011000000: color_data = Z;
		19'b0011011010011000001: color_data = Z;
		19'b0011011010011000010: color_data = Z;
		19'b0011011010011000011: color_data = Z;
		19'b0011011010011000100: color_data = Z;
		19'b0011011010011000101: color_data = Z;
		19'b0011011010011000110: color_data = Z;
		19'b0011011010011000111: color_data = Z;
		19'b0011011010011001000: color_data = Z;
		19'b0011011010011001001: color_data = Z;
		19'b0011011010011001010: color_data = Z;
		19'b0011011010011001011: color_data = Z;
		19'b0011011010011001100: color_data = Z;
		19'b0011011010011001101: color_data = Z;
		19'b0011011010011001110: color_data = Z;
		19'b0011011010011001111: color_data = Z;
		19'b0011011010011010000: color_data = Z;
		19'b0011011010011010001: color_data = Z;
		19'b0011011010011010010: color_data = Z;
		19'b0011011010011010011: color_data = Z;
		19'b0011011010011010100: color_data = Z;
		19'b0011011010011010101: color_data = Z;
		19'b0011011010011010110: color_data = Z;
		19'b0011011010011010111: color_data = Z;
		19'b0011011010011011000: color_data = Z;
		19'b0011011010011011001: color_data = Z;
		19'b0011011010011011010: color_data = Z;
		19'b0011011010011011011: color_data = Z;
		19'b0011011010011011100: color_data = Z;
		19'b0011011010011011101: color_data = Z;
		19'b0011011010011011110: color_data = Z;
		19'b0011011010011011111: color_data = Z;
		19'b0011011010011100000: color_data = Z;
		19'b0011011010011100001: color_data = Z;
		19'b0011011010011100010: color_data = Z;
		19'b0011011010011100011: color_data = Z;
		19'b0011011010011100100: color_data = Z;
		19'b0011011010011100101: color_data = Z;
		19'b0011011010011100110: color_data = Z;
		19'b0011011010011100111: color_data = Z;
		19'b0011011010011101000: color_data = Z;
		19'b0011011010011101001: color_data = Z;
		19'b0011011010011101010: color_data = Z;
		19'b0011011010011101011: color_data = Z;
		19'b0011011010011101100: color_data = Z;
		19'b0011011010011101101: color_data = Z;
		19'b0011011010011101110: color_data = Z;
		19'b0011011010011101111: color_data = Z;
		19'b0011011010011110000: color_data = Z;
		19'b0011011010011110001: color_data = Z;
		19'b0011011010011110010: color_data = Z;
		19'b0011011010011110011: color_data = Z;
		19'b0011011010011110100: color_data = Z;
		19'b0011011010011110101: color_data = Z;
		19'b0011011010011110110: color_data = Z;
		19'b0011011010011110111: color_data = Z;
		19'b0011011010011111000: color_data = Z;
		19'b0011011010011111001: color_data = Z;
		19'b0011011010011111010: color_data = Z;
		19'b0011011010011111011: color_data = Z;
		19'b0011011010011111100: color_data = Z;
		19'b0011011010011111101: color_data = Z;
		19'b0011011010011111110: color_data = Z;
		19'b0011011010011111111: color_data = Z;
		19'b0011011010100000000: color_data = Z;
		19'b0011011010100000001: color_data = Z;
		19'b0011011010100000010: color_data = Z;
		19'b0011011010100000011: color_data = Z;
		19'b0011011010100000100: color_data = Z;
		19'b0011011010100000101: color_data = Z;
		19'b0011011010100000110: color_data = Z;
		19'b0011011010100000111: color_data = Z;
		19'b0011011010100001000: color_data = Z;
		19'b0011011010100001001: color_data = Z;
		19'b0011011010100001010: color_data = Z;
		19'b0011011010100001011: color_data = Z;
		19'b0011011010100001100: color_data = Z;
		19'b0011011010100001101: color_data = Z;
		19'b0011011010100001110: color_data = Z;
		19'b0011011010100001111: color_data = Z;
		19'b0011011010100010000: color_data = Z;
		19'b0011011010100010001: color_data = Z;
		19'b0011011010100010010: color_data = Z;
		19'b0011011010100010011: color_data = Z;
		19'b0011011010100010100: color_data = Z;
		19'b0011011010100010101: color_data = Z;
		19'b0011011010100010110: color_data = Z;
		19'b0011011010100010111: color_data = Z;
		19'b0011011010100011000: color_data = Z;
		19'b0011011010100011001: color_data = Z;
		19'b0011011010100011010: color_data = Z;
		19'b0011011010100011011: color_data = Z;
		19'b0011011010100011100: color_data = Z;
		19'b0011011010100011101: color_data = Z;
		19'b0011011010100011110: color_data = Z;
		19'b0011011010100011111: color_data = Z;
		19'b0011011010100100000: color_data = Z;
		19'b0011011010100100001: color_data = Z;
		19'b0011011010100100010: color_data = Z;
		19'b0011011010100100011: color_data = Z;
		19'b0011011010100100100: color_data = Z;
		19'b0011011010100100101: color_data = Z;
		19'b0011011010100100110: color_data = Z;
		19'b0011011010100100111: color_data = Z;
		19'b0011011010100101000: color_data = Z;
		19'b0011011010100101001: color_data = Z;
		19'b0011011010100101010: color_data = Z;
		19'b0011011010100101011: color_data = Z;
		19'b0011011010100101100: color_data = Z;
		19'b0011011010100101101: color_data = Z;
		19'b0011011010100101110: color_data = Z;
		19'b0011011010100101111: color_data = Z;
		19'b0011011010100110000: color_data = Z;
		19'b0011011010100110001: color_data = Z;
		19'b0011011010100110010: color_data = Z;
		19'b0011011010100110011: color_data = Z;
		19'b0011011010100110100: color_data = Z;
		19'b0011011010100110101: color_data = Z;
		19'b0011011010100110110: color_data = Z;
		19'b0011011010100110111: color_data = Z;
		19'b0011011010100111000: color_data = Z;
		19'b0011011010100111001: color_data = Z;
		19'b0011011010100111010: color_data = Z;
		19'b0011011010100111011: color_data = Z;
		19'b0011011010100111100: color_data = Z;
		19'b0011011010100111101: color_data = Z;
		19'b0011011010100111110: color_data = Z;
		19'b0011011010100111111: color_data = Z;
		19'b0011011010101000000: color_data = Z;
		19'b0011011010101000001: color_data = Z;
		19'b0011011010101000010: color_data = Z;
		19'b0011011010101000011: color_data = Z;
		19'b0011011010101000100: color_data = Z;
		19'b0011011010101000101: color_data = Z;
		19'b0011011010101000110: color_data = Z;
		19'b0011011010101000111: color_data = Z;
		19'b0011011010101001000: color_data = Z;
		19'b0011011010101001001: color_data = Z;
		19'b0011011010101001010: color_data = Z;
		19'b0011011010101001011: color_data = Z;
		19'b0011011010101001100: color_data = Z;
		19'b0011011010101001101: color_data = Z;
		19'b0011011010101001110: color_data = Z;
		19'b0011011010101001111: color_data = Z;
		19'b0011011010101010000: color_data = Z;
		19'b0011011010101010001: color_data = Z;
		19'b0011011010101010010: color_data = Z;
		19'b0011011010101010011: color_data = Z;
		19'b0011011010101010100: color_data = Z;
		19'b0011011010101010101: color_data = Z;
		19'b0011011010101010110: color_data = Z;
		19'b0011011010101010111: color_data = Z;
		19'b0011011010101011000: color_data = Z;
		19'b0011011010101011001: color_data = Z;
		19'b0011011010101011010: color_data = Z;
		19'b0011011010101011011: color_data = Z;
		19'b0011011010101011100: color_data = Z;
		19'b0011011010101011101: color_data = Z;
		19'b0011011010101011110: color_data = Z;
		19'b0011011010101011111: color_data = Z;
		19'b0011011010101100000: color_data = Z;
		19'b0011011010101100001: color_data = Z;
		19'b0011011010101100010: color_data = Z;
		19'b0011011010101100011: color_data = Z;
		19'b0011011010101100100: color_data = Z;
		19'b0011011010101100101: color_data = Z;
		19'b0011011010101100110: color_data = Z;
		19'b0011011010101100111: color_data = Z;
		19'b0011011010101101000: color_data = Z;
		19'b0011011010101101001: color_data = Z;
		19'b0011011010101101010: color_data = Z;
		19'b0011011010101101011: color_data = Z;
		19'b0011011010101101100: color_data = Z;
		19'b0011011010101101101: color_data = Z;
		19'b0011011010101101110: color_data = Z;
		19'b0011011010101101111: color_data = Z;
		19'b0011011010101110000: color_data = Z;
		19'b0011011010101110001: color_data = Z;
		19'b0011011010101110010: color_data = Z;
		19'b0011011010101110011: color_data = Z;
		19'b0011011010101110100: color_data = Z;
		19'b0011011010101110101: color_data = Z;
		19'b0011011010101110110: color_data = Z;
		19'b0011011010101110111: color_data = Z;
		19'b0011011010101111000: color_data = Z;
		19'b0011011010101111001: color_data = Z;
		19'b0011011010101111010: color_data = Z;
		19'b0011011010101111011: color_data = Z;
		19'b0011011010101111100: color_data = Z;
		19'b0011011010101111101: color_data = Z;
		19'b0011011010101111110: color_data = Z;
		19'b0011011010101111111: color_data = Z;
		19'b0011011010110000000: color_data = Z;
		19'b0011011010110000001: color_data = Z;
		19'b0011011010110000010: color_data = Z;
		19'b0011011010110000011: color_data = Z;
		19'b0011011010110000100: color_data = Z;
		19'b0011011010110000101: color_data = Z;
		19'b0011011010110000110: color_data = Z;
		19'b0011011010110000111: color_data = Z;
		19'b0011011010110001000: color_data = Z;
		19'b0011011010110001001: color_data = Z;
		19'b0011011010110001010: color_data = Z;
		19'b0011011010110001011: color_data = Z;
		19'b0011011010110001100: color_data = Z;
		19'b0011011010110001101: color_data = Z;
		19'b0011011010110001110: color_data = Z;
		19'b0011011010110001111: color_data = Z;
		19'b0011011010110010000: color_data = Z;
		19'b0011011010110010001: color_data = Z;
		19'b0011011010110010010: color_data = Z;
		19'b0011011010110010011: color_data = Z;
		19'b0011011010110010100: color_data = Z;
		19'b0011011010110010101: color_data = Z;
		19'b0011011010110010110: color_data = Z;
		19'b0011011010110111001: color_data = Z;
		19'b0011011010110111010: color_data = Z;
		19'b0011011010110111011: color_data = Z;
		19'b0011011010110111100: color_data = Z;
		19'b0011011010111011100: color_data = Z;
		19'b0011011100010101110: color_data = Z;
		19'b0011011100010101111: color_data = Z;
		19'b0011011100010110000: color_data = Z;
		19'b0011011100010110001: color_data = Z;
		19'b0011011100010110010: color_data = Z;
		19'b0011011100010110011: color_data = Z;
		19'b0011011100010110100: color_data = Z;
		19'b0011011100010110101: color_data = Z;
		19'b0011011100010110110: color_data = Z;
		19'b0011011100010110111: color_data = Z;
		19'b0011011100010111000: color_data = Z;
		19'b0011011100010111001: color_data = Z;
		19'b0011011100010111010: color_data = Z;
		19'b0011011100010111011: color_data = Z;
		19'b0011011100010111100: color_data = Z;
		19'b0011011100010111101: color_data = Z;
		19'b0011011100010111110: color_data = Z;
		19'b0011011100010111111: color_data = Z;
		19'b0011011100011000000: color_data = Z;
		19'b0011011100011000001: color_data = Z;
		19'b0011011100011000010: color_data = Z;
		19'b0011011100011000011: color_data = Z;
		19'b0011011100011000100: color_data = Z;
		19'b0011011100011000101: color_data = Z;
		19'b0011011100011000110: color_data = Z;
		19'b0011011100011000111: color_data = Z;
		19'b0011011100011001000: color_data = Z;
		19'b0011011100011001001: color_data = Z;
		19'b0011011100011001010: color_data = Z;
		19'b0011011100011001011: color_data = Z;
		19'b0011011100011001100: color_data = Z;
		19'b0011011100011001101: color_data = Z;
		19'b0011011100011001110: color_data = Z;
		19'b0011011100011001111: color_data = Z;
		19'b0011011100011010000: color_data = Z;
		19'b0011011100011010001: color_data = Z;
		19'b0011011100011010010: color_data = Z;
		19'b0011011100011010011: color_data = Z;
		19'b0011011100011010100: color_data = Z;
		19'b0011011100011010101: color_data = Z;
		19'b0011011100011010110: color_data = Z;
		19'b0011011100011010111: color_data = Z;
		19'b0011011100011011000: color_data = Z;
		19'b0011011100011011001: color_data = Z;
		19'b0011011100011011010: color_data = Z;
		19'b0011011100011011011: color_data = Z;
		19'b0011011100011011100: color_data = Z;
		19'b0011011100011011101: color_data = Z;
		19'b0011011100011011110: color_data = Z;
		19'b0011011100011011111: color_data = Z;
		19'b0011011100011100000: color_data = Z;
		19'b0011011100011100001: color_data = Z;
		19'b0011011100011100010: color_data = Z;
		19'b0011011100011100011: color_data = Z;
		19'b0011011100011100100: color_data = Z;
		19'b0011011100011100101: color_data = Z;
		19'b0011011100011100110: color_data = Z;
		19'b0011011100011100111: color_data = Z;
		19'b0011011100011101000: color_data = Z;
		19'b0011011100011101001: color_data = Z;
		19'b0011011100011101010: color_data = Z;
		19'b0011011100011101011: color_data = Z;
		19'b0011011100011101100: color_data = Z;
		19'b0011011100011101101: color_data = Z;
		19'b0011011100011101110: color_data = Z;
		19'b0011011100011101111: color_data = Z;
		19'b0011011100011110000: color_data = Z;
		19'b0011011100011110001: color_data = Z;
		19'b0011011100011110010: color_data = Z;
		19'b0011011100011110011: color_data = Z;
		19'b0011011100011110100: color_data = Z;
		19'b0011011100011110101: color_data = Z;
		19'b0011011100011110110: color_data = Z;
		19'b0011011100011110111: color_data = Z;
		19'b0011011100011111000: color_data = Z;
		19'b0011011100011111001: color_data = Z;
		19'b0011011100011111010: color_data = Z;
		19'b0011011100011111011: color_data = Z;
		19'b0011011100011111100: color_data = Z;
		19'b0011011100011111101: color_data = Z;
		19'b0011011100011111110: color_data = Z;
		19'b0011011100011111111: color_data = Z;
		19'b0011011100100000000: color_data = Z;
		19'b0011011100100000001: color_data = Z;
		19'b0011011100100000010: color_data = Z;
		19'b0011011100100000011: color_data = Z;
		19'b0011011100100000100: color_data = Z;
		19'b0011011100100000101: color_data = Z;
		19'b0011011100100000110: color_data = Z;
		19'b0011011100100000111: color_data = Z;
		19'b0011011100100001000: color_data = Z;
		19'b0011011100100001001: color_data = Z;
		19'b0011011100100001010: color_data = Z;
		19'b0011011100100001011: color_data = Z;
		19'b0011011100100001100: color_data = Z;
		19'b0011011100100001101: color_data = Z;
		19'b0011011100100001110: color_data = Z;
		19'b0011011100100001111: color_data = Z;
		19'b0011011100100010000: color_data = Z;
		19'b0011011100100010001: color_data = Z;
		19'b0011011100100010010: color_data = Z;
		19'b0011011100100010011: color_data = Z;
		19'b0011011100100010100: color_data = Z;
		19'b0011011100100010101: color_data = Z;
		19'b0011011100100010110: color_data = Z;
		19'b0011011100100010111: color_data = Z;
		19'b0011011100100011000: color_data = Z;
		19'b0011011100100011001: color_data = Z;
		19'b0011011100100011010: color_data = Z;
		19'b0011011100100011011: color_data = Z;
		19'b0011011100100011100: color_data = Z;
		19'b0011011100100011101: color_data = Z;
		19'b0011011100100011110: color_data = Z;
		19'b0011011100100011111: color_data = Z;
		19'b0011011100100100000: color_data = Z;
		19'b0011011100100100001: color_data = Z;
		19'b0011011100100100010: color_data = Z;
		19'b0011011100100100011: color_data = Z;
		19'b0011011100100100100: color_data = Z;
		19'b0011011100100100101: color_data = Z;
		19'b0011011100100100110: color_data = Z;
		19'b0011011100100100111: color_data = Z;
		19'b0011011100100101000: color_data = Z;
		19'b0011011100100101001: color_data = Z;
		19'b0011011100100101010: color_data = Z;
		19'b0011011100100101011: color_data = Z;
		19'b0011011100100101100: color_data = Z;
		19'b0011011100100101101: color_data = Z;
		19'b0011011100100101110: color_data = Z;
		19'b0011011100100101111: color_data = Z;
		19'b0011011100100110000: color_data = Z;
		19'b0011011100100110001: color_data = Z;
		19'b0011011100100110010: color_data = Z;
		19'b0011011100100110011: color_data = Z;
		19'b0011011100100110100: color_data = Z;
		19'b0011011100100110101: color_data = Z;
		19'b0011011100100110110: color_data = Z;
		19'b0011011100100110111: color_data = Z;
		19'b0011011100100111000: color_data = Z;
		19'b0011011100100111001: color_data = Z;
		19'b0011011100100111010: color_data = Z;
		19'b0011011100100111011: color_data = Z;
		19'b0011011100100111100: color_data = Z;
		19'b0011011100100111101: color_data = Z;
		19'b0011011100100111110: color_data = Z;
		19'b0011011100100111111: color_data = Z;
		19'b0011011100101000000: color_data = Z;
		19'b0011011100101000001: color_data = Z;
		19'b0011011100101000010: color_data = Z;
		19'b0011011100101000011: color_data = Z;
		19'b0011011100101000100: color_data = Z;
		19'b0011011100101000101: color_data = Z;
		19'b0011011100101000110: color_data = Z;
		19'b0011011100101000111: color_data = Z;
		19'b0011011100101001000: color_data = Z;
		19'b0011011100101001001: color_data = Z;
		19'b0011011100101001010: color_data = Z;
		19'b0011011100101001011: color_data = Z;
		19'b0011011100101001100: color_data = Z;
		19'b0011011100101001101: color_data = Z;
		19'b0011011100101001110: color_data = Z;
		19'b0011011100101001111: color_data = Z;
		19'b0011011100101010000: color_data = Z;
		19'b0011011100101010001: color_data = Z;
		19'b0011011100101010010: color_data = Z;
		19'b0011011100101010011: color_data = Z;
		19'b0011011100101010100: color_data = Z;
		19'b0011011100101010101: color_data = Z;
		19'b0011011100101010110: color_data = Z;
		19'b0011011100101010111: color_data = Z;
		19'b0011011100101011000: color_data = Z;
		19'b0011011100101011001: color_data = Z;
		19'b0011011100101011010: color_data = Z;
		19'b0011011100101011011: color_data = Z;
		19'b0011011100101011100: color_data = Z;
		19'b0011011100101011101: color_data = Z;
		19'b0011011100101011110: color_data = Z;
		19'b0011011100101011111: color_data = Z;
		19'b0011011100101100000: color_data = Z;
		19'b0011011100101100001: color_data = Z;
		19'b0011011100101100010: color_data = Z;
		19'b0011011100101100011: color_data = Z;
		19'b0011011100101100100: color_data = Z;
		19'b0011011100101100101: color_data = Z;
		19'b0011011100101100110: color_data = Z;
		19'b0011011100101100111: color_data = Z;
		19'b0011011100101101000: color_data = Z;
		19'b0011011100101101001: color_data = Z;
		19'b0011011100101101010: color_data = Z;
		19'b0011011100101101011: color_data = Z;
		19'b0011011100101101100: color_data = Z;
		19'b0011011100101101101: color_data = Z;
		19'b0011011100101101110: color_data = Z;
		19'b0011011100101101111: color_data = Z;
		19'b0011011100101110000: color_data = Z;
		19'b0011011100101110001: color_data = Z;
		19'b0011011100101110010: color_data = Z;
		19'b0011011100101110011: color_data = Z;
		19'b0011011100101110100: color_data = Z;
		19'b0011011100101110101: color_data = Z;
		19'b0011011100101110110: color_data = Z;
		19'b0011011100101110111: color_data = Z;
		19'b0011011100101111000: color_data = Z;
		19'b0011011100101111001: color_data = Z;
		19'b0011011100101111010: color_data = Z;
		19'b0011011100101111011: color_data = Z;
		19'b0011011100101111100: color_data = Z;
		19'b0011011100101111101: color_data = Z;
		19'b0011011100101111110: color_data = Z;
		19'b0011011100101111111: color_data = Z;
		19'b0011011100110000000: color_data = Z;
		19'b0011011100110000001: color_data = Z;
		19'b0011011100110000010: color_data = Z;
		19'b0011011100110000011: color_data = Z;
		19'b0011011100110000100: color_data = Z;
		19'b0011011100110000101: color_data = Z;
		19'b0011011100110000110: color_data = Z;
		19'b0011011100110000111: color_data = Z;
		19'b0011011100110001000: color_data = Z;
		19'b0011011100110001001: color_data = Z;
		19'b0011011100110001010: color_data = Z;
		19'b0011011100110001011: color_data = Z;
		19'b0011011100110001100: color_data = Z;
		19'b0011011100110001101: color_data = Z;
		19'b0011011100110001110: color_data = Z;
		19'b0011011100110001111: color_data = Z;
		19'b0011011100110010000: color_data = Z;
		19'b0011011100110010001: color_data = Z;
		19'b0011011100110010010: color_data = Z;
		19'b0011011100110010011: color_data = Z;
		19'b0011011100110010100: color_data = Z;
		19'b0011011100110111001: color_data = Z;
		19'b0011011100110111010: color_data = Z;
		19'b0011011100110111011: color_data = Z;
		19'b0011011100110111100: color_data = Z;
		19'b0011011100110111101: color_data = Z;
		19'b0011011100111011100: color_data = Z;
		19'b0011011110010101110: color_data = Z;
		19'b0011011110010101111: color_data = Z;
		19'b0011011110010110000: color_data = Z;
		19'b0011011110010110001: color_data = Z;
		19'b0011011110010110010: color_data = Z;
		19'b0011011110010110011: color_data = Z;
		19'b0011011110010110100: color_data = Z;
		19'b0011011110010110101: color_data = Z;
		19'b0011011110010110110: color_data = Z;
		19'b0011011110010110111: color_data = Z;
		19'b0011011110010111000: color_data = Z;
		19'b0011011110010111001: color_data = Z;
		19'b0011011110010111010: color_data = Z;
		19'b0011011110010111011: color_data = Z;
		19'b0011011110010111100: color_data = Z;
		19'b0011011110010111101: color_data = Z;
		19'b0011011110010111110: color_data = Z;
		19'b0011011110010111111: color_data = Z;
		19'b0011011110011000000: color_data = Z;
		19'b0011011110011000001: color_data = Z;
		19'b0011011110011000010: color_data = Z;
		19'b0011011110011000011: color_data = Z;
		19'b0011011110011000100: color_data = Z;
		19'b0011011110011000101: color_data = Z;
		19'b0011011110011000110: color_data = Z;
		19'b0011011110011000111: color_data = Z;
		19'b0011011110011001000: color_data = Z;
		19'b0011011110011001001: color_data = Z;
		19'b0011011110011001010: color_data = Z;
		19'b0011011110011001011: color_data = Z;
		19'b0011011110011001100: color_data = Z;
		19'b0011011110011001101: color_data = Z;
		19'b0011011110011001110: color_data = Z;
		19'b0011011110011001111: color_data = Z;
		19'b0011011110011010000: color_data = Z;
		19'b0011011110011010001: color_data = Z;
		19'b0011011110011010010: color_data = Z;
		19'b0011011110011010011: color_data = Z;
		19'b0011011110011010100: color_data = Z;
		19'b0011011110011010101: color_data = Z;
		19'b0011011110011010110: color_data = Z;
		19'b0011011110011010111: color_data = Z;
		19'b0011011110011011000: color_data = Z;
		19'b0011011110011011001: color_data = Z;
		19'b0011011110011011010: color_data = Z;
		19'b0011011110011011011: color_data = Z;
		19'b0011011110011011100: color_data = Z;
		19'b0011011110011011101: color_data = Z;
		19'b0011011110011011110: color_data = Z;
		19'b0011011110011011111: color_data = Z;
		19'b0011011110011100000: color_data = Z;
		19'b0011011110011100001: color_data = Z;
		19'b0011011110011100010: color_data = Z;
		19'b0011011110011100011: color_data = Z;
		19'b0011011110011100100: color_data = Z;
		19'b0011011110011100101: color_data = Z;
		19'b0011011110011100110: color_data = Z;
		19'b0011011110011100111: color_data = Z;
		19'b0011011110011101000: color_data = Z;
		19'b0011011110011101001: color_data = Z;
		19'b0011011110011101010: color_data = Z;
		19'b0011011110011101011: color_data = Z;
		19'b0011011110011101100: color_data = Z;
		19'b0011011110011101101: color_data = Z;
		19'b0011011110011101110: color_data = Z;
		19'b0011011110011101111: color_data = Z;
		19'b0011011110011110000: color_data = Z;
		19'b0011011110011110001: color_data = Z;
		19'b0011011110011110010: color_data = Z;
		19'b0011011110011110011: color_data = Z;
		19'b0011011110011110100: color_data = Z;
		19'b0011011110011110101: color_data = Z;
		19'b0011011110011110110: color_data = Z;
		19'b0011011110011110111: color_data = Z;
		19'b0011011110011111000: color_data = Z;
		19'b0011011110011111001: color_data = Z;
		19'b0011011110011111010: color_data = Z;
		19'b0011011110011111011: color_data = Z;
		19'b0011011110011111100: color_data = Z;
		19'b0011011110011111101: color_data = Z;
		19'b0011011110011111110: color_data = Z;
		19'b0011011110011111111: color_data = Z;
		19'b0011011110100000000: color_data = Z;
		19'b0011011110100000001: color_data = Z;
		19'b0011011110100000010: color_data = Z;
		19'b0011011110100000011: color_data = Z;
		19'b0011011110100000100: color_data = Z;
		19'b0011011110100000101: color_data = Z;
		19'b0011011110100000110: color_data = Z;
		19'b0011011110100000111: color_data = Z;
		19'b0011011110100001000: color_data = Z;
		19'b0011011110100001001: color_data = Z;
		19'b0011011110100001010: color_data = Z;
		19'b0011011110100001011: color_data = Z;
		19'b0011011110100001100: color_data = Z;
		19'b0011011110100001101: color_data = Z;
		19'b0011011110100001110: color_data = Z;
		19'b0011011110100001111: color_data = Z;
		19'b0011011110100010000: color_data = Z;
		19'b0011011110100010001: color_data = Z;
		19'b0011011110100010010: color_data = Z;
		19'b0011011110100010011: color_data = Z;
		19'b0011011110100010100: color_data = Z;
		19'b0011011110100010101: color_data = Z;
		19'b0011011110100010110: color_data = Z;
		19'b0011011110100010111: color_data = Z;
		19'b0011011110100011000: color_data = Z;
		19'b0011011110100011001: color_data = Z;
		19'b0011011110100011010: color_data = Z;
		19'b0011011110100011011: color_data = Z;
		19'b0011011110100011100: color_data = Z;
		19'b0011011110100011101: color_data = Z;
		19'b0011011110100011110: color_data = Z;
		19'b0011011110100011111: color_data = Z;
		19'b0011011110100100000: color_data = Z;
		19'b0011011110100100001: color_data = Z;
		19'b0011011110100100010: color_data = Z;
		19'b0011011110100100011: color_data = Z;
		19'b0011011110100100100: color_data = Z;
		19'b0011011110100100101: color_data = Z;
		19'b0011011110100100110: color_data = Z;
		19'b0011011110100100111: color_data = Z;
		19'b0011011110100101000: color_data = Z;
		19'b0011011110100101001: color_data = Z;
		19'b0011011110100101010: color_data = Z;
		19'b0011011110100101011: color_data = Z;
		19'b0011011110100101100: color_data = Z;
		19'b0011011110100101101: color_data = Z;
		19'b0011011110100101110: color_data = Z;
		19'b0011011110100101111: color_data = Z;
		19'b0011011110100110000: color_data = Z;
		19'b0011011110100110001: color_data = Z;
		19'b0011011110100110010: color_data = Z;
		19'b0011011110100110011: color_data = Z;
		19'b0011011110100110100: color_data = Z;
		19'b0011011110100110101: color_data = Z;
		19'b0011011110100110110: color_data = Z;
		19'b0011011110100110111: color_data = Z;
		19'b0011011110100111000: color_data = Z;
		19'b0011011110100111001: color_data = Z;
		19'b0011011110100111010: color_data = Z;
		19'b0011011110100111011: color_data = Z;
		19'b0011011110100111100: color_data = Z;
		19'b0011011110100111101: color_data = Z;
		19'b0011011110100111110: color_data = Z;
		19'b0011011110100111111: color_data = Z;
		19'b0011011110101000000: color_data = Z;
		19'b0011011110101000001: color_data = Z;
		19'b0011011110101000010: color_data = Z;
		19'b0011011110101000011: color_data = Z;
		19'b0011011110101000100: color_data = Z;
		19'b0011011110101000101: color_data = Z;
		19'b0011011110101000110: color_data = Z;
		19'b0011011110101000111: color_data = Z;
		19'b0011011110101001000: color_data = Z;
		19'b0011011110101001001: color_data = Z;
		19'b0011011110101001010: color_data = Z;
		19'b0011011110101001011: color_data = Z;
		19'b0011011110101001100: color_data = Z;
		19'b0011011110101001101: color_data = Z;
		19'b0011011110101001110: color_data = Z;
		19'b0011011110101001111: color_data = Z;
		19'b0011011110101010000: color_data = Z;
		19'b0011011110101010001: color_data = Z;
		19'b0011011110101010010: color_data = Z;
		19'b0011011110101010011: color_data = Z;
		19'b0011011110101010100: color_data = Z;
		19'b0011011110101010101: color_data = Z;
		19'b0011011110101010110: color_data = Z;
		19'b0011011110101010111: color_data = Z;
		19'b0011011110101011000: color_data = Z;
		19'b0011011110101011001: color_data = Z;
		19'b0011011110101011010: color_data = Z;
		19'b0011011110101011011: color_data = Z;
		19'b0011011110101011100: color_data = Z;
		19'b0011011110101011101: color_data = Z;
		19'b0011011110101011110: color_data = Z;
		19'b0011011110101011111: color_data = Z;
		19'b0011011110101100000: color_data = Z;
		19'b0011011110101100001: color_data = Z;
		19'b0011011110101100010: color_data = Z;
		19'b0011011110101100011: color_data = Z;
		19'b0011011110101100100: color_data = Z;
		19'b0011011110101100101: color_data = Z;
		19'b0011011110101100110: color_data = Z;
		19'b0011011110101100111: color_data = Z;
		19'b0011011110101101000: color_data = Z;
		19'b0011011110101101001: color_data = Z;
		19'b0011011110101101010: color_data = Z;
		19'b0011011110101101011: color_data = Z;
		19'b0011011110101101100: color_data = Z;
		19'b0011011110101101101: color_data = Z;
		19'b0011011110101101110: color_data = Z;
		19'b0011011110101101111: color_data = Z;
		19'b0011011110101110000: color_data = Z;
		19'b0011011110101110001: color_data = Z;
		19'b0011011110101110010: color_data = Z;
		19'b0011011110101110011: color_data = Z;
		19'b0011011110101110100: color_data = Z;
		19'b0011011110101110101: color_data = Z;
		19'b0011011110101110110: color_data = Z;
		19'b0011011110101110111: color_data = Z;
		19'b0011011110101111000: color_data = Z;
		19'b0011011110101111001: color_data = Z;
		19'b0011011110101111010: color_data = Z;
		19'b0011011110101111011: color_data = Z;
		19'b0011011110101111100: color_data = Z;
		19'b0011011110101111101: color_data = Z;
		19'b0011011110101111110: color_data = Z;
		19'b0011011110101111111: color_data = Z;
		19'b0011011110110000000: color_data = Z;
		19'b0011011110110000001: color_data = Z;
		19'b0011011110110000010: color_data = Z;
		19'b0011011110110000011: color_data = Z;
		19'b0011011110110000100: color_data = Z;
		19'b0011011110110000101: color_data = Z;
		19'b0011011110110000110: color_data = Z;
		19'b0011011110110000111: color_data = Z;
		19'b0011011110110001000: color_data = Z;
		19'b0011011110110001001: color_data = Z;
		19'b0011011110110001010: color_data = Z;
		19'b0011011110110001011: color_data = Z;
		19'b0011011110110001100: color_data = Z;
		19'b0011011110110001101: color_data = Z;
		19'b0011011110110001110: color_data = Z;
		19'b0011011110110001111: color_data = Z;
		19'b0011011110110010000: color_data = Z;
		19'b0011011110110010001: color_data = Z;
		19'b0011011110110010010: color_data = Z;
		19'b0011011110110010011: color_data = Z;
		19'b0011011110110010100: color_data = Z;
		19'b0011011110110111001: color_data = Z;
		19'b0011011110110111010: color_data = Z;
		19'b0011011110110111011: color_data = Z;
		19'b0011011110110111100: color_data = Z;
		19'b0011011110110111101: color_data = Z;
		19'b0011011110111011100: color_data = Z;
		19'b0011100000010101110: color_data = Z;
		19'b0011100000010101111: color_data = Z;
		19'b0011100000010110000: color_data = Z;
		19'b0011100000010110001: color_data = Z;
		19'b0011100000010110010: color_data = Z;
		19'b0011100000010110011: color_data = Z;
		19'b0011100000010110100: color_data = Z;
		19'b0011100000010110101: color_data = Z;
		19'b0011100000010110110: color_data = Z;
		19'b0011100000010110111: color_data = Z;
		19'b0011100000010111000: color_data = Z;
		19'b0011100000010111001: color_data = Z;
		19'b0011100000010111010: color_data = Z;
		19'b0011100000010111011: color_data = Z;
		19'b0011100000010111100: color_data = Z;
		19'b0011100000010111101: color_data = Z;
		19'b0011100000010111110: color_data = Z;
		19'b0011100000010111111: color_data = Z;
		19'b0011100000011000000: color_data = Z;
		19'b0011100000011000001: color_data = Z;
		19'b0011100000011000010: color_data = Z;
		19'b0011100000011000011: color_data = Z;
		19'b0011100000011000100: color_data = Z;
		19'b0011100000011000101: color_data = Z;
		19'b0011100000011000110: color_data = Z;
		19'b0011100000011000111: color_data = Z;
		19'b0011100000011001000: color_data = Z;
		19'b0011100000011001001: color_data = Z;
		19'b0011100000011001010: color_data = Z;
		19'b0011100000011001011: color_data = Z;
		19'b0011100000011001100: color_data = Z;
		19'b0011100000011001101: color_data = Z;
		19'b0011100000011001110: color_data = Z;
		19'b0011100000011001111: color_data = Z;
		19'b0011100000011010000: color_data = Z;
		19'b0011100000011010001: color_data = Z;
		19'b0011100000011010010: color_data = Z;
		19'b0011100000011010011: color_data = Z;
		19'b0011100000011010100: color_data = Z;
		19'b0011100000011010101: color_data = Z;
		19'b0011100000011010110: color_data = Z;
		19'b0011100000011010111: color_data = Z;
		19'b0011100000011011000: color_data = Z;
		19'b0011100000011011001: color_data = Z;
		19'b0011100000011011010: color_data = Z;
		19'b0011100000011011011: color_data = Z;
		19'b0011100000011011100: color_data = Z;
		19'b0011100000011011101: color_data = Z;
		19'b0011100000011011110: color_data = Z;
		19'b0011100000011011111: color_data = Z;
		19'b0011100000011100000: color_data = Z;
		19'b0011100000011100001: color_data = Z;
		19'b0011100000011100010: color_data = Z;
		19'b0011100000011100011: color_data = Z;
		19'b0011100000011100100: color_data = Z;
		19'b0011100000011100101: color_data = Z;
		19'b0011100000011100110: color_data = Z;
		19'b0011100000011100111: color_data = Z;
		19'b0011100000011101000: color_data = Z;
		19'b0011100000011101001: color_data = Z;
		19'b0011100000011101010: color_data = Z;
		19'b0011100000011101011: color_data = Z;
		19'b0011100000011101100: color_data = Z;
		19'b0011100000011101101: color_data = Z;
		19'b0011100000011101110: color_data = Z;
		19'b0011100000011101111: color_data = Z;
		19'b0011100000011110000: color_data = Z;
		19'b0011100000011110001: color_data = Z;
		19'b0011100000011110010: color_data = Z;
		19'b0011100000011110011: color_data = Z;
		19'b0011100000011110100: color_data = Z;
		19'b0011100000011110101: color_data = Z;
		19'b0011100000011110110: color_data = Z;
		19'b0011100000011110111: color_data = Z;
		19'b0011100000011111000: color_data = Z;
		19'b0011100000011111001: color_data = Z;
		19'b0011100000011111010: color_data = Z;
		19'b0011100000011111011: color_data = Z;
		19'b0011100000011111100: color_data = Z;
		19'b0011100000011111101: color_data = Z;
		19'b0011100000011111110: color_data = Z;
		19'b0011100000011111111: color_data = Z;
		19'b0011100000100000000: color_data = Z;
		19'b0011100000100000001: color_data = Z;
		19'b0011100000100000010: color_data = Z;
		19'b0011100000100000011: color_data = Z;
		19'b0011100000100000100: color_data = Z;
		19'b0011100000100000101: color_data = Z;
		19'b0011100000100000110: color_data = Z;
		19'b0011100000100000111: color_data = Z;
		19'b0011100000100001000: color_data = Z;
		19'b0011100000100001001: color_data = Z;
		19'b0011100000100001010: color_data = Z;
		19'b0011100000100001011: color_data = Z;
		19'b0011100000100001100: color_data = Z;
		19'b0011100000100001101: color_data = Z;
		19'b0011100000100001110: color_data = Z;
		19'b0011100000100001111: color_data = Z;
		19'b0011100000100010000: color_data = Z;
		19'b0011100000100010001: color_data = Z;
		19'b0011100000100010010: color_data = Z;
		19'b0011100000100010011: color_data = Z;
		19'b0011100000100010100: color_data = Z;
		19'b0011100000100010101: color_data = Z;
		19'b0011100000100010110: color_data = Z;
		19'b0011100000100010111: color_data = Z;
		19'b0011100000100011000: color_data = Z;
		19'b0011100000100011001: color_data = Z;
		19'b0011100000100011010: color_data = Z;
		19'b0011100000100011011: color_data = Z;
		19'b0011100000100011100: color_data = Z;
		19'b0011100000100011101: color_data = Z;
		19'b0011100000100011110: color_data = Z;
		19'b0011100000100011111: color_data = Z;
		19'b0011100000100100000: color_data = Z;
		19'b0011100000100100001: color_data = Z;
		19'b0011100000100100010: color_data = Z;
		19'b0011100000100100011: color_data = Z;
		19'b0011100000100100100: color_data = Z;
		19'b0011100000100100101: color_data = Z;
		19'b0011100000100100110: color_data = Z;
		19'b0011100000100100111: color_data = Z;
		19'b0011100000100101000: color_data = Z;
		19'b0011100000100101001: color_data = Z;
		19'b0011100000100101010: color_data = Z;
		19'b0011100000100101011: color_data = Z;
		19'b0011100000100101100: color_data = Z;
		19'b0011100000100101101: color_data = Z;
		19'b0011100000100101110: color_data = Z;
		19'b0011100000100101111: color_data = Z;
		19'b0011100000100110000: color_data = Z;
		19'b0011100000100110001: color_data = Z;
		19'b0011100000100110010: color_data = Z;
		19'b0011100000100110011: color_data = Z;
		19'b0011100000100110100: color_data = Z;
		19'b0011100000100110101: color_data = Z;
		19'b0011100000100110110: color_data = Z;
		19'b0011100000100110111: color_data = Z;
		19'b0011100000100111000: color_data = Z;
		19'b0011100000100111001: color_data = Z;
		19'b0011100000100111010: color_data = Z;
		19'b0011100000100111011: color_data = Z;
		19'b0011100000100111100: color_data = Z;
		19'b0011100000100111101: color_data = Z;
		19'b0011100000100111110: color_data = Z;
		19'b0011100000100111111: color_data = Z;
		19'b0011100000101000000: color_data = Z;
		19'b0011100000101000001: color_data = Z;
		19'b0011100000101000010: color_data = Z;
		19'b0011100000101000011: color_data = Z;
		19'b0011100000101000100: color_data = Z;
		19'b0011100000101000101: color_data = Z;
		19'b0011100000101000110: color_data = Z;
		19'b0011100000101000111: color_data = Z;
		19'b0011100000101001000: color_data = Z;
		19'b0011100000101001001: color_data = Z;
		19'b0011100000101001010: color_data = Z;
		19'b0011100000101001011: color_data = Z;
		19'b0011100000101001100: color_data = Z;
		19'b0011100000101001101: color_data = Z;
		19'b0011100000101001110: color_data = Z;
		19'b0011100000101001111: color_data = Z;
		19'b0011100000101010000: color_data = Z;
		19'b0011100000101010001: color_data = Z;
		19'b0011100000101010010: color_data = Z;
		19'b0011100000101010011: color_data = Z;
		19'b0011100000101010100: color_data = Z;
		19'b0011100000101010101: color_data = Z;
		19'b0011100000101010110: color_data = Z;
		19'b0011100000101010111: color_data = Z;
		19'b0011100000101011000: color_data = Z;
		19'b0011100000101011001: color_data = Z;
		19'b0011100000101011010: color_data = Z;
		19'b0011100000101011011: color_data = Z;
		19'b0011100000101011100: color_data = Z;
		19'b0011100000101011101: color_data = Z;
		19'b0011100000101011110: color_data = Z;
		19'b0011100000101011111: color_data = Z;
		19'b0011100000101100000: color_data = Z;
		19'b0011100000101100001: color_data = Z;
		19'b0011100000101100010: color_data = Z;
		19'b0011100000101100011: color_data = Z;
		19'b0011100000101100100: color_data = Z;
		19'b0011100000101100101: color_data = Z;
		19'b0011100000101100110: color_data = Z;
		19'b0011100000101100111: color_data = Z;
		19'b0011100000101101000: color_data = Z;
		19'b0011100000101101001: color_data = Z;
		19'b0011100000101101010: color_data = Z;
		19'b0011100000101101011: color_data = Z;
		19'b0011100000101101100: color_data = Z;
		19'b0011100000101101101: color_data = Z;
		19'b0011100000101101110: color_data = Z;
		19'b0011100000101101111: color_data = Z;
		19'b0011100000101110000: color_data = Z;
		19'b0011100000101110001: color_data = Z;
		19'b0011100000101110010: color_data = Z;
		19'b0011100000101110011: color_data = Z;
		19'b0011100000101110100: color_data = Z;
		19'b0011100000101110101: color_data = Z;
		19'b0011100000101110110: color_data = Z;
		19'b0011100000101110111: color_data = Z;
		19'b0011100000101111000: color_data = Z;
		19'b0011100000101111001: color_data = Z;
		19'b0011100000101111010: color_data = Z;
		19'b0011100000101111011: color_data = Z;
		19'b0011100000101111100: color_data = Z;
		19'b0011100000101111101: color_data = Z;
		19'b0011100000101111110: color_data = Z;
		19'b0011100000101111111: color_data = Z;
		19'b0011100000110000000: color_data = Z;
		19'b0011100000110000001: color_data = Z;
		19'b0011100000110000010: color_data = Z;
		19'b0011100000110000011: color_data = Z;
		19'b0011100000110000100: color_data = Z;
		19'b0011100000110000101: color_data = Z;
		19'b0011100000110000110: color_data = Z;
		19'b0011100000110000111: color_data = Z;
		19'b0011100000110001000: color_data = Z;
		19'b0011100000110001001: color_data = Z;
		19'b0011100000110001010: color_data = Z;
		19'b0011100000110001011: color_data = Z;
		19'b0011100000110001100: color_data = Z;
		19'b0011100000110001101: color_data = Z;
		19'b0011100000110001110: color_data = Z;
		19'b0011100000110001111: color_data = Z;
		19'b0011100000110010000: color_data = Z;
		19'b0011100000110010001: color_data = Z;
		19'b0011100000110010010: color_data = Z;
		19'b0011100000110010011: color_data = Z;
		19'b0011100000110111001: color_data = Z;
		19'b0011100000110111010: color_data = Z;
		19'b0011100000110111011: color_data = Z;
		19'b0011100000110111100: color_data = Z;
		19'b0011100000110111101: color_data = Z;
		19'b0011100000110111110: color_data = Z;
		19'b0011100000110111111: color_data = Z;
		19'b0011100010010101101: color_data = Z;
		19'b0011100010010101110: color_data = Z;
		19'b0011100010010101111: color_data = Z;
		19'b0011100010010110000: color_data = Z;
		19'b0011100010010110001: color_data = Z;
		19'b0011100010010110010: color_data = Z;
		19'b0011100010010110011: color_data = Z;
		19'b0011100010010110100: color_data = Z;
		19'b0011100010010110101: color_data = Z;
		19'b0011100010010110110: color_data = Z;
		19'b0011100010010110111: color_data = Z;
		19'b0011100010010111000: color_data = Z;
		19'b0011100010010111001: color_data = Z;
		19'b0011100010010111010: color_data = Z;
		19'b0011100010010111011: color_data = Z;
		19'b0011100010010111100: color_data = Z;
		19'b0011100010010111101: color_data = Z;
		19'b0011100010010111110: color_data = Z;
		19'b0011100010010111111: color_data = Z;
		19'b0011100010011000000: color_data = Z;
		19'b0011100010011000001: color_data = Z;
		19'b0011100010011000010: color_data = Z;
		19'b0011100010011000011: color_data = Z;
		19'b0011100010011000100: color_data = Z;
		19'b0011100010011000101: color_data = Z;
		19'b0011100010011000110: color_data = Z;
		19'b0011100010011000111: color_data = Z;
		19'b0011100010011001000: color_data = Z;
		19'b0011100010011001001: color_data = Z;
		19'b0011100010011001010: color_data = Z;
		19'b0011100010011001011: color_data = Z;
		19'b0011100010011001100: color_data = Z;
		19'b0011100010011001101: color_data = Z;
		19'b0011100010011001110: color_data = Z;
		19'b0011100010011001111: color_data = Z;
		19'b0011100010011010000: color_data = Z;
		19'b0011100010011010001: color_data = Z;
		19'b0011100010011010010: color_data = Z;
		19'b0011100010011010011: color_data = Z;
		19'b0011100010011010100: color_data = Z;
		19'b0011100010011010101: color_data = Z;
		19'b0011100010011010110: color_data = Z;
		19'b0011100010011010111: color_data = Z;
		19'b0011100010011011000: color_data = Z;
		19'b0011100010011011001: color_data = Z;
		19'b0011100010011011010: color_data = Z;
		19'b0011100010011011011: color_data = Z;
		19'b0011100010011011100: color_data = Z;
		19'b0011100010011011101: color_data = Z;
		19'b0011100010011011110: color_data = Z;
		19'b0011100010011011111: color_data = Z;
		19'b0011100010011100000: color_data = Z;
		19'b0011100010011100001: color_data = Z;
		19'b0011100010011100010: color_data = Z;
		19'b0011100010011100011: color_data = Z;
		19'b0011100010011100100: color_data = Z;
		19'b0011100010011100101: color_data = Z;
		19'b0011100010011100110: color_data = Z;
		19'b0011100010011100111: color_data = Z;
		19'b0011100010011101000: color_data = Z;
		19'b0011100010011101001: color_data = Z;
		19'b0011100010011101010: color_data = Z;
		19'b0011100010011101011: color_data = Z;
		19'b0011100010011101100: color_data = Z;
		19'b0011100010011101101: color_data = Z;
		19'b0011100010011101110: color_data = Z;
		19'b0011100010011101111: color_data = Z;
		19'b0011100010011110000: color_data = Z;
		19'b0011100010011110001: color_data = Z;
		19'b0011100010011110010: color_data = Z;
		19'b0011100010011110011: color_data = Z;
		19'b0011100010011110100: color_data = Z;
		19'b0011100010011110101: color_data = Z;
		19'b0011100010011110110: color_data = Z;
		19'b0011100010011110111: color_data = Z;
		19'b0011100010011111000: color_data = Z;
		19'b0011100010011111001: color_data = Z;
		19'b0011100010011111010: color_data = Z;
		19'b0011100010011111011: color_data = Z;
		19'b0011100010011111100: color_data = Z;
		19'b0011100010011111101: color_data = Z;
		19'b0011100010011111110: color_data = Z;
		19'b0011100010011111111: color_data = Z;
		19'b0011100010100000000: color_data = Z;
		19'b0011100010100000001: color_data = Z;
		19'b0011100010100000010: color_data = Z;
		19'b0011100010100000011: color_data = Z;
		19'b0011100010100000100: color_data = Z;
		19'b0011100010100000101: color_data = Z;
		19'b0011100010100000110: color_data = Z;
		19'b0011100010100000111: color_data = Z;
		19'b0011100010100001000: color_data = Z;
		19'b0011100010100001001: color_data = Z;
		19'b0011100010100001010: color_data = Z;
		19'b0011100010100001011: color_data = Z;
		19'b0011100010100001100: color_data = Z;
		19'b0011100010100001101: color_data = Z;
		19'b0011100010100001110: color_data = Z;
		19'b0011100010100001111: color_data = Z;
		19'b0011100010100010000: color_data = Z;
		19'b0011100010100010001: color_data = Z;
		19'b0011100010100010010: color_data = Z;
		19'b0011100010100010011: color_data = Z;
		19'b0011100010100010100: color_data = Z;
		19'b0011100010100010101: color_data = Z;
		19'b0011100010100010110: color_data = Z;
		19'b0011100010100010111: color_data = Z;
		19'b0011100010100011000: color_data = Z;
		19'b0011100010100011001: color_data = Z;
		19'b0011100010100011010: color_data = Z;
		19'b0011100010100011011: color_data = Z;
		19'b0011100010100011100: color_data = Z;
		19'b0011100010100011101: color_data = Z;
		19'b0011100010100011110: color_data = Z;
		19'b0011100010100011111: color_data = Z;
		19'b0011100010100100000: color_data = Z;
		19'b0011100010100100001: color_data = Z;
		19'b0011100010100100010: color_data = Z;
		19'b0011100010100100011: color_data = Z;
		19'b0011100010100100100: color_data = Z;
		19'b0011100010100100101: color_data = Z;
		19'b0011100010100100110: color_data = Z;
		19'b0011100010100100111: color_data = Z;
		19'b0011100010100101000: color_data = Z;
		19'b0011100010100101001: color_data = Z;
		19'b0011100010100101010: color_data = Z;
		19'b0011100010100101011: color_data = Z;
		19'b0011100010100101100: color_data = Z;
		19'b0011100010100101101: color_data = Z;
		19'b0011100010100101110: color_data = Z;
		19'b0011100010100101111: color_data = Z;
		19'b0011100010100110000: color_data = Z;
		19'b0011100010100110001: color_data = Z;
		19'b0011100010100110010: color_data = Z;
		19'b0011100010100110011: color_data = Z;
		19'b0011100010100110100: color_data = Z;
		19'b0011100010100110101: color_data = Z;
		19'b0011100010100110110: color_data = Z;
		19'b0011100010100110111: color_data = Z;
		19'b0011100010100111000: color_data = Z;
		19'b0011100010100111001: color_data = Z;
		19'b0011100010100111010: color_data = Z;
		19'b0011100010100111011: color_data = Z;
		19'b0011100010100111100: color_data = Z;
		19'b0011100010100111101: color_data = Z;
		19'b0011100010100111110: color_data = Z;
		19'b0011100010100111111: color_data = Z;
		19'b0011100010101000000: color_data = Z;
		19'b0011100010101000001: color_data = Z;
		19'b0011100010101000010: color_data = Z;
		19'b0011100010101000011: color_data = Z;
		19'b0011100010101000100: color_data = Z;
		19'b0011100010101000101: color_data = Z;
		19'b0011100010101000110: color_data = Z;
		19'b0011100010101000111: color_data = Z;
		19'b0011100010101001000: color_data = Z;
		19'b0011100010101001001: color_data = Z;
		19'b0011100010101001010: color_data = Z;
		19'b0011100010101001011: color_data = Z;
		19'b0011100010101001100: color_data = Z;
		19'b0011100010101001101: color_data = Z;
		19'b0011100010101001110: color_data = Z;
		19'b0011100010101001111: color_data = Z;
		19'b0011100010101010000: color_data = Z;
		19'b0011100010101010001: color_data = Z;
		19'b0011100010101010010: color_data = Z;
		19'b0011100010101010011: color_data = Z;
		19'b0011100010101010100: color_data = Z;
		19'b0011100010101010101: color_data = Z;
		19'b0011100010101010110: color_data = Z;
		19'b0011100010101010111: color_data = Z;
		19'b0011100010101011000: color_data = Z;
		19'b0011100010101011001: color_data = Z;
		19'b0011100010101011010: color_data = Z;
		19'b0011100010101011011: color_data = Z;
		19'b0011100010101011100: color_data = Z;
		19'b0011100010101011101: color_data = Z;
		19'b0011100010101011110: color_data = Z;
		19'b0011100010101011111: color_data = Z;
		19'b0011100010101100000: color_data = Z;
		19'b0011100010101100001: color_data = Z;
		19'b0011100010101100010: color_data = Z;
		19'b0011100010101100011: color_data = Z;
		19'b0011100010101100100: color_data = Z;
		19'b0011100010101100101: color_data = Z;
		19'b0011100010101100110: color_data = Z;
		19'b0011100010101100111: color_data = Z;
		19'b0011100010101101000: color_data = Z;
		19'b0011100010101101001: color_data = Z;
		19'b0011100010101101010: color_data = Z;
		19'b0011100010101101011: color_data = Z;
		19'b0011100010101101100: color_data = Z;
		19'b0011100010101101101: color_data = Z;
		19'b0011100010101101110: color_data = Z;
		19'b0011100010101101111: color_data = Z;
		19'b0011100010101110000: color_data = Z;
		19'b0011100010101110001: color_data = Z;
		19'b0011100010101110010: color_data = Z;
		19'b0011100010101110011: color_data = Z;
		19'b0011100010101110100: color_data = Z;
		19'b0011100010101110101: color_data = Z;
		19'b0011100010101110110: color_data = Z;
		19'b0011100010101110111: color_data = Z;
		19'b0011100010101111000: color_data = Z;
		19'b0011100010101111001: color_data = Z;
		19'b0011100010101111010: color_data = Z;
		19'b0011100010101111011: color_data = Z;
		19'b0011100010101111100: color_data = Z;
		19'b0011100010101111101: color_data = Z;
		19'b0011100010101111110: color_data = Z;
		19'b0011100010101111111: color_data = Z;
		19'b0011100010110000000: color_data = Z;
		19'b0011100010110000001: color_data = Z;
		19'b0011100010110000010: color_data = Z;
		19'b0011100010110000011: color_data = Z;
		19'b0011100010110000100: color_data = Z;
		19'b0011100010110000101: color_data = Z;
		19'b0011100010110000110: color_data = Z;
		19'b0011100010110000111: color_data = Z;
		19'b0011100010110001000: color_data = Z;
		19'b0011100010110001001: color_data = Z;
		19'b0011100010110001010: color_data = Z;
		19'b0011100010110001011: color_data = Z;
		19'b0011100010110001100: color_data = Z;
		19'b0011100010110001101: color_data = Z;
		19'b0011100010110001110: color_data = Z;
		19'b0011100010110001111: color_data = Z;
		19'b0011100010110010000: color_data = Z;
		19'b0011100010110010001: color_data = Z;
		19'b0011100010110010010: color_data = Z;
		19'b0011100010110111010: color_data = Z;
		19'b0011100010110111011: color_data = Z;
		19'b0011100010110111100: color_data = Z;
		19'b0011100010110111101: color_data = Z;
		19'b0011100010110111110: color_data = Z;
		19'b0011100010110111111: color_data = Z;
		19'b0011100010111000000: color_data = Z;
		19'b0011100010111011101: color_data = Z;
		19'b0011100100010101110: color_data = Z;
		19'b0011100100010101111: color_data = Z;
		19'b0011100100010110100: color_data = Z;
		19'b0011100100010110101: color_data = Z;
		19'b0011100100010110110: color_data = Z;
		19'b0011100100010110111: color_data = Z;
		19'b0011100100010111000: color_data = Z;
		19'b0011100100010111001: color_data = Z;
		19'b0011100100010111010: color_data = Z;
		19'b0011100100010111011: color_data = Z;
		19'b0011100100010111100: color_data = Z;
		19'b0011100100010111101: color_data = Z;
		19'b0011100100010111110: color_data = Z;
		19'b0011100100010111111: color_data = Z;
		19'b0011100100011000000: color_data = Z;
		19'b0011100100011000001: color_data = Z;
		19'b0011100100011000010: color_data = Z;
		19'b0011100100011000011: color_data = Z;
		19'b0011100100011000100: color_data = Z;
		19'b0011100100011000101: color_data = Z;
		19'b0011100100011000110: color_data = Z;
		19'b0011100100011000111: color_data = Z;
		19'b0011100100011001000: color_data = Z;
		19'b0011100100011001001: color_data = Z;
		19'b0011100100011001010: color_data = Z;
		19'b0011100100011001011: color_data = Z;
		19'b0011100100011001100: color_data = Z;
		19'b0011100100011001101: color_data = Z;
		19'b0011100100011001110: color_data = Z;
		19'b0011100100011001111: color_data = Z;
		19'b0011100100011010000: color_data = Z;
		19'b0011100100011010001: color_data = Z;
		19'b0011100100011010010: color_data = Z;
		19'b0011100100011010011: color_data = Z;
		19'b0011100100011010100: color_data = Z;
		19'b0011100100011010101: color_data = Z;
		19'b0011100100011010110: color_data = Z;
		19'b0011100100011010111: color_data = Z;
		19'b0011100100011011000: color_data = Z;
		19'b0011100100011011001: color_data = Z;
		19'b0011100100011011010: color_data = Z;
		19'b0011100100011011011: color_data = Z;
		19'b0011100100011011100: color_data = Z;
		19'b0011100100011011101: color_data = Z;
		19'b0011100100011011110: color_data = Z;
		19'b0011100100011011111: color_data = Z;
		19'b0011100100011100000: color_data = Z;
		19'b0011100100011100001: color_data = Z;
		19'b0011100100011100010: color_data = Z;
		19'b0011100100011100011: color_data = Z;
		19'b0011100100011100100: color_data = Z;
		19'b0011100100011100101: color_data = Z;
		19'b0011100100011100110: color_data = Z;
		19'b0011100100011100111: color_data = Z;
		19'b0011100100011101000: color_data = Z;
		19'b0011100100011101001: color_data = Z;
		19'b0011100100011101010: color_data = Z;
		19'b0011100100011101011: color_data = Z;
		19'b0011100100011101100: color_data = Z;
		19'b0011100100011101101: color_data = Z;
		19'b0011100100011101110: color_data = Z;
		19'b0011100100011101111: color_data = Z;
		19'b0011100100011110000: color_data = Z;
		19'b0011100100011110001: color_data = Z;
		19'b0011100100011110010: color_data = Z;
		19'b0011100100011110011: color_data = Z;
		19'b0011100100011110100: color_data = Z;
		19'b0011100100011110101: color_data = Z;
		19'b0011100100011110110: color_data = Z;
		19'b0011100100011110111: color_data = Z;
		19'b0011100100011111000: color_data = Z;
		19'b0011100100011111001: color_data = Z;
		19'b0011100100011111010: color_data = Z;
		19'b0011100100011111011: color_data = Z;
		19'b0011100100011111100: color_data = Z;
		19'b0011100100011111101: color_data = Z;
		19'b0011100100011111110: color_data = Z;
		19'b0011100100011111111: color_data = Z;
		19'b0011100100100000000: color_data = Z;
		19'b0011100100100000001: color_data = Z;
		19'b0011100100100000010: color_data = Z;
		19'b0011100100100000011: color_data = Z;
		19'b0011100100100000100: color_data = Z;
		19'b0011100100100000101: color_data = Z;
		19'b0011100100100000110: color_data = Z;
		19'b0011100100100000111: color_data = Z;
		19'b0011100100100001000: color_data = Z;
		19'b0011100100100001001: color_data = Z;
		19'b0011100100100001010: color_data = Z;
		19'b0011100100100001011: color_data = Z;
		19'b0011100100100001100: color_data = Z;
		19'b0011100100100001101: color_data = Z;
		19'b0011100100100001110: color_data = Z;
		19'b0011100100100001111: color_data = Z;
		19'b0011100100100010000: color_data = Z;
		19'b0011100100100010001: color_data = Z;
		19'b0011100100100010010: color_data = Z;
		19'b0011100100100010011: color_data = Z;
		19'b0011100100100010100: color_data = Z;
		19'b0011100100100010101: color_data = Z;
		19'b0011100100100010110: color_data = Z;
		19'b0011100100100010111: color_data = Z;
		19'b0011100100100011000: color_data = Z;
		19'b0011100100100011001: color_data = Z;
		19'b0011100100100011010: color_data = Z;
		19'b0011100100100011011: color_data = Z;
		19'b0011100100100011100: color_data = Z;
		19'b0011100100100011101: color_data = Z;
		19'b0011100100100011110: color_data = Z;
		19'b0011100100100011111: color_data = Z;
		19'b0011100100100100000: color_data = Z;
		19'b0011100100100100001: color_data = Z;
		19'b0011100100100100010: color_data = Z;
		19'b0011100100100100011: color_data = Z;
		19'b0011100100100100100: color_data = Z;
		19'b0011100100100100101: color_data = Z;
		19'b0011100100100100110: color_data = Z;
		19'b0011100100100100111: color_data = Z;
		19'b0011100100100101000: color_data = Z;
		19'b0011100100100101001: color_data = Z;
		19'b0011100100100101010: color_data = Z;
		19'b0011100100100101011: color_data = Z;
		19'b0011100100100101100: color_data = Z;
		19'b0011100100100101101: color_data = Z;
		19'b0011100100100101110: color_data = Z;
		19'b0011100100100101111: color_data = Z;
		19'b0011100100100110000: color_data = Z;
		19'b0011100100100110001: color_data = Z;
		19'b0011100100100110010: color_data = Z;
		19'b0011100100100110011: color_data = Z;
		19'b0011100100100110100: color_data = Z;
		19'b0011100100100110101: color_data = Z;
		19'b0011100100100110110: color_data = Z;
		19'b0011100100100110111: color_data = Z;
		19'b0011100100100111000: color_data = Z;
		19'b0011100100100111001: color_data = Z;
		19'b0011100100100111010: color_data = Z;
		19'b0011100100100111011: color_data = Z;
		19'b0011100100100111100: color_data = Z;
		19'b0011100100100111101: color_data = Z;
		19'b0011100100100111110: color_data = Z;
		19'b0011100100100111111: color_data = Z;
		19'b0011100100101000000: color_data = Z;
		19'b0011100100101000001: color_data = Z;
		19'b0011100100101000010: color_data = Z;
		19'b0011100100101000011: color_data = Z;
		19'b0011100100101000100: color_data = Z;
		19'b0011100100101000101: color_data = Z;
		19'b0011100100101000110: color_data = Z;
		19'b0011100100101000111: color_data = Z;
		19'b0011100100101001000: color_data = Z;
		19'b0011100100101001001: color_data = Z;
		19'b0011100100101001010: color_data = Z;
		19'b0011100100101001011: color_data = Z;
		19'b0011100100101001100: color_data = Z;
		19'b0011100100101001101: color_data = Z;
		19'b0011100100101001110: color_data = Z;
		19'b0011100100101001111: color_data = Z;
		19'b0011100100101010000: color_data = Z;
		19'b0011100100101010001: color_data = Z;
		19'b0011100100101010010: color_data = Z;
		19'b0011100100101010011: color_data = Z;
		19'b0011100100101010100: color_data = Z;
		19'b0011100100101010101: color_data = Z;
		19'b0011100100101010110: color_data = Z;
		19'b0011100100101010111: color_data = Z;
		19'b0011100100101011000: color_data = Z;
		19'b0011100100101011001: color_data = Z;
		19'b0011100100101011010: color_data = Z;
		19'b0011100100101011011: color_data = Z;
		19'b0011100100101011100: color_data = Z;
		19'b0011100100101011101: color_data = Z;
		19'b0011100100101011110: color_data = Z;
		19'b0011100100101011111: color_data = Z;
		19'b0011100100101100000: color_data = Z;
		19'b0011100100101100001: color_data = Z;
		19'b0011100100101100010: color_data = Z;
		19'b0011100100101100011: color_data = Z;
		19'b0011100100101100100: color_data = Z;
		19'b0011100100101100101: color_data = Z;
		19'b0011100100101100110: color_data = Z;
		19'b0011100100101100111: color_data = Z;
		19'b0011100100101101000: color_data = Z;
		19'b0011100100101101001: color_data = Z;
		19'b0011100100101101010: color_data = Z;
		19'b0011100100101101011: color_data = Z;
		19'b0011100100101101100: color_data = Z;
		19'b0011100100101101101: color_data = Z;
		19'b0011100100101101110: color_data = Z;
		19'b0011100100101101111: color_data = Z;
		19'b0011100100101110000: color_data = Z;
		19'b0011100100101110001: color_data = Z;
		19'b0011100100101110010: color_data = Z;
		19'b0011100100101110011: color_data = Z;
		19'b0011100100101110100: color_data = Z;
		19'b0011100100101110101: color_data = Z;
		19'b0011100100101110110: color_data = Z;
		19'b0011100100101110111: color_data = Z;
		19'b0011100100101111000: color_data = Z;
		19'b0011100100101111001: color_data = Z;
		19'b0011100100101111010: color_data = Z;
		19'b0011100100101111011: color_data = Z;
		19'b0011100100101111100: color_data = Z;
		19'b0011100100101111101: color_data = Z;
		19'b0011100100101111110: color_data = Z;
		19'b0011100100101111111: color_data = Z;
		19'b0011100100110000000: color_data = Z;
		19'b0011100100110000001: color_data = Z;
		19'b0011100100110000010: color_data = Z;
		19'b0011100100110000011: color_data = Z;
		19'b0011100100110000100: color_data = Z;
		19'b0011100100110000101: color_data = Z;
		19'b0011100100110000110: color_data = Z;
		19'b0011100100110000111: color_data = Z;
		19'b0011100100110001000: color_data = Z;
		19'b0011100100110001001: color_data = Z;
		19'b0011100100110001010: color_data = Z;
		19'b0011100100110001011: color_data = Z;
		19'b0011100100110001100: color_data = Z;
		19'b0011100100110001101: color_data = Z;
		19'b0011100100110001110: color_data = Z;
		19'b0011100100110001111: color_data = Z;
		19'b0011100100110010000: color_data = Z;
		19'b0011100100110010001: color_data = Z;
		19'b0011100100110010010: color_data = Z;
		19'b0011100100110111011: color_data = Z;
		19'b0011100100110111100: color_data = Z;
		19'b0011100100110111101: color_data = Z;
		19'b0011100100110111110: color_data = Z;
		19'b0011100100110111111: color_data = Z;
		19'b0011100100111000000: color_data = Z;
		19'b0011100100111000001: color_data = Z;
		19'b0011100100111011101: color_data = Z;
		19'b0011100110010110100: color_data = Z;
		19'b0011100110010110101: color_data = Z;
		19'b0011100110010110110: color_data = Z;
		19'b0011100110010110111: color_data = Z;
		19'b0011100110010111000: color_data = Z;
		19'b0011100110010111001: color_data = Z;
		19'b0011100110010111010: color_data = Z;
		19'b0011100110010111011: color_data = Z;
		19'b0011100110010111100: color_data = Z;
		19'b0011100110010111101: color_data = Z;
		19'b0011100110010111110: color_data = Z;
		19'b0011100110010111111: color_data = Z;
		19'b0011100110011000000: color_data = Z;
		19'b0011100110011000001: color_data = Z;
		19'b0011100110011000010: color_data = Z;
		19'b0011100110011000011: color_data = Z;
		19'b0011100110011000100: color_data = Z;
		19'b0011100110011000101: color_data = Z;
		19'b0011100110011000110: color_data = Z;
		19'b0011100110011000111: color_data = Z;
		19'b0011100110011001000: color_data = Z;
		19'b0011100110011001001: color_data = Z;
		19'b0011100110011001010: color_data = Z;
		19'b0011100110011001011: color_data = Z;
		19'b0011100110011001100: color_data = Z;
		19'b0011100110011001101: color_data = Z;
		19'b0011100110011001110: color_data = Z;
		19'b0011100110011001111: color_data = Z;
		19'b0011100110011010000: color_data = Z;
		19'b0011100110011010001: color_data = Z;
		19'b0011100110011010010: color_data = Z;
		19'b0011100110011010011: color_data = Z;
		19'b0011100110011010100: color_data = Z;
		19'b0011100110011010101: color_data = Z;
		19'b0011100110011010110: color_data = Z;
		19'b0011100110011010111: color_data = Z;
		19'b0011100110011011000: color_data = Z;
		19'b0011100110011011001: color_data = Z;
		19'b0011100110011011010: color_data = Z;
		19'b0011100110011011011: color_data = Z;
		19'b0011100110011011100: color_data = Z;
		19'b0011100110011011101: color_data = Z;
		19'b0011100110011011110: color_data = Z;
		19'b0011100110011011111: color_data = Z;
		19'b0011100110011100000: color_data = Z;
		19'b0011100110011100001: color_data = Z;
		19'b0011100110011100010: color_data = Z;
		19'b0011100110011100011: color_data = Z;
		19'b0011100110011100100: color_data = Z;
		19'b0011100110011100101: color_data = Z;
		19'b0011100110011100110: color_data = Z;
		19'b0011100110011100111: color_data = Z;
		19'b0011100110011101000: color_data = Z;
		19'b0011100110011101001: color_data = Z;
		19'b0011100110011101010: color_data = Z;
		19'b0011100110011101011: color_data = Z;
		19'b0011100110011101100: color_data = Z;
		19'b0011100110011101101: color_data = Z;
		19'b0011100110011101110: color_data = Z;
		19'b0011100110011101111: color_data = Z;
		19'b0011100110011110000: color_data = Z;
		19'b0011100110011110001: color_data = Z;
		19'b0011100110011110010: color_data = Z;
		19'b0011100110011110011: color_data = Z;
		19'b0011100110011110100: color_data = Z;
		19'b0011100110011110101: color_data = Z;
		19'b0011100110011110110: color_data = Z;
		19'b0011100110011110111: color_data = Z;
		19'b0011100110011111000: color_data = Z;
		19'b0011100110011111001: color_data = Z;
		19'b0011100110011111010: color_data = Z;
		19'b0011100110011111011: color_data = Z;
		19'b0011100110011111100: color_data = Z;
		19'b0011100110011111101: color_data = Z;
		19'b0011100110011111110: color_data = Z;
		19'b0011100110011111111: color_data = Z;
		19'b0011100110100000000: color_data = Z;
		19'b0011100110100000001: color_data = Z;
		19'b0011100110100000010: color_data = Z;
		19'b0011100110100000011: color_data = Z;
		19'b0011100110100000100: color_data = Z;
		19'b0011100110100000101: color_data = Z;
		19'b0011100110100000110: color_data = Z;
		19'b0011100110100000111: color_data = Z;
		19'b0011100110100001000: color_data = Z;
		19'b0011100110100001001: color_data = Z;
		19'b0011100110100001010: color_data = Z;
		19'b0011100110100001011: color_data = Z;
		19'b0011100110100001100: color_data = Z;
		19'b0011100110100001101: color_data = Z;
		19'b0011100110100001110: color_data = Z;
		19'b0011100110100001111: color_data = Z;
		19'b0011100110100010000: color_data = Z;
		19'b0011100110100010001: color_data = Z;
		19'b0011100110100010010: color_data = Z;
		19'b0011100110100010011: color_data = Z;
		19'b0011100110100010100: color_data = Z;
		19'b0011100110100010101: color_data = Z;
		19'b0011100110100010110: color_data = Z;
		19'b0011100110100010111: color_data = Z;
		19'b0011100110100011000: color_data = Z;
		19'b0011100110100011001: color_data = Z;
		19'b0011100110100011010: color_data = Z;
		19'b0011100110100011011: color_data = Z;
		19'b0011100110100011100: color_data = Z;
		19'b0011100110100011101: color_data = Z;
		19'b0011100110100011110: color_data = Z;
		19'b0011100110100011111: color_data = Z;
		19'b0011100110100100000: color_data = Z;
		19'b0011100110100100001: color_data = Z;
		19'b0011100110100100010: color_data = Z;
		19'b0011100110100100011: color_data = Z;
		19'b0011100110100100100: color_data = Z;
		19'b0011100110100100101: color_data = Z;
		19'b0011100110100100110: color_data = Z;
		19'b0011100110100100111: color_data = Z;
		19'b0011100110100101000: color_data = Z;
		19'b0011100110100101001: color_data = Z;
		19'b0011100110100101010: color_data = Z;
		19'b0011100110100101011: color_data = Z;
		19'b0011100110100101100: color_data = Z;
		19'b0011100110100101101: color_data = Z;
		19'b0011100110100101110: color_data = Z;
		19'b0011100110100101111: color_data = Z;
		19'b0011100110100110000: color_data = Z;
		19'b0011100110100110001: color_data = Z;
		19'b0011100110100110010: color_data = Z;
		19'b0011100110100110011: color_data = Z;
		19'b0011100110100110100: color_data = Z;
		19'b0011100110100110101: color_data = Z;
		19'b0011100110100110110: color_data = Z;
		19'b0011100110100110111: color_data = Z;
		19'b0011100110100111000: color_data = Z;
		19'b0011100110100111001: color_data = Z;
		19'b0011100110100111010: color_data = Z;
		19'b0011100110100111011: color_data = Z;
		19'b0011100110100111100: color_data = Z;
		19'b0011100110100111101: color_data = Z;
		19'b0011100110100111110: color_data = Z;
		19'b0011100110100111111: color_data = Z;
		19'b0011100110101000000: color_data = Z;
		19'b0011100110101000001: color_data = Z;
		19'b0011100110101000010: color_data = Z;
		19'b0011100110101000011: color_data = Z;
		19'b0011100110101000100: color_data = Z;
		19'b0011100110101000101: color_data = Z;
		19'b0011100110101000110: color_data = Z;
		19'b0011100110101000111: color_data = Z;
		19'b0011100110101001000: color_data = Z;
		19'b0011100110101001001: color_data = Z;
		19'b0011100110101001010: color_data = Z;
		19'b0011100110101001011: color_data = Z;
		19'b0011100110101001100: color_data = Z;
		19'b0011100110101001101: color_data = Z;
		19'b0011100110101001110: color_data = Z;
		19'b0011100110101001111: color_data = Z;
		19'b0011100110101010000: color_data = Z;
		19'b0011100110101010001: color_data = Z;
		19'b0011100110101010010: color_data = Z;
		19'b0011100110101010011: color_data = Z;
		19'b0011100110101010100: color_data = Z;
		19'b0011100110101010101: color_data = Z;
		19'b0011100110101010110: color_data = Z;
		19'b0011100110101010111: color_data = Z;
		19'b0011100110101011000: color_data = Z;
		19'b0011100110101011001: color_data = Z;
		19'b0011100110101011010: color_data = Z;
		19'b0011100110101011011: color_data = Z;
		19'b0011100110101011100: color_data = Z;
		19'b0011100110101011101: color_data = Z;
		19'b0011100110101011110: color_data = Z;
		19'b0011100110101011111: color_data = Z;
		19'b0011100110101100000: color_data = Z;
		19'b0011100110101100001: color_data = Z;
		19'b0011100110101100010: color_data = Z;
		19'b0011100110101100011: color_data = Z;
		19'b0011100110101100100: color_data = Z;
		19'b0011100110101100101: color_data = Z;
		19'b0011100110101100110: color_data = Z;
		19'b0011100110101100111: color_data = Z;
		19'b0011100110101101000: color_data = Z;
		19'b0011100110101101001: color_data = Z;
		19'b0011100110101101010: color_data = Z;
		19'b0011100110101101011: color_data = Z;
		19'b0011100110101101100: color_data = Z;
		19'b0011100110101101101: color_data = Z;
		19'b0011100110101101110: color_data = Z;
		19'b0011100110101101111: color_data = Z;
		19'b0011100110101110000: color_data = Z;
		19'b0011100110101110001: color_data = Z;
		19'b0011100110101110010: color_data = Z;
		19'b0011100110101110011: color_data = Z;
		19'b0011100110101110100: color_data = Z;
		19'b0011100110101110101: color_data = Z;
		19'b0011100110101110110: color_data = Z;
		19'b0011100110101110111: color_data = Z;
		19'b0011100110101111000: color_data = Z;
		19'b0011100110101111001: color_data = Z;
		19'b0011100110101111010: color_data = Z;
		19'b0011100110101111011: color_data = Z;
		19'b0011100110101111100: color_data = Z;
		19'b0011100110101111101: color_data = Z;
		19'b0011100110101111110: color_data = Z;
		19'b0011100110101111111: color_data = Z;
		19'b0011100110110000000: color_data = Z;
		19'b0011100110110000001: color_data = Z;
		19'b0011100110110000010: color_data = Z;
		19'b0011100110110000011: color_data = Z;
		19'b0011100110110000100: color_data = Z;
		19'b0011100110110000101: color_data = Z;
		19'b0011100110110000110: color_data = Z;
		19'b0011100110110000111: color_data = Z;
		19'b0011100110110001000: color_data = Z;
		19'b0011100110110001001: color_data = Z;
		19'b0011100110110001010: color_data = Z;
		19'b0011100110110001011: color_data = Z;
		19'b0011100110110001100: color_data = Z;
		19'b0011100110110001101: color_data = Z;
		19'b0011100110110001110: color_data = Z;
		19'b0011100110110001111: color_data = Z;
		19'b0011100110110010000: color_data = Z;
		19'b0011100110110010001: color_data = Z;
		19'b0011100110110111011: color_data = Z;
		19'b0011100110110111100: color_data = Z;
		19'b0011100110110111101: color_data = Z;
		19'b0011100110110111110: color_data = Z;
		19'b0011100110110111111: color_data = Z;
		19'b0011100110111000000: color_data = Z;
		19'b0011100110111000001: color_data = Z;
		19'b0011100110111000010: color_data = Z;
		19'b0011100110111000100: color_data = Z;
		19'b0011100110111000101: color_data = Z;
		19'b0011101000010110011: color_data = Z;
		19'b0011101000010110100: color_data = Z;
		19'b0011101000010110101: color_data = Z;
		19'b0011101000010110110: color_data = Z;
		19'b0011101000010110111: color_data = Z;
		19'b0011101000010111000: color_data = Z;
		19'b0011101000010111001: color_data = Z;
		19'b0011101000010111010: color_data = Z;
		19'b0011101000010111011: color_data = Z;
		19'b0011101000010111100: color_data = Z;
		19'b0011101000010111101: color_data = Z;
		19'b0011101000010111110: color_data = Z;
		19'b0011101000010111111: color_data = Z;
		19'b0011101000011000000: color_data = Z;
		19'b0011101000011000001: color_data = Z;
		19'b0011101000011000010: color_data = Z;
		19'b0011101000011000011: color_data = Z;
		19'b0011101000011000100: color_data = Z;
		19'b0011101000011000101: color_data = Z;
		19'b0011101000011000110: color_data = Z;
		19'b0011101000011000111: color_data = Z;
		19'b0011101000011001000: color_data = Z;
		19'b0011101000011001001: color_data = Z;
		19'b0011101000011001010: color_data = Z;
		19'b0011101000011001011: color_data = Z;
		19'b0011101000011001100: color_data = Z;
		19'b0011101000011001101: color_data = Z;
		19'b0011101000011001110: color_data = Z;
		19'b0011101000011001111: color_data = Z;
		19'b0011101000011010000: color_data = Z;
		19'b0011101000011010001: color_data = Z;
		19'b0011101000011010010: color_data = Z;
		19'b0011101000011010011: color_data = Z;
		19'b0011101000011010100: color_data = Z;
		19'b0011101000011010101: color_data = Z;
		19'b0011101000011010110: color_data = Z;
		19'b0011101000011010111: color_data = Z;
		19'b0011101000011011000: color_data = Z;
		19'b0011101000011011001: color_data = Z;
		19'b0011101000011011010: color_data = Z;
		19'b0011101000011011011: color_data = Z;
		19'b0011101000011011100: color_data = Z;
		19'b0011101000011011101: color_data = Z;
		19'b0011101000011011110: color_data = Z;
		19'b0011101000011011111: color_data = Z;
		19'b0011101000011100000: color_data = Z;
		19'b0011101000011100001: color_data = Z;
		19'b0011101000011100010: color_data = Z;
		19'b0011101000011100011: color_data = Z;
		19'b0011101000011100100: color_data = Z;
		19'b0011101000011100101: color_data = Z;
		19'b0011101000011100110: color_data = Z;
		19'b0011101000011100111: color_data = Z;
		19'b0011101000011101000: color_data = Z;
		19'b0011101000011101001: color_data = Z;
		19'b0011101000011101010: color_data = Z;
		19'b0011101000011101011: color_data = Z;
		19'b0011101000011101100: color_data = Z;
		19'b0011101000011101101: color_data = Z;
		19'b0011101000011101110: color_data = Z;
		19'b0011101000011101111: color_data = Z;
		19'b0011101000011110000: color_data = Z;
		19'b0011101000011110001: color_data = Z;
		19'b0011101000011110010: color_data = Z;
		19'b0011101000011110011: color_data = Z;
		19'b0011101000011110100: color_data = Z;
		19'b0011101000011110101: color_data = Z;
		19'b0011101000011110110: color_data = Z;
		19'b0011101000011110111: color_data = Z;
		19'b0011101000011111000: color_data = Z;
		19'b0011101000011111001: color_data = Z;
		19'b0011101000011111010: color_data = Z;
		19'b0011101000011111011: color_data = Z;
		19'b0011101000011111100: color_data = Z;
		19'b0011101000011111101: color_data = Z;
		19'b0011101000011111110: color_data = Z;
		19'b0011101000011111111: color_data = Z;
		19'b0011101000100000000: color_data = Z;
		19'b0011101000100000001: color_data = Z;
		19'b0011101000100000010: color_data = Z;
		19'b0011101000100000011: color_data = Z;
		19'b0011101000100000100: color_data = Z;
		19'b0011101000100000101: color_data = Z;
		19'b0011101000100000110: color_data = Z;
		19'b0011101000100000111: color_data = Z;
		19'b0011101000100001000: color_data = Z;
		19'b0011101000100001001: color_data = Z;
		19'b0011101000100001010: color_data = Z;
		19'b0011101000100001011: color_data = Z;
		19'b0011101000100001100: color_data = Z;
		19'b0011101000100001101: color_data = Z;
		19'b0011101000100001110: color_data = Z;
		19'b0011101000100001111: color_data = Z;
		19'b0011101000100010000: color_data = Z;
		19'b0011101000100010001: color_data = Z;
		19'b0011101000100010010: color_data = Z;
		19'b0011101000100010011: color_data = Z;
		19'b0011101000100010100: color_data = Z;
		19'b0011101000100010101: color_data = Z;
		19'b0011101000100010110: color_data = Z;
		19'b0011101000100010111: color_data = Z;
		19'b0011101000100011000: color_data = Z;
		19'b0011101000100011001: color_data = Z;
		19'b0011101000100011010: color_data = Z;
		19'b0011101000100011011: color_data = Z;
		19'b0011101000100011100: color_data = Z;
		19'b0011101000100011101: color_data = Z;
		19'b0011101000100011110: color_data = Z;
		19'b0011101000100011111: color_data = Z;
		19'b0011101000100100000: color_data = Z;
		19'b0011101000100100001: color_data = Z;
		19'b0011101000100100010: color_data = Z;
		19'b0011101000100100011: color_data = Z;
		19'b0011101000100100100: color_data = Z;
		19'b0011101000100100101: color_data = Z;
		19'b0011101000100100110: color_data = Z;
		19'b0011101000100100111: color_data = Z;
		19'b0011101000100101000: color_data = Z;
		19'b0011101000100101001: color_data = Z;
		19'b0011101000100101010: color_data = Z;
		19'b0011101000100101011: color_data = Z;
		19'b0011101000100101100: color_data = Z;
		19'b0011101000100101101: color_data = Z;
		19'b0011101000100101110: color_data = Z;
		19'b0011101000100101111: color_data = Z;
		19'b0011101000100110000: color_data = Z;
		19'b0011101000100110001: color_data = Z;
		19'b0011101000100110010: color_data = Z;
		19'b0011101000100110011: color_data = Z;
		19'b0011101000100110100: color_data = Z;
		19'b0011101000100110101: color_data = Z;
		19'b0011101000100110110: color_data = Z;
		19'b0011101000100110111: color_data = Z;
		19'b0011101000100111000: color_data = Z;
		19'b0011101000100111001: color_data = Z;
		19'b0011101000100111010: color_data = Z;
		19'b0011101000100111011: color_data = Z;
		19'b0011101000100111100: color_data = Z;
		19'b0011101000100111101: color_data = Z;
		19'b0011101000100111110: color_data = Z;
		19'b0011101000100111111: color_data = Z;
		19'b0011101000101000000: color_data = Z;
		19'b0011101000101000001: color_data = Z;
		19'b0011101000101000010: color_data = Z;
		19'b0011101000101000011: color_data = Z;
		19'b0011101000101000100: color_data = Z;
		19'b0011101000101000101: color_data = Z;
		19'b0011101000101000110: color_data = Z;
		19'b0011101000101000111: color_data = Z;
		19'b0011101000101001000: color_data = Z;
		19'b0011101000101001001: color_data = Z;
		19'b0011101000101001010: color_data = Z;
		19'b0011101000101001011: color_data = Z;
		19'b0011101000101001100: color_data = Z;
		19'b0011101000101001101: color_data = Z;
		19'b0011101000101001110: color_data = Z;
		19'b0011101000101001111: color_data = Z;
		19'b0011101000101010000: color_data = Z;
		19'b0011101000101010001: color_data = Z;
		19'b0011101000101010010: color_data = Z;
		19'b0011101000101010011: color_data = Z;
		19'b0011101000101010100: color_data = Z;
		19'b0011101000101010101: color_data = Z;
		19'b0011101000101010110: color_data = Z;
		19'b0011101000101010111: color_data = Z;
		19'b0011101000101011000: color_data = Z;
		19'b0011101000101011001: color_data = Z;
		19'b0011101000101011010: color_data = Z;
		19'b0011101000101011011: color_data = Z;
		19'b0011101000101011100: color_data = Z;
		19'b0011101000101011101: color_data = Z;
		19'b0011101000101011110: color_data = Z;
		19'b0011101000101011111: color_data = Z;
		19'b0011101000101100000: color_data = Z;
		19'b0011101000101100001: color_data = Z;
		19'b0011101000101100010: color_data = Z;
		19'b0011101000101100011: color_data = Z;
		19'b0011101000101100100: color_data = Z;
		19'b0011101000101100101: color_data = Z;
		19'b0011101000101100110: color_data = Z;
		19'b0011101000101100111: color_data = Z;
		19'b0011101000101101000: color_data = Z;
		19'b0011101000101101001: color_data = Z;
		19'b0011101000101101010: color_data = Z;
		19'b0011101000101101011: color_data = Z;
		19'b0011101000101101100: color_data = Z;
		19'b0011101000101101101: color_data = Z;
		19'b0011101000101101110: color_data = Z;
		19'b0011101000101101111: color_data = Z;
		19'b0011101000101110000: color_data = Z;
		19'b0011101000101110001: color_data = Z;
		19'b0011101000101110010: color_data = Z;
		19'b0011101000101110011: color_data = Z;
		19'b0011101000101110100: color_data = Z;
		19'b0011101000101110101: color_data = Z;
		19'b0011101000101110110: color_data = Z;
		19'b0011101000101110111: color_data = Z;
		19'b0011101000101111000: color_data = Z;
		19'b0011101000101111001: color_data = Z;
		19'b0011101000101111010: color_data = Z;
		19'b0011101000101111011: color_data = Z;
		19'b0011101000101111100: color_data = Z;
		19'b0011101000101111101: color_data = Z;
		19'b0011101000101111110: color_data = Z;
		19'b0011101000101111111: color_data = Z;
		19'b0011101000110000000: color_data = Z;
		19'b0011101000110000001: color_data = Z;
		19'b0011101000110000010: color_data = Z;
		19'b0011101000110000011: color_data = Z;
		19'b0011101000110000100: color_data = Z;
		19'b0011101000110000101: color_data = Z;
		19'b0011101000110000110: color_data = Z;
		19'b0011101000110000111: color_data = Z;
		19'b0011101000110001000: color_data = Z;
		19'b0011101000110001001: color_data = Z;
		19'b0011101000110001010: color_data = Z;
		19'b0011101000110001011: color_data = Z;
		19'b0011101000110001100: color_data = Z;
		19'b0011101000110001101: color_data = Z;
		19'b0011101000110001110: color_data = Z;
		19'b0011101000110001111: color_data = Z;
		19'b0011101000110010000: color_data = Z;
		19'b0011101000110111100: color_data = Z;
		19'b0011101000110111101: color_data = Z;
		19'b0011101000110111110: color_data = Z;
		19'b0011101000110111111: color_data = Z;
		19'b0011101000111000000: color_data = Z;
		19'b0011101000111000001: color_data = Z;
		19'b0011101000111000010: color_data = Z;
		19'b0011101000111000011: color_data = Z;
		19'b0011101000111000100: color_data = Z;
		19'b0011101000111000101: color_data = Z;
		19'b0011101000111000110: color_data = Z;
		19'b0011101000111000111: color_data = Z;
		19'b0011101000111011110: color_data = Z;
		19'b0011101010010110011: color_data = Z;
		19'b0011101010010110100: color_data = Z;
		19'b0011101010010110101: color_data = Z;
		19'b0011101010010110110: color_data = Z;
		19'b0011101010010110111: color_data = Z;
		19'b0011101010010111000: color_data = Z;
		19'b0011101010010111001: color_data = Z;
		19'b0011101010010111010: color_data = Z;
		19'b0011101010010111011: color_data = Z;
		19'b0011101010010111100: color_data = Z;
		19'b0011101010010111101: color_data = Z;
		19'b0011101010010111110: color_data = Z;
		19'b0011101010010111111: color_data = Z;
		19'b0011101010011000000: color_data = Z;
		19'b0011101010011000001: color_data = Z;
		19'b0011101010011000010: color_data = Z;
		19'b0011101010011000011: color_data = Z;
		19'b0011101010011000100: color_data = Z;
		19'b0011101010011000101: color_data = Z;
		19'b0011101010011000110: color_data = Z;
		19'b0011101010011000111: color_data = Z;
		19'b0011101010011001000: color_data = Z;
		19'b0011101010011001001: color_data = Z;
		19'b0011101010011001010: color_data = Z;
		19'b0011101010011001011: color_data = Z;
		19'b0011101010011001100: color_data = Z;
		19'b0011101010011001101: color_data = Z;
		19'b0011101010011001110: color_data = Z;
		19'b0011101010011001111: color_data = Z;
		19'b0011101010011010000: color_data = Z;
		19'b0011101010011010001: color_data = Z;
		19'b0011101010011010010: color_data = Z;
		19'b0011101010011010011: color_data = Z;
		19'b0011101010011010100: color_data = Z;
		19'b0011101010011010101: color_data = Z;
		19'b0011101010011010110: color_data = Z;
		19'b0011101010011010111: color_data = Z;
		19'b0011101010011011000: color_data = Z;
		19'b0011101010011011001: color_data = Z;
		19'b0011101010011011010: color_data = Z;
		19'b0011101010011011011: color_data = Z;
		19'b0011101010011011100: color_data = Z;
		19'b0011101010011011101: color_data = Z;
		19'b0011101010011011110: color_data = Z;
		19'b0011101010011011111: color_data = Z;
		19'b0011101010011100000: color_data = Z;
		19'b0011101010011100001: color_data = Z;
		19'b0011101010011100010: color_data = Z;
		19'b0011101010011100011: color_data = Z;
		19'b0011101010011100100: color_data = Z;
		19'b0011101010011100101: color_data = Z;
		19'b0011101010011100110: color_data = Z;
		19'b0011101010011100111: color_data = Z;
		19'b0011101010011101000: color_data = Z;
		19'b0011101010011101001: color_data = Z;
		19'b0011101010011101010: color_data = Z;
		19'b0011101010011101011: color_data = Z;
		19'b0011101010011101100: color_data = Z;
		19'b0011101010011101101: color_data = Z;
		19'b0011101010011101110: color_data = Z;
		19'b0011101010011101111: color_data = Z;
		19'b0011101010011110000: color_data = Z;
		19'b0011101010011110001: color_data = Z;
		19'b0011101010011110010: color_data = Z;
		19'b0011101010011110011: color_data = Z;
		19'b0011101010011110100: color_data = Z;
		19'b0011101010011110101: color_data = Z;
		19'b0011101010011110110: color_data = Z;
		19'b0011101010011110111: color_data = Z;
		19'b0011101010011111000: color_data = Z;
		19'b0011101010011111001: color_data = Z;
		19'b0011101010011111010: color_data = Z;
		19'b0011101010011111011: color_data = Z;
		19'b0011101010011111100: color_data = Z;
		19'b0011101010011111101: color_data = Z;
		19'b0011101010011111110: color_data = Z;
		19'b0011101010011111111: color_data = Z;
		19'b0011101010100000000: color_data = Z;
		19'b0011101010100000001: color_data = Z;
		19'b0011101010100000010: color_data = Z;
		19'b0011101010100000011: color_data = Z;
		19'b0011101010100000100: color_data = Z;
		19'b0011101010100000101: color_data = Z;
		19'b0011101010100000110: color_data = Z;
		19'b0011101010100000111: color_data = Z;
		19'b0011101010100001000: color_data = Z;
		19'b0011101010100001001: color_data = Z;
		19'b0011101010100001010: color_data = Z;
		19'b0011101010100001011: color_data = Z;
		19'b0011101010100001100: color_data = Z;
		19'b0011101010100001101: color_data = Z;
		19'b0011101010100001110: color_data = Z;
		19'b0011101010100001111: color_data = Z;
		19'b0011101010100010000: color_data = Z;
		19'b0011101010100010001: color_data = Z;
		19'b0011101010100010010: color_data = Z;
		19'b0011101010100010011: color_data = Z;
		19'b0011101010100010100: color_data = Z;
		19'b0011101010100010101: color_data = Z;
		19'b0011101010100010110: color_data = Z;
		19'b0011101010100010111: color_data = Z;
		19'b0011101010100011000: color_data = Z;
		19'b0011101010100011001: color_data = Z;
		19'b0011101010100011010: color_data = Z;
		19'b0011101010100011011: color_data = Z;
		19'b0011101010100011100: color_data = Z;
		19'b0011101010100011101: color_data = Z;
		19'b0011101010100011110: color_data = Z;
		19'b0011101010100011111: color_data = Z;
		19'b0011101010100100000: color_data = Z;
		19'b0011101010100100001: color_data = Z;
		19'b0011101010100100010: color_data = Z;
		19'b0011101010100100011: color_data = Z;
		19'b0011101010100100100: color_data = Z;
		19'b0011101010100100101: color_data = Z;
		19'b0011101010100100110: color_data = Z;
		19'b0011101010100100111: color_data = Z;
		19'b0011101010100101000: color_data = Z;
		19'b0011101010100101001: color_data = Z;
		19'b0011101010100101010: color_data = Z;
		19'b0011101010100101011: color_data = Z;
		19'b0011101010100101100: color_data = Z;
		19'b0011101010100101101: color_data = Z;
		19'b0011101010100101110: color_data = Z;
		19'b0011101010100101111: color_data = Z;
		19'b0011101010100110000: color_data = Z;
		19'b0011101010100110001: color_data = Z;
		19'b0011101010100110010: color_data = Z;
		19'b0011101010100110011: color_data = Z;
		19'b0011101010100110100: color_data = Z;
		19'b0011101010100110101: color_data = Z;
		19'b0011101010100110110: color_data = Z;
		19'b0011101010100110111: color_data = Z;
		19'b0011101010100111000: color_data = Z;
		19'b0011101010100111001: color_data = Z;
		19'b0011101010100111010: color_data = Z;
		19'b0011101010100111011: color_data = Z;
		19'b0011101010100111100: color_data = Z;
		19'b0011101010100111101: color_data = Z;
		19'b0011101010100111110: color_data = Z;
		19'b0011101010100111111: color_data = Z;
		19'b0011101010101000000: color_data = Z;
		19'b0011101010101000001: color_data = Z;
		19'b0011101010101000010: color_data = Z;
		19'b0011101010101000011: color_data = Z;
		19'b0011101010101000100: color_data = Z;
		19'b0011101010101000101: color_data = Z;
		19'b0011101010101000110: color_data = Z;
		19'b0011101010101000111: color_data = Z;
		19'b0011101010101001000: color_data = Z;
		19'b0011101010101001001: color_data = Z;
		19'b0011101010101001010: color_data = Z;
		19'b0011101010101001011: color_data = Z;
		19'b0011101010101001100: color_data = Z;
		19'b0011101010101001101: color_data = Z;
		19'b0011101010101001110: color_data = Z;
		19'b0011101010101001111: color_data = Z;
		19'b0011101010101010000: color_data = Z;
		19'b0011101010101010001: color_data = Z;
		19'b0011101010101010010: color_data = Z;
		19'b0011101010101010011: color_data = Z;
		19'b0011101010101010100: color_data = Z;
		19'b0011101010101010101: color_data = Z;
		19'b0011101010101010110: color_data = Z;
		19'b0011101010101010111: color_data = Z;
		19'b0011101010101011000: color_data = Z;
		19'b0011101010101011001: color_data = Z;
		19'b0011101010101011010: color_data = Z;
		19'b0011101010101011011: color_data = Z;
		19'b0011101010101011100: color_data = Z;
		19'b0011101010101011101: color_data = Z;
		19'b0011101010101011110: color_data = Z;
		19'b0011101010101011111: color_data = Z;
		19'b0011101010101100000: color_data = Z;
		19'b0011101010101100001: color_data = Z;
		19'b0011101010101100010: color_data = Z;
		19'b0011101010101100011: color_data = Z;
		19'b0011101010101100100: color_data = Z;
		19'b0011101010101100101: color_data = Z;
		19'b0011101010101100110: color_data = Z;
		19'b0011101010101100111: color_data = Z;
		19'b0011101010101101000: color_data = Z;
		19'b0011101010101101001: color_data = Z;
		19'b0011101010101101010: color_data = Z;
		19'b0011101010101101011: color_data = Z;
		19'b0011101010101101100: color_data = Z;
		19'b0011101010101101101: color_data = Z;
		19'b0011101010101101110: color_data = Z;
		19'b0011101010101101111: color_data = Z;
		19'b0011101010101110000: color_data = Z;
		19'b0011101010101110001: color_data = Z;
		19'b0011101010101110010: color_data = Z;
		19'b0011101010101110011: color_data = Z;
		19'b0011101010101110100: color_data = Z;
		19'b0011101010101110101: color_data = Z;
		19'b0011101010101110110: color_data = Z;
		19'b0011101010101110111: color_data = Z;
		19'b0011101010101111000: color_data = Z;
		19'b0011101010101111001: color_data = Z;
		19'b0011101010101111010: color_data = Z;
		19'b0011101010101111011: color_data = Z;
		19'b0011101010101111100: color_data = Z;
		19'b0011101010101111101: color_data = Z;
		19'b0011101010101111110: color_data = Z;
		19'b0011101010101111111: color_data = Z;
		19'b0011101010110000000: color_data = Z;
		19'b0011101010110000001: color_data = Z;
		19'b0011101010110000010: color_data = Z;
		19'b0011101010110000011: color_data = Z;
		19'b0011101010110000100: color_data = Z;
		19'b0011101010110000101: color_data = Z;
		19'b0011101010110000110: color_data = Z;
		19'b0011101010110000111: color_data = Z;
		19'b0011101010110001000: color_data = Z;
		19'b0011101010110001001: color_data = Z;
		19'b0011101010110001010: color_data = Z;
		19'b0011101010110001011: color_data = Z;
		19'b0011101010110001100: color_data = Z;
		19'b0011101010110001101: color_data = Z;
		19'b0011101010110001110: color_data = Z;
		19'b0011101010110001111: color_data = Z;
		19'b0011101010110010000: color_data = Z;
		19'b0011101010110111101: color_data = Z;
		19'b0011101010110111110: color_data = Z;
		19'b0011101010110111111: color_data = Z;
		19'b0011101010111000000: color_data = Z;
		19'b0011101010111000001: color_data = Z;
		19'b0011101010111000010: color_data = Z;
		19'b0011101010111000011: color_data = Z;
		19'b0011101010111000100: color_data = Z;
		19'b0011101010111000101: color_data = Z;
		19'b0011101010111000110: color_data = Z;
		19'b0011101010111000111: color_data = Z;
		19'b0011101100010110101: color_data = Z;
		19'b0011101100010110110: color_data = Z;
		19'b0011101100010110111: color_data = Z;
		19'b0011101100010111000: color_data = Z;
		19'b0011101100010111001: color_data = Z;
		19'b0011101100010111010: color_data = Z;
		19'b0011101100010111011: color_data = Z;
		19'b0011101100010111100: color_data = Z;
		19'b0011101100010111101: color_data = Z;
		19'b0011101100010111110: color_data = Z;
		19'b0011101100010111111: color_data = Z;
		19'b0011101100011000000: color_data = Z;
		19'b0011101100011000001: color_data = Z;
		19'b0011101100011000010: color_data = Z;
		19'b0011101100011000011: color_data = Z;
		19'b0011101100011000100: color_data = Z;
		19'b0011101100011000101: color_data = Z;
		19'b0011101100011000110: color_data = Z;
		19'b0011101100011000111: color_data = Z;
		19'b0011101100011001000: color_data = Z;
		19'b0011101100011001001: color_data = Z;
		19'b0011101100011001010: color_data = Z;
		19'b0011101100011001011: color_data = Z;
		19'b0011101100011001100: color_data = Z;
		19'b0011101100011001101: color_data = Z;
		19'b0011101100011001110: color_data = Z;
		19'b0011101100011001111: color_data = Z;
		19'b0011101100011010000: color_data = Z;
		19'b0011101100011010001: color_data = Z;
		19'b0011101100011010010: color_data = Z;
		19'b0011101100011010011: color_data = Z;
		19'b0011101100011010100: color_data = Z;
		19'b0011101100011010101: color_data = Z;
		19'b0011101100011010110: color_data = Z;
		19'b0011101100011010111: color_data = Z;
		19'b0011101100011011000: color_data = Z;
		19'b0011101100011011001: color_data = Z;
		19'b0011101100011011010: color_data = Z;
		19'b0011101100011011011: color_data = Z;
		19'b0011101100011011100: color_data = Z;
		19'b0011101100011011101: color_data = Z;
		19'b0011101100011011110: color_data = Z;
		19'b0011101100011011111: color_data = Z;
		19'b0011101100011100000: color_data = Z;
		19'b0011101100011100001: color_data = Z;
		19'b0011101100011100010: color_data = Z;
		19'b0011101100011100011: color_data = Z;
		19'b0011101100011100100: color_data = Z;
		19'b0011101100011100101: color_data = Z;
		19'b0011101100011100110: color_data = Z;
		19'b0011101100011100111: color_data = Z;
		19'b0011101100011101000: color_data = Z;
		19'b0011101100011101001: color_data = Z;
		19'b0011101100011101010: color_data = Z;
		19'b0011101100011101011: color_data = Z;
		19'b0011101100011101100: color_data = Z;
		19'b0011101100011101101: color_data = Z;
		19'b0011101100011101110: color_data = Z;
		19'b0011101100011101111: color_data = Z;
		19'b0011101100011110000: color_data = Z;
		19'b0011101100011110001: color_data = Z;
		19'b0011101100011110010: color_data = Z;
		19'b0011101100011110011: color_data = Z;
		19'b0011101100011110100: color_data = Z;
		19'b0011101100011110101: color_data = Z;
		19'b0011101100011110110: color_data = Z;
		19'b0011101100011110111: color_data = Z;
		19'b0011101100011111000: color_data = Z;
		19'b0011101100011111001: color_data = Z;
		19'b0011101100011111010: color_data = Z;
		19'b0011101100011111011: color_data = Z;
		19'b0011101100011111100: color_data = Z;
		19'b0011101100011111101: color_data = Z;
		19'b0011101100011111110: color_data = Z;
		19'b0011101100011111111: color_data = Z;
		19'b0011101100100000000: color_data = Z;
		19'b0011101100100000001: color_data = Z;
		19'b0011101100100000010: color_data = Z;
		19'b0011101100100000011: color_data = Z;
		19'b0011101100100000100: color_data = Z;
		19'b0011101100100000101: color_data = Z;
		19'b0011101100100000110: color_data = Z;
		19'b0011101100100000111: color_data = Z;
		19'b0011101100100001000: color_data = Z;
		19'b0011101100100001001: color_data = Z;
		19'b0011101100100001010: color_data = Z;
		19'b0011101100100001011: color_data = Z;
		19'b0011101100100001100: color_data = Z;
		19'b0011101100100001101: color_data = Z;
		19'b0011101100100001110: color_data = Z;
		19'b0011101100100001111: color_data = Z;
		19'b0011101100100010000: color_data = Z;
		19'b0011101100100010001: color_data = Z;
		19'b0011101100100010010: color_data = Z;
		19'b0011101100100010011: color_data = Z;
		19'b0011101100100010100: color_data = Z;
		19'b0011101100100010101: color_data = Z;
		19'b0011101100100010110: color_data = Z;
		19'b0011101100100010111: color_data = Z;
		19'b0011101100100011000: color_data = Z;
		19'b0011101100100011001: color_data = Z;
		19'b0011101100100011010: color_data = Z;
		19'b0011101100100011011: color_data = Z;
		19'b0011101100100011100: color_data = Z;
		19'b0011101100100011101: color_data = Z;
		19'b0011101100100011110: color_data = Z;
		19'b0011101100100011111: color_data = Z;
		19'b0011101100100100000: color_data = Z;
		19'b0011101100100100001: color_data = Z;
		19'b0011101100100100010: color_data = Z;
		19'b0011101100100100011: color_data = Z;
		19'b0011101100100100100: color_data = Z;
		19'b0011101100100100101: color_data = Z;
		19'b0011101100100100110: color_data = Z;
		19'b0011101100100100111: color_data = Z;
		19'b0011101100100101000: color_data = Z;
		19'b0011101100100101001: color_data = Z;
		19'b0011101100100101010: color_data = Z;
		19'b0011101100100101011: color_data = Z;
		19'b0011101100100101100: color_data = Z;
		19'b0011101100100101101: color_data = Z;
		19'b0011101100100101110: color_data = Z;
		19'b0011101100100101111: color_data = Z;
		19'b0011101100100110000: color_data = Z;
		19'b0011101100100110001: color_data = Z;
		19'b0011101100100110010: color_data = Z;
		19'b0011101100100110011: color_data = Z;
		19'b0011101100100110100: color_data = Z;
		19'b0011101100100110101: color_data = Z;
		19'b0011101100100110110: color_data = Z;
		19'b0011101100100110111: color_data = Z;
		19'b0011101100100111000: color_data = Z;
		19'b0011101100100111001: color_data = Z;
		19'b0011101100100111010: color_data = Z;
		19'b0011101100100111011: color_data = Z;
		19'b0011101100100111100: color_data = Z;
		19'b0011101100100111101: color_data = Z;
		19'b0011101100100111110: color_data = Z;
		19'b0011101100100111111: color_data = Z;
		19'b0011101100101000000: color_data = Z;
		19'b0011101100101000001: color_data = Z;
		19'b0011101100101000010: color_data = Z;
		19'b0011101100101000011: color_data = Z;
		19'b0011101100101000100: color_data = Z;
		19'b0011101100101000101: color_data = Z;
		19'b0011101100101000110: color_data = Z;
		19'b0011101100101000111: color_data = Z;
		19'b0011101100101001000: color_data = Z;
		19'b0011101100101001001: color_data = Z;
		19'b0011101100101001010: color_data = Z;
		19'b0011101100101001011: color_data = Z;
		19'b0011101100101001100: color_data = Z;
		19'b0011101100101001101: color_data = Z;
		19'b0011101100101001110: color_data = Z;
		19'b0011101100101001111: color_data = Z;
		19'b0011101100101010000: color_data = Z;
		19'b0011101100101010001: color_data = Z;
		19'b0011101100101010010: color_data = Z;
		19'b0011101100101010011: color_data = Z;
		19'b0011101100101010100: color_data = Z;
		19'b0011101100101010101: color_data = Z;
		19'b0011101100101010110: color_data = Z;
		19'b0011101100101010111: color_data = Z;
		19'b0011101100101011000: color_data = Z;
		19'b0011101100101011001: color_data = Z;
		19'b0011101100101011010: color_data = Z;
		19'b0011101100101011011: color_data = Z;
		19'b0011101100101011100: color_data = Z;
		19'b0011101100101011101: color_data = Z;
		19'b0011101100101011110: color_data = Z;
		19'b0011101100101011111: color_data = Z;
		19'b0011101100101100000: color_data = Z;
		19'b0011101100101100001: color_data = Z;
		19'b0011101100101100010: color_data = Z;
		19'b0011101100101100011: color_data = Z;
		19'b0011101100101100100: color_data = Z;
		19'b0011101100101100101: color_data = Z;
		19'b0011101100101100110: color_data = Z;
		19'b0011101100101100111: color_data = Z;
		19'b0011101100101101000: color_data = Z;
		19'b0011101100101101001: color_data = Z;
		19'b0011101100101101010: color_data = Z;
		19'b0011101100101101011: color_data = Z;
		19'b0011101100101101100: color_data = Z;
		19'b0011101100101101101: color_data = Z;
		19'b0011101100101101110: color_data = Z;
		19'b0011101100101101111: color_data = Z;
		19'b0011101100101110000: color_data = Z;
		19'b0011101100101110001: color_data = Z;
		19'b0011101100101110010: color_data = Z;
		19'b0011101100101110011: color_data = Z;
		19'b0011101100101110100: color_data = Z;
		19'b0011101100101110101: color_data = Z;
		19'b0011101100101110110: color_data = Z;
		19'b0011101100101110111: color_data = Z;
		19'b0011101100101111000: color_data = Z;
		19'b0011101100101111001: color_data = Z;
		19'b0011101100101111010: color_data = Z;
		19'b0011101100101111011: color_data = Z;
		19'b0011101100101111100: color_data = Z;
		19'b0011101100101111101: color_data = Z;
		19'b0011101100101111110: color_data = Z;
		19'b0011101100101111111: color_data = Z;
		19'b0011101100110000000: color_data = Z;
		19'b0011101100110000001: color_data = Z;
		19'b0011101100110000010: color_data = Z;
		19'b0011101100110000011: color_data = Z;
		19'b0011101100110000100: color_data = Z;
		19'b0011101100110000101: color_data = Z;
		19'b0011101100110000110: color_data = Z;
		19'b0011101100110000111: color_data = Z;
		19'b0011101100110001000: color_data = Z;
		19'b0011101100110001001: color_data = Z;
		19'b0011101100110001010: color_data = Z;
		19'b0011101100110001011: color_data = Z;
		19'b0011101100110001100: color_data = Z;
		19'b0011101100110001101: color_data = Z;
		19'b0011101100110001110: color_data = Z;
		19'b0011101100110001111: color_data = Z;
		19'b0011101100110111111: color_data = Z;
		19'b0011101100111000000: color_data = Z;
		19'b0011101100111000001: color_data = Z;
		19'b0011101100111000010: color_data = Z;
		19'b0011101100111000011: color_data = Z;
		19'b0011101100111000100: color_data = Z;
		19'b0011101100111000101: color_data = Z;
		19'b0011101100111000110: color_data = Z;
		19'b0011101100111000111: color_data = Z;
		19'b0011101100111011100: color_data = Z;
		19'b0011101100111011110: color_data = Z;
		19'b0011101110010110101: color_data = Z;
		19'b0011101110010110110: color_data = Z;
		19'b0011101110010110111: color_data = Z;
		19'b0011101110010111000: color_data = Z;
		19'b0011101110010111001: color_data = Z;
		19'b0011101110010111010: color_data = Z;
		19'b0011101110010111011: color_data = Z;
		19'b0011101110010111100: color_data = Z;
		19'b0011101110010111101: color_data = Z;
		19'b0011101110010111110: color_data = Z;
		19'b0011101110010111111: color_data = Z;
		19'b0011101110011000000: color_data = Z;
		19'b0011101110011000001: color_data = Z;
		19'b0011101110011000010: color_data = Z;
		19'b0011101110011000011: color_data = Z;
		19'b0011101110011000100: color_data = Z;
		19'b0011101110011000101: color_data = Z;
		19'b0011101110011000110: color_data = Z;
		19'b0011101110011000111: color_data = Z;
		19'b0011101110011001000: color_data = Z;
		19'b0011101110011001001: color_data = Z;
		19'b0011101110011001010: color_data = Z;
		19'b0011101110011001011: color_data = Z;
		19'b0011101110011001100: color_data = Z;
		19'b0011101110011001101: color_data = Z;
		19'b0011101110011001110: color_data = Z;
		19'b0011101110011001111: color_data = Z;
		19'b0011101110011010000: color_data = Z;
		19'b0011101110011010001: color_data = Z;
		19'b0011101110011010010: color_data = Z;
		19'b0011101110011010011: color_data = Z;
		19'b0011101110011010100: color_data = Z;
		19'b0011101110011010101: color_data = Z;
		19'b0011101110011010110: color_data = Z;
		19'b0011101110011010111: color_data = Z;
		19'b0011101110011011000: color_data = Z;
		19'b0011101110011011001: color_data = Z;
		19'b0011101110011011010: color_data = Z;
		19'b0011101110011011011: color_data = Z;
		19'b0011101110011011100: color_data = Z;
		19'b0011101110011011101: color_data = Z;
		19'b0011101110011011110: color_data = Z;
		19'b0011101110011011111: color_data = Z;
		19'b0011101110011100000: color_data = Z;
		19'b0011101110011100001: color_data = Z;
		19'b0011101110011100010: color_data = Z;
		19'b0011101110011100011: color_data = Z;
		19'b0011101110011100100: color_data = Z;
		19'b0011101110011100101: color_data = Z;
		19'b0011101110011100110: color_data = Z;
		19'b0011101110011100111: color_data = Z;
		19'b0011101110011101000: color_data = Z;
		19'b0011101110011101001: color_data = Z;
		19'b0011101110011101010: color_data = Z;
		19'b0011101110011101011: color_data = Z;
		19'b0011101110011101100: color_data = Z;
		19'b0011101110011101101: color_data = Z;
		19'b0011101110011101110: color_data = Z;
		19'b0011101110011101111: color_data = Z;
		19'b0011101110011110000: color_data = Z;
		19'b0011101110011110001: color_data = Z;
		19'b0011101110011110010: color_data = Z;
		19'b0011101110011110011: color_data = Z;
		19'b0011101110011110100: color_data = Z;
		19'b0011101110011110101: color_data = Z;
		19'b0011101110011110110: color_data = Z;
		19'b0011101110011110111: color_data = Z;
		19'b0011101110011111000: color_data = Z;
		19'b0011101110011111001: color_data = Z;
		19'b0011101110011111010: color_data = Z;
		19'b0011101110011111011: color_data = Z;
		19'b0011101110011111100: color_data = Z;
		19'b0011101110011111101: color_data = Z;
		19'b0011101110011111110: color_data = Z;
		19'b0011101110011111111: color_data = Z;
		19'b0011101110100000000: color_data = Z;
		19'b0011101110100000001: color_data = Z;
		19'b0011101110100000010: color_data = Z;
		19'b0011101110100000011: color_data = Z;
		19'b0011101110100000100: color_data = Z;
		19'b0011101110100000101: color_data = Z;
		19'b0011101110100000110: color_data = Z;
		19'b0011101110100000111: color_data = Z;
		19'b0011101110100001000: color_data = Z;
		19'b0011101110100001001: color_data = Z;
		19'b0011101110100001010: color_data = Z;
		19'b0011101110100001011: color_data = Z;
		19'b0011101110100001100: color_data = Z;
		19'b0011101110100001101: color_data = Z;
		19'b0011101110100001110: color_data = Z;
		19'b0011101110100001111: color_data = Z;
		19'b0011101110100010000: color_data = Z;
		19'b0011101110100010001: color_data = Z;
		19'b0011101110100010010: color_data = Z;
		19'b0011101110100010011: color_data = Z;
		19'b0011101110100010100: color_data = Z;
		19'b0011101110100010101: color_data = Z;
		19'b0011101110100010110: color_data = Z;
		19'b0011101110100010111: color_data = Z;
		19'b0011101110100011000: color_data = Z;
		19'b0011101110100011001: color_data = Z;
		19'b0011101110100011010: color_data = Z;
		19'b0011101110100011011: color_data = Z;
		19'b0011101110100011100: color_data = Z;
		19'b0011101110100011101: color_data = Z;
		19'b0011101110100011110: color_data = Z;
		19'b0011101110100011111: color_data = Z;
		19'b0011101110100100000: color_data = Z;
		19'b0011101110100100001: color_data = Z;
		19'b0011101110100100010: color_data = Z;
		19'b0011101110100100011: color_data = Z;
		19'b0011101110100100100: color_data = Z;
		19'b0011101110100100101: color_data = Z;
		19'b0011101110100100110: color_data = Z;
		19'b0011101110100100111: color_data = Z;
		19'b0011101110100101000: color_data = Z;
		19'b0011101110100101001: color_data = Z;
		19'b0011101110100101010: color_data = Z;
		19'b0011101110100101011: color_data = Z;
		19'b0011101110100101100: color_data = Z;
		19'b0011101110100101101: color_data = Z;
		19'b0011101110100101110: color_data = Z;
		19'b0011101110100101111: color_data = Z;
		19'b0011101110100110000: color_data = Z;
		19'b0011101110100110001: color_data = Z;
		19'b0011101110100110010: color_data = Z;
		19'b0011101110100110011: color_data = Z;
		19'b0011101110100110100: color_data = Z;
		19'b0011101110100110101: color_data = Z;
		19'b0011101110100110110: color_data = Z;
		19'b0011101110100110111: color_data = Z;
		19'b0011101110100111000: color_data = Z;
		19'b0011101110100111001: color_data = Z;
		19'b0011101110100111010: color_data = Z;
		19'b0011101110100111011: color_data = Z;
		19'b0011101110100111100: color_data = Z;
		19'b0011101110100111101: color_data = Z;
		19'b0011101110100111110: color_data = Z;
		19'b0011101110100111111: color_data = Z;
		19'b0011101110101000000: color_data = Z;
		19'b0011101110101000001: color_data = Z;
		19'b0011101110101000010: color_data = Z;
		19'b0011101110101000011: color_data = Z;
		19'b0011101110101000100: color_data = Z;
		19'b0011101110101000101: color_data = Z;
		19'b0011101110101000110: color_data = Z;
		19'b0011101110101000111: color_data = Z;
		19'b0011101110101001000: color_data = Z;
		19'b0011101110101001001: color_data = Z;
		19'b0011101110101001010: color_data = Z;
		19'b0011101110101001011: color_data = Z;
		19'b0011101110101001100: color_data = Z;
		19'b0011101110101001101: color_data = Z;
		19'b0011101110101001110: color_data = Z;
		19'b0011101110101001111: color_data = Z;
		19'b0011101110101010000: color_data = Z;
		19'b0011101110101010001: color_data = Z;
		19'b0011101110101010010: color_data = Z;
		19'b0011101110101010011: color_data = Z;
		19'b0011101110101010100: color_data = Z;
		19'b0011101110101010101: color_data = Z;
		19'b0011101110101010110: color_data = Z;
		19'b0011101110101010111: color_data = Z;
		19'b0011101110101011000: color_data = Z;
		19'b0011101110101011001: color_data = Z;
		19'b0011101110101011010: color_data = Z;
		19'b0011101110101011011: color_data = Z;
		19'b0011101110101011100: color_data = Z;
		19'b0011101110101011101: color_data = Z;
		19'b0011101110101011110: color_data = Z;
		19'b0011101110101011111: color_data = Z;
		19'b0011101110101100000: color_data = Z;
		19'b0011101110101100001: color_data = Z;
		19'b0011101110101100010: color_data = Z;
		19'b0011101110101100011: color_data = Z;
		19'b0011101110101100100: color_data = Z;
		19'b0011101110101100101: color_data = Z;
		19'b0011101110101100110: color_data = Z;
		19'b0011101110101100111: color_data = Z;
		19'b0011101110101101000: color_data = Z;
		19'b0011101110101101001: color_data = Z;
		19'b0011101110101101010: color_data = Z;
		19'b0011101110101101011: color_data = Z;
		19'b0011101110101101100: color_data = Z;
		19'b0011101110101101101: color_data = Z;
		19'b0011101110101101110: color_data = Z;
		19'b0011101110101101111: color_data = Z;
		19'b0011101110101110000: color_data = Z;
		19'b0011101110101110001: color_data = Z;
		19'b0011101110101110010: color_data = Z;
		19'b0011101110101110011: color_data = Z;
		19'b0011101110101110100: color_data = Z;
		19'b0011101110101110101: color_data = Z;
		19'b0011101110101110110: color_data = Z;
		19'b0011101110101110111: color_data = Z;
		19'b0011101110101111000: color_data = Z;
		19'b0011101110101111001: color_data = Z;
		19'b0011101110101111010: color_data = Z;
		19'b0011101110101111011: color_data = Z;
		19'b0011101110101111100: color_data = Z;
		19'b0011101110101111101: color_data = Z;
		19'b0011101110101111110: color_data = Z;
		19'b0011101110101111111: color_data = Z;
		19'b0011101110110000000: color_data = Z;
		19'b0011101110110000001: color_data = Z;
		19'b0011101110110000010: color_data = Z;
		19'b0011101110110000011: color_data = Z;
		19'b0011101110110000100: color_data = Z;
		19'b0011101110110000101: color_data = Z;
		19'b0011101110110000110: color_data = Z;
		19'b0011101110110000111: color_data = Z;
		19'b0011101110110001000: color_data = Z;
		19'b0011101110110001001: color_data = Z;
		19'b0011101110110001010: color_data = Z;
		19'b0011101110110001011: color_data = Z;
		19'b0011101110110001100: color_data = Z;
		19'b0011101110110001101: color_data = Z;
		19'b0011101110110001110: color_data = Z;
		19'b0011101110111000010: color_data = Z;
		19'b0011101110111000011: color_data = Z;
		19'b0011101110111000100: color_data = Z;
		19'b0011101110111000101: color_data = Z;
		19'b0011101110111000110: color_data = Z;
		19'b0011101110111000111: color_data = Z;
		19'b0011101110111001000: color_data = Z;
		19'b0011101110111001001: color_data = Z;
		19'b0011101110111001010: color_data = Z;
		19'b0011101110111001011: color_data = Z;
		19'b0011101110111011010: color_data = Z;
		19'b0011101110111011011: color_data = Z;
		19'b0011101110111011100: color_data = Z;
		19'b0011101110111011101: color_data = Z;
		19'b0011101110111011110: color_data = Z;
		19'b0011101110111011111: color_data = Z;
		19'b0011110000010110100: color_data = Z;
		19'b0011110000010110101: color_data = Z;
		19'b0011110000010110110: color_data = Z;
		19'b0011110000010110111: color_data = Z;
		19'b0011110000010111000: color_data = Z;
		19'b0011110000010111001: color_data = Z;
		19'b0011110000010111010: color_data = Z;
		19'b0011110000010111011: color_data = Z;
		19'b0011110000010111100: color_data = Z;
		19'b0011110000010111101: color_data = Z;
		19'b0011110000010111110: color_data = Z;
		19'b0011110000010111111: color_data = Z;
		19'b0011110000011000000: color_data = Z;
		19'b0011110000011000001: color_data = Z;
		19'b0011110000011000010: color_data = Z;
		19'b0011110000011000011: color_data = Z;
		19'b0011110000011000100: color_data = Z;
		19'b0011110000011000101: color_data = Z;
		19'b0011110000011000110: color_data = Z;
		19'b0011110000011000111: color_data = Z;
		19'b0011110000011001000: color_data = Z;
		19'b0011110000011001001: color_data = Z;
		19'b0011110000011001010: color_data = Z;
		19'b0011110000011001011: color_data = Z;
		19'b0011110000011010010: color_data = Z;
		19'b0011110000011010011: color_data = Z;
		19'b0011110000011010100: color_data = Z;
		19'b0011110000011010101: color_data = Z;
		19'b0011110000011010110: color_data = Z;
		19'b0011110000011010111: color_data = Z;
		19'b0011110000011011000: color_data = Z;
		19'b0011110000011011001: color_data = Z;
		19'b0011110000011011010: color_data = Z;
		19'b0011110000011011011: color_data = Z;
		19'b0011110000011011100: color_data = Z;
		19'b0011110000011011101: color_data = Z;
		19'b0011110000011011110: color_data = Z;
		19'b0011110000011011111: color_data = Z;
		19'b0011110000011100000: color_data = Z;
		19'b0011110000011100001: color_data = Z;
		19'b0011110000011100010: color_data = Z;
		19'b0011110000011100011: color_data = Z;
		19'b0011110000011100100: color_data = Z;
		19'b0011110000011100101: color_data = Z;
		19'b0011110000011100110: color_data = Z;
		19'b0011110000011100111: color_data = Z;
		19'b0011110000011101000: color_data = Z;
		19'b0011110000011101001: color_data = Z;
		19'b0011110000011101010: color_data = Z;
		19'b0011110000011101011: color_data = Z;
		19'b0011110000011101100: color_data = Z;
		19'b0011110000011101101: color_data = Z;
		19'b0011110000011101110: color_data = Z;
		19'b0011110000011101111: color_data = Z;
		19'b0011110000011110000: color_data = Z;
		19'b0011110000011110001: color_data = Z;
		19'b0011110000011110010: color_data = Z;
		19'b0011110000011110011: color_data = Z;
		19'b0011110000011110100: color_data = Z;
		19'b0011110000011110101: color_data = Z;
		19'b0011110000011110110: color_data = Z;
		19'b0011110000011110111: color_data = Z;
		19'b0011110000011111000: color_data = Z;
		19'b0011110000011111001: color_data = Z;
		19'b0011110000011111010: color_data = Z;
		19'b0011110000011111011: color_data = Z;
		19'b0011110000011111100: color_data = Z;
		19'b0011110000011111101: color_data = Z;
		19'b0011110000011111110: color_data = Z;
		19'b0011110000011111111: color_data = Z;
		19'b0011110000100000000: color_data = Z;
		19'b0011110000100000001: color_data = Z;
		19'b0011110000100000010: color_data = Z;
		19'b0011110000100000011: color_data = Z;
		19'b0011110000100000100: color_data = Z;
		19'b0011110000100000101: color_data = Z;
		19'b0011110000100000110: color_data = Z;
		19'b0011110000100000111: color_data = Z;
		19'b0011110000100001000: color_data = Z;
		19'b0011110000100001001: color_data = Z;
		19'b0011110000100001010: color_data = Z;
		19'b0011110000100001011: color_data = Z;
		19'b0011110000100001100: color_data = Z;
		19'b0011110000100001101: color_data = Z;
		19'b0011110000100001110: color_data = Z;
		19'b0011110000100001111: color_data = Z;
		19'b0011110000100010000: color_data = Z;
		19'b0011110000100010001: color_data = Z;
		19'b0011110000100010010: color_data = Z;
		19'b0011110000100010011: color_data = Z;
		19'b0011110000100010100: color_data = Z;
		19'b0011110000100010101: color_data = Z;
		19'b0011110000100010110: color_data = Z;
		19'b0011110000100010111: color_data = Z;
		19'b0011110000100011000: color_data = Z;
		19'b0011110000100011001: color_data = Z;
		19'b0011110000100011010: color_data = Z;
		19'b0011110000100011011: color_data = Z;
		19'b0011110000100011100: color_data = Z;
		19'b0011110000100011101: color_data = Z;
		19'b0011110000100011110: color_data = Z;
		19'b0011110000100011111: color_data = Z;
		19'b0011110000100100000: color_data = Z;
		19'b0011110000100100001: color_data = Z;
		19'b0011110000100100010: color_data = Z;
		19'b0011110000100100011: color_data = Z;
		19'b0011110000100100100: color_data = Z;
		19'b0011110000100100101: color_data = Z;
		19'b0011110000100100110: color_data = Z;
		19'b0011110000100100111: color_data = Z;
		19'b0011110000100101000: color_data = Z;
		19'b0011110000100101001: color_data = Z;
		19'b0011110000100101010: color_data = Z;
		19'b0011110000100101011: color_data = Z;
		19'b0011110000100101100: color_data = Z;
		19'b0011110000100101101: color_data = Z;
		19'b0011110000100101110: color_data = Z;
		19'b0011110000100101111: color_data = Z;
		19'b0011110000100110000: color_data = Z;
		19'b0011110000100110001: color_data = Z;
		19'b0011110000100110010: color_data = Z;
		19'b0011110000100110011: color_data = Z;
		19'b0011110000100110100: color_data = Z;
		19'b0011110000100110101: color_data = Z;
		19'b0011110000100110110: color_data = Z;
		19'b0011110000100110111: color_data = Z;
		19'b0011110000100111000: color_data = Z;
		19'b0011110000100111001: color_data = Z;
		19'b0011110000100111010: color_data = Z;
		19'b0011110000100111011: color_data = Z;
		19'b0011110000100111100: color_data = Z;
		19'b0011110000100111101: color_data = Z;
		19'b0011110000100111110: color_data = Z;
		19'b0011110000100111111: color_data = Z;
		19'b0011110000101000000: color_data = Z;
		19'b0011110000101000001: color_data = Z;
		19'b0011110000101000010: color_data = Z;
		19'b0011110000101000011: color_data = Z;
		19'b0011110000101000100: color_data = Z;
		19'b0011110000101000101: color_data = Z;
		19'b0011110000101000110: color_data = Z;
		19'b0011110000101000111: color_data = Z;
		19'b0011110000101001000: color_data = Z;
		19'b0011110000101001001: color_data = Z;
		19'b0011110000101001010: color_data = Z;
		19'b0011110000101001011: color_data = Z;
		19'b0011110000101001100: color_data = Z;
		19'b0011110000101001101: color_data = Z;
		19'b0011110000101001110: color_data = Z;
		19'b0011110000101001111: color_data = Z;
		19'b0011110000101010000: color_data = Z;
		19'b0011110000101010001: color_data = Z;
		19'b0011110000101010010: color_data = Z;
		19'b0011110000101010011: color_data = Z;
		19'b0011110000101010100: color_data = Z;
		19'b0011110000101010101: color_data = Z;
		19'b0011110000101010110: color_data = Z;
		19'b0011110000101010111: color_data = Z;
		19'b0011110000101011000: color_data = Z;
		19'b0011110000101011001: color_data = Z;
		19'b0011110000101011010: color_data = Z;
		19'b0011110000101011011: color_data = Z;
		19'b0011110000101011100: color_data = Z;
		19'b0011110000101011101: color_data = Z;
		19'b0011110000101011110: color_data = Z;
		19'b0011110000101011111: color_data = Z;
		19'b0011110000101100000: color_data = Z;
		19'b0011110000101100001: color_data = Z;
		19'b0011110000101100010: color_data = Z;
		19'b0011110000101100011: color_data = Z;
		19'b0011110000101100100: color_data = Z;
		19'b0011110000101100101: color_data = Z;
		19'b0011110000101100110: color_data = Z;
		19'b0011110000101100111: color_data = Z;
		19'b0011110000101101000: color_data = Z;
		19'b0011110000101101001: color_data = Z;
		19'b0011110000101101010: color_data = Z;
		19'b0011110000101101011: color_data = Z;
		19'b0011110000101101100: color_data = Z;
		19'b0011110000101101101: color_data = Z;
		19'b0011110000101101110: color_data = Z;
		19'b0011110000101101111: color_data = Z;
		19'b0011110000101110000: color_data = Z;
		19'b0011110000101110001: color_data = Z;
		19'b0011110000101110010: color_data = Z;
		19'b0011110000101110011: color_data = Z;
		19'b0011110000101110100: color_data = Z;
		19'b0011110000101110101: color_data = Z;
		19'b0011110000101110110: color_data = Z;
		19'b0011110000101110111: color_data = Z;
		19'b0011110000101111000: color_data = Z;
		19'b0011110000101111001: color_data = Z;
		19'b0011110000101111010: color_data = Z;
		19'b0011110000101111011: color_data = Z;
		19'b0011110000101111100: color_data = Z;
		19'b0011110000101111101: color_data = Z;
		19'b0011110000101111110: color_data = Z;
		19'b0011110000101111111: color_data = Z;
		19'b0011110000110000000: color_data = Z;
		19'b0011110000110000001: color_data = Z;
		19'b0011110000110000010: color_data = Z;
		19'b0011110000110000011: color_data = Z;
		19'b0011110000110000100: color_data = Z;
		19'b0011110000110000101: color_data = Z;
		19'b0011110000110000110: color_data = Z;
		19'b0011110000110000111: color_data = Z;
		19'b0011110000110001000: color_data = Z;
		19'b0011110000110001001: color_data = Z;
		19'b0011110000110001010: color_data = Z;
		19'b0011110000110001011: color_data = Z;
		19'b0011110000110001100: color_data = Z;
		19'b0011110000110001101: color_data = Z;
		19'b0011110000111000011: color_data = Z;
		19'b0011110000111000100: color_data = Z;
		19'b0011110000111000101: color_data = Z;
		19'b0011110000111000110: color_data = Z;
		19'b0011110000111000111: color_data = Z;
		19'b0011110000111001000: color_data = Z;
		19'b0011110000111011010: color_data = Z;
		19'b0011110000111011011: color_data = Z;
		19'b0011110000111011100: color_data = Z;
		19'b0011110000111011101: color_data = Z;
		19'b0011110000111011110: color_data = Z;
		19'b0011110000111011111: color_data = Z;
		19'b0011110010010110011: color_data = Z;
		19'b0011110010010110100: color_data = Z;
		19'b0011110010010110101: color_data = Z;
		19'b0011110010010110110: color_data = Z;
		19'b0011110010010111000: color_data = Z;
		19'b0011110010010111001: color_data = Z;
		19'b0011110010010111010: color_data = Z;
		19'b0011110010010111011: color_data = Z;
		19'b0011110010010111100: color_data = Z;
		19'b0011110010010111101: color_data = Z;
		19'b0011110010010111110: color_data = Z;
		19'b0011110010010111111: color_data = Z;
		19'b0011110010011000000: color_data = Z;
		19'b0011110010011000001: color_data = Z;
		19'b0011110010011000010: color_data = Z;
		19'b0011110010011000011: color_data = Z;
		19'b0011110010011000100: color_data = Z;
		19'b0011110010011000101: color_data = Z;
		19'b0011110010011000110: color_data = Z;
		19'b0011110010011000111: color_data = Z;
		19'b0011110010011001000: color_data = Z;
		19'b0011110010011001001: color_data = Z;
		19'b0011110010011001010: color_data = Z;
		19'b0011110010011010010: color_data = Z;
		19'b0011110010011010011: color_data = Z;
		19'b0011110010011010100: color_data = Z;
		19'b0011110010011010101: color_data = Z;
		19'b0011110010011010110: color_data = Z;
		19'b0011110010011010111: color_data = Z;
		19'b0011110010011011000: color_data = Z;
		19'b0011110010011011001: color_data = Z;
		19'b0011110010011011010: color_data = Z;
		19'b0011110010011011011: color_data = Z;
		19'b0011110010011011100: color_data = Z;
		19'b0011110010011011101: color_data = Z;
		19'b0011110010011011110: color_data = Z;
		19'b0011110010011011111: color_data = Z;
		19'b0011110010011100000: color_data = Z;
		19'b0011110010011100001: color_data = Z;
		19'b0011110010011100010: color_data = Z;
		19'b0011110010011100011: color_data = Z;
		19'b0011110010011100100: color_data = Z;
		19'b0011110010011100101: color_data = Z;
		19'b0011110010011100110: color_data = Z;
		19'b0011110010011100111: color_data = Z;
		19'b0011110010011101000: color_data = Z;
		19'b0011110010011101001: color_data = Z;
		19'b0011110010011101010: color_data = Z;
		19'b0011110010011101011: color_data = Z;
		19'b0011110010011101100: color_data = Z;
		19'b0011110010011101101: color_data = Z;
		19'b0011110010011101110: color_data = Z;
		19'b0011110010011101111: color_data = Z;
		19'b0011110010011110000: color_data = Z;
		19'b0011110010011110001: color_data = Z;
		19'b0011110010011110010: color_data = Z;
		19'b0011110010011110011: color_data = Z;
		19'b0011110010011110100: color_data = Z;
		19'b0011110010011110101: color_data = Z;
		19'b0011110010011110110: color_data = Z;
		19'b0011110010011110111: color_data = Z;
		19'b0011110010011111000: color_data = Z;
		19'b0011110010011111001: color_data = Z;
		19'b0011110010011111010: color_data = Z;
		19'b0011110010011111011: color_data = Z;
		19'b0011110010011111100: color_data = Z;
		19'b0011110010011111101: color_data = Z;
		19'b0011110010011111110: color_data = Z;
		19'b0011110010011111111: color_data = Z;
		19'b0011110010100000000: color_data = Z;
		19'b0011110010100000001: color_data = Z;
		19'b0011110010100000010: color_data = Z;
		19'b0011110010100000011: color_data = Z;
		19'b0011110010100000100: color_data = Z;
		19'b0011110010100000101: color_data = Z;
		19'b0011110010100000110: color_data = Z;
		19'b0011110010100000111: color_data = Z;
		19'b0011110010100001000: color_data = Z;
		19'b0011110010100001001: color_data = Z;
		19'b0011110010100001010: color_data = Z;
		19'b0011110010100001011: color_data = Z;
		19'b0011110010100001100: color_data = Z;
		19'b0011110010100001101: color_data = Z;
		19'b0011110010100001110: color_data = Z;
		19'b0011110010100001111: color_data = Z;
		19'b0011110010100010000: color_data = Z;
		19'b0011110010100010001: color_data = Z;
		19'b0011110010100010010: color_data = Z;
		19'b0011110010100010011: color_data = Z;
		19'b0011110010100010100: color_data = Z;
		19'b0011110010100010101: color_data = Z;
		19'b0011110010100010110: color_data = Z;
		19'b0011110010100010111: color_data = Z;
		19'b0011110010100011000: color_data = Z;
		19'b0011110010100011001: color_data = Z;
		19'b0011110010100011010: color_data = Z;
		19'b0011110010100011011: color_data = Z;
		19'b0011110010100011100: color_data = Z;
		19'b0011110010100011101: color_data = Z;
		19'b0011110010100011110: color_data = Z;
		19'b0011110010100011111: color_data = Z;
		19'b0011110010100100000: color_data = Z;
		19'b0011110010100100001: color_data = Z;
		19'b0011110010100100010: color_data = Z;
		19'b0011110010100100011: color_data = Z;
		19'b0011110010100100100: color_data = Z;
		19'b0011110010100100101: color_data = Z;
		19'b0011110010100100110: color_data = Z;
		19'b0011110010100100111: color_data = Z;
		19'b0011110010100101000: color_data = Z;
		19'b0011110010100101001: color_data = Z;
		19'b0011110010100101010: color_data = Z;
		19'b0011110010100101011: color_data = Z;
		19'b0011110010100101100: color_data = Z;
		19'b0011110010100101101: color_data = Z;
		19'b0011110010100101110: color_data = Z;
		19'b0011110010100101111: color_data = Z;
		19'b0011110010100110000: color_data = Z;
		19'b0011110010100110001: color_data = Z;
		19'b0011110010100110010: color_data = Z;
		19'b0011110010100110011: color_data = Z;
		19'b0011110010100110100: color_data = Z;
		19'b0011110010100110101: color_data = Z;
		19'b0011110010100110110: color_data = Z;
		19'b0011110010100110111: color_data = Z;
		19'b0011110010100111000: color_data = Z;
		19'b0011110010100111001: color_data = Z;
		19'b0011110010100111010: color_data = Z;
		19'b0011110010100111011: color_data = Z;
		19'b0011110010100111100: color_data = Z;
		19'b0011110010100111101: color_data = Z;
		19'b0011110010100111110: color_data = Z;
		19'b0011110010100111111: color_data = Z;
		19'b0011110010101000000: color_data = Z;
		19'b0011110010101000001: color_data = Z;
		19'b0011110010101000010: color_data = Z;
		19'b0011110010101000011: color_data = Z;
		19'b0011110010101000100: color_data = Z;
		19'b0011110010101000101: color_data = Z;
		19'b0011110010101000110: color_data = Z;
		19'b0011110010101000111: color_data = Z;
		19'b0011110010101001000: color_data = Z;
		19'b0011110010101001001: color_data = Z;
		19'b0011110010101001010: color_data = Z;
		19'b0011110010101001011: color_data = Z;
		19'b0011110010101001100: color_data = Z;
		19'b0011110010101001101: color_data = Z;
		19'b0011110010101001110: color_data = Z;
		19'b0011110010101001111: color_data = Z;
		19'b0011110010101010000: color_data = Z;
		19'b0011110010101010001: color_data = Z;
		19'b0011110010101010010: color_data = Z;
		19'b0011110010101010011: color_data = Z;
		19'b0011110010101010100: color_data = Z;
		19'b0011110010101010101: color_data = Z;
		19'b0011110010101010110: color_data = Z;
		19'b0011110010101010111: color_data = Z;
		19'b0011110010101011000: color_data = Z;
		19'b0011110010101011001: color_data = Z;
		19'b0011110010101011010: color_data = Z;
		19'b0011110010101011011: color_data = Z;
		19'b0011110010101011100: color_data = Z;
		19'b0011110010101011101: color_data = Z;
		19'b0011110010101011110: color_data = Z;
		19'b0011110010101011111: color_data = Z;
		19'b0011110010101100000: color_data = Z;
		19'b0011110010101100001: color_data = Z;
		19'b0011110010101100010: color_data = Z;
		19'b0011110010101100011: color_data = Z;
		19'b0011110010101100100: color_data = Z;
		19'b0011110010101100101: color_data = Z;
		19'b0011110010101100110: color_data = Z;
		19'b0011110010101100111: color_data = Z;
		19'b0011110010101101000: color_data = Z;
		19'b0011110010101101001: color_data = Z;
		19'b0011110010101101010: color_data = Z;
		19'b0011110010101101011: color_data = Z;
		19'b0011110010101101100: color_data = Z;
		19'b0011110010101101101: color_data = Z;
		19'b0011110010101101110: color_data = Z;
		19'b0011110010101101111: color_data = Z;
		19'b0011110010101110000: color_data = Z;
		19'b0011110010101110001: color_data = Z;
		19'b0011110010101110010: color_data = Z;
		19'b0011110010101110011: color_data = Z;
		19'b0011110010101110100: color_data = Z;
		19'b0011110010101110101: color_data = Z;
		19'b0011110010101110110: color_data = Z;
		19'b0011110010101110111: color_data = Z;
		19'b0011110010101111000: color_data = Z;
		19'b0011110010101111001: color_data = Z;
		19'b0011110010101111010: color_data = Z;
		19'b0011110010101111011: color_data = Z;
		19'b0011110010101111100: color_data = Z;
		19'b0011110010101111101: color_data = Z;
		19'b0011110010101111110: color_data = Z;
		19'b0011110010101111111: color_data = Z;
		19'b0011110010110000000: color_data = Z;
		19'b0011110010110000001: color_data = Z;
		19'b0011110010110000010: color_data = Z;
		19'b0011110010110000011: color_data = Z;
		19'b0011110010110000100: color_data = Z;
		19'b0011110010110000101: color_data = Z;
		19'b0011110010110000110: color_data = Z;
		19'b0011110010110000111: color_data = Z;
		19'b0011110010110001000: color_data = Z;
		19'b0011110010110001001: color_data = Z;
		19'b0011110010110001010: color_data = Z;
		19'b0011110010110001011: color_data = Z;
		19'b0011110010110001100: color_data = Z;
		19'b0011110010110001101: color_data = Z;
		19'b0011110010111000100: color_data = Z;
		19'b0011110010111000101: color_data = Z;
		19'b0011110010111000110: color_data = Z;
		19'b0011110010111011010: color_data = Z;
		19'b0011110010111011011: color_data = Z;
		19'b0011110010111011101: color_data = Z;
		19'b0011110010111011110: color_data = Z;
		19'b0011110010111011111: color_data = Z;
		19'b0011110100010110010: color_data = Z;
		19'b0011110100010110011: color_data = Z;
		19'b0011110100010110100: color_data = Z;
		19'b0011110100010110101: color_data = Z;
		19'b0011110100010110110: color_data = Z;
		19'b0011110100010111000: color_data = Z;
		19'b0011110100010111001: color_data = Z;
		19'b0011110100010111010: color_data = Z;
		19'b0011110100010111011: color_data = Z;
		19'b0011110100010111100: color_data = Z;
		19'b0011110100010111101: color_data = Z;
		19'b0011110100010111110: color_data = Z;
		19'b0011110100010111111: color_data = Z;
		19'b0011110100011000000: color_data = Z;
		19'b0011110100011000001: color_data = Z;
		19'b0011110100011000010: color_data = Z;
		19'b0011110100011000011: color_data = Z;
		19'b0011110100011000100: color_data = Z;
		19'b0011110100011000101: color_data = Z;
		19'b0011110100011000110: color_data = Z;
		19'b0011110100011000111: color_data = Z;
		19'b0011110100011001000: color_data = Z;
		19'b0011110100011010010: color_data = Z;
		19'b0011110100011010011: color_data = Z;
		19'b0011110100011010100: color_data = Z;
		19'b0011110100011010101: color_data = Z;
		19'b0011110100011010110: color_data = Z;
		19'b0011110100011011001: color_data = Z;
		19'b0011110100011011010: color_data = Z;
		19'b0011110100011011011: color_data = Z;
		19'b0011110100011011100: color_data = Z;
		19'b0011110100011011101: color_data = Z;
		19'b0011110100011011110: color_data = Z;
		19'b0011110100011011111: color_data = Z;
		19'b0011110100011100000: color_data = Z;
		19'b0011110100011100001: color_data = Z;
		19'b0011110100011100010: color_data = Z;
		19'b0011110100011100011: color_data = Z;
		19'b0011110100011100100: color_data = Z;
		19'b0011110100011100101: color_data = Z;
		19'b0011110100011100110: color_data = Z;
		19'b0011110100011100111: color_data = Z;
		19'b0011110100011101000: color_data = Z;
		19'b0011110100011101001: color_data = Z;
		19'b0011110100011101010: color_data = Z;
		19'b0011110100011101011: color_data = Z;
		19'b0011110100011101100: color_data = Z;
		19'b0011110100011101101: color_data = Z;
		19'b0011110100011101110: color_data = Z;
		19'b0011110100011101111: color_data = Z;
		19'b0011110100011110000: color_data = Z;
		19'b0011110100011110001: color_data = Z;
		19'b0011110100011110010: color_data = Z;
		19'b0011110100011110011: color_data = Z;
		19'b0011110100011110100: color_data = Z;
		19'b0011110100011110101: color_data = Z;
		19'b0011110100011110110: color_data = Z;
		19'b0011110100011110111: color_data = Z;
		19'b0011110100011111000: color_data = Z;
		19'b0011110100011111001: color_data = Z;
		19'b0011110100011111010: color_data = Z;
		19'b0011110100011111011: color_data = Z;
		19'b0011110100011111100: color_data = Z;
		19'b0011110100011111101: color_data = Z;
		19'b0011110100011111110: color_data = Z;
		19'b0011110100011111111: color_data = Z;
		19'b0011110100100000000: color_data = Z;
		19'b0011110100100000001: color_data = Z;
		19'b0011110100100000010: color_data = Z;
		19'b0011110100100000011: color_data = Z;
		19'b0011110100100000100: color_data = Z;
		19'b0011110100100000101: color_data = Z;
		19'b0011110100100000110: color_data = Z;
		19'b0011110100100000111: color_data = Z;
		19'b0011110100100001000: color_data = Z;
		19'b0011110100100001001: color_data = Z;
		19'b0011110100100001010: color_data = Z;
		19'b0011110100100001011: color_data = Z;
		19'b0011110100100001100: color_data = Z;
		19'b0011110100100001101: color_data = Z;
		19'b0011110100100001110: color_data = Z;
		19'b0011110100100001111: color_data = Z;
		19'b0011110100100010000: color_data = Z;
		19'b0011110100100010001: color_data = Z;
		19'b0011110100100010010: color_data = Z;
		19'b0011110100100010011: color_data = Z;
		19'b0011110100100010100: color_data = Z;
		19'b0011110100100010101: color_data = Z;
		19'b0011110100100010110: color_data = Z;
		19'b0011110100100010111: color_data = Z;
		19'b0011110100100011000: color_data = Z;
		19'b0011110100100011001: color_data = Z;
		19'b0011110100100011010: color_data = Z;
		19'b0011110100100011011: color_data = Z;
		19'b0011110100100011100: color_data = Z;
		19'b0011110100100011101: color_data = Z;
		19'b0011110100100011110: color_data = Z;
		19'b0011110100100011111: color_data = Z;
		19'b0011110100100100000: color_data = Z;
		19'b0011110100100100001: color_data = Z;
		19'b0011110100100100010: color_data = Z;
		19'b0011110100100100011: color_data = Z;
		19'b0011110100100100100: color_data = Z;
		19'b0011110100100100101: color_data = Z;
		19'b0011110100100100110: color_data = Z;
		19'b0011110100100100111: color_data = Z;
		19'b0011110100100101000: color_data = Z;
		19'b0011110100100101001: color_data = Z;
		19'b0011110100100101010: color_data = Z;
		19'b0011110100100101011: color_data = Z;
		19'b0011110100100101100: color_data = Z;
		19'b0011110100100101101: color_data = Z;
		19'b0011110100100101110: color_data = Z;
		19'b0011110100100101111: color_data = Z;
		19'b0011110100100110000: color_data = Z;
		19'b0011110100100110001: color_data = Z;
		19'b0011110100100110010: color_data = Z;
		19'b0011110100100110011: color_data = Z;
		19'b0011110100100110100: color_data = Z;
		19'b0011110100100110101: color_data = Z;
		19'b0011110100100110110: color_data = Z;
		19'b0011110100100110111: color_data = Z;
		19'b0011110100100111000: color_data = Z;
		19'b0011110100100111001: color_data = Z;
		19'b0011110100100111010: color_data = Z;
		19'b0011110100100111011: color_data = Z;
		19'b0011110100100111100: color_data = Z;
		19'b0011110100100111101: color_data = Z;
		19'b0011110100100111110: color_data = Z;
		19'b0011110100100111111: color_data = Z;
		19'b0011110100101000000: color_data = Z;
		19'b0011110100101000001: color_data = Z;
		19'b0011110100101000010: color_data = Z;
		19'b0011110100101000011: color_data = Z;
		19'b0011110100101000100: color_data = Z;
		19'b0011110100101000101: color_data = Z;
		19'b0011110100101000110: color_data = Z;
		19'b0011110100101000111: color_data = Z;
		19'b0011110100101001000: color_data = Z;
		19'b0011110100101001001: color_data = Z;
		19'b0011110100101001010: color_data = Z;
		19'b0011110100101001011: color_data = Z;
		19'b0011110100101001100: color_data = Z;
		19'b0011110100101001101: color_data = Z;
		19'b0011110100101001110: color_data = Z;
		19'b0011110100101001111: color_data = Z;
		19'b0011110100101010000: color_data = Z;
		19'b0011110100101010001: color_data = Z;
		19'b0011110100101010010: color_data = Z;
		19'b0011110100101010011: color_data = Z;
		19'b0011110100101010100: color_data = Z;
		19'b0011110100101010101: color_data = Z;
		19'b0011110100101010110: color_data = Z;
		19'b0011110100101010111: color_data = Z;
		19'b0011110100101011000: color_data = Z;
		19'b0011110100101011001: color_data = Z;
		19'b0011110100101011010: color_data = Z;
		19'b0011110100101011011: color_data = Z;
		19'b0011110100101011100: color_data = Z;
		19'b0011110100101011101: color_data = Z;
		19'b0011110100101011110: color_data = Z;
		19'b0011110100101011111: color_data = Z;
		19'b0011110100101100000: color_data = Z;
		19'b0011110100101100001: color_data = Z;
		19'b0011110100101100010: color_data = Z;
		19'b0011110100101100011: color_data = Z;
		19'b0011110100101100100: color_data = Z;
		19'b0011110100101100101: color_data = Z;
		19'b0011110100101100110: color_data = Z;
		19'b0011110100101100111: color_data = Z;
		19'b0011110100101101000: color_data = Z;
		19'b0011110100101101001: color_data = Z;
		19'b0011110100101101010: color_data = Z;
		19'b0011110100101101011: color_data = Z;
		19'b0011110100101101100: color_data = Z;
		19'b0011110100101101101: color_data = Z;
		19'b0011110100101101110: color_data = Z;
		19'b0011110100101101111: color_data = Z;
		19'b0011110100101110000: color_data = Z;
		19'b0011110100101110001: color_data = Z;
		19'b0011110100101110010: color_data = Z;
		19'b0011110100101110011: color_data = Z;
		19'b0011110100101110100: color_data = Z;
		19'b0011110100101110101: color_data = Z;
		19'b0011110100101110110: color_data = Z;
		19'b0011110100101110111: color_data = Z;
		19'b0011110100101111000: color_data = Z;
		19'b0011110100101111001: color_data = Z;
		19'b0011110100101111010: color_data = Z;
		19'b0011110100101111011: color_data = Z;
		19'b0011110100101111100: color_data = Z;
		19'b0011110100101111101: color_data = Z;
		19'b0011110100101111110: color_data = Z;
		19'b0011110100101111111: color_data = Z;
		19'b0011110100110000000: color_data = Z;
		19'b0011110100110000001: color_data = Z;
		19'b0011110100110000010: color_data = Z;
		19'b0011110100110000011: color_data = Z;
		19'b0011110100110000100: color_data = Z;
		19'b0011110100110000101: color_data = Z;
		19'b0011110100110000110: color_data = Z;
		19'b0011110100110000111: color_data = Z;
		19'b0011110100110001000: color_data = Z;
		19'b0011110100110001001: color_data = Z;
		19'b0011110100110001010: color_data = Z;
		19'b0011110100110001011: color_data = Z;
		19'b0011110100110001100: color_data = Z;
		19'b0011110100111000101: color_data = Z;
		19'b0011110100111000110: color_data = Z;
		19'b0011110100111001001: color_data = Z;
		19'b0011110100111001010: color_data = Z;
		19'b0011110100111001011: color_data = Z;
		19'b0011110100111011010: color_data = Z;
		19'b0011110100111011011: color_data = Z;
		19'b0011110100111011101: color_data = Z;
		19'b0011110100111011110: color_data = Z;
		19'b0011110100111011111: color_data = Z;
		19'b0011110100111100000: color_data = Z;
		19'b0011110110010110001: color_data = Z;
		19'b0011110110010110010: color_data = Z;
		19'b0011110110010110011: color_data = Z;
		19'b0011110110010110100: color_data = Z;
		19'b0011110110010110101: color_data = Z;
		19'b0011110110010110111: color_data = Z;
		19'b0011110110010111000: color_data = Z;
		19'b0011110110010111001: color_data = Z;
		19'b0011110110010111010: color_data = Z;
		19'b0011110110010111011: color_data = Z;
		19'b0011110110010111100: color_data = Z;
		19'b0011110110010111101: color_data = Z;
		19'b0011110110010111110: color_data = Z;
		19'b0011110110010111111: color_data = Z;
		19'b0011110110011000000: color_data = Z;
		19'b0011110110011000001: color_data = Z;
		19'b0011110110011000010: color_data = Z;
		19'b0011110110011000011: color_data = Z;
		19'b0011110110011000100: color_data = Z;
		19'b0011110110011000101: color_data = Z;
		19'b0011110110011000110: color_data = Z;
		19'b0011110110011010001: color_data = Z;
		19'b0011110110011010010: color_data = Z;
		19'b0011110110011010011: color_data = Z;
		19'b0011110110011010100: color_data = Z;
		19'b0011110110011011001: color_data = Z;
		19'b0011110110011011010: color_data = Z;
		19'b0011110110011011011: color_data = Z;
		19'b0011110110011011100: color_data = Z;
		19'b0011110110011011101: color_data = Z;
		19'b0011110110011011110: color_data = Z;
		19'b0011110110011011111: color_data = Z;
		19'b0011110110011100000: color_data = Z;
		19'b0011110110011100001: color_data = Z;
		19'b0011110110011100010: color_data = Z;
		19'b0011110110011100011: color_data = Z;
		19'b0011110110011100100: color_data = Z;
		19'b0011110110011100101: color_data = Z;
		19'b0011110110011100110: color_data = Z;
		19'b0011110110011100111: color_data = Z;
		19'b0011110110011101000: color_data = Z;
		19'b0011110110011101001: color_data = Z;
		19'b0011110110011101010: color_data = Z;
		19'b0011110110011101011: color_data = Z;
		19'b0011110110011101100: color_data = Z;
		19'b0011110110011101101: color_data = Z;
		19'b0011110110011101110: color_data = Z;
		19'b0011110110011101111: color_data = Z;
		19'b0011110110011110000: color_data = Z;
		19'b0011110110011110001: color_data = Z;
		19'b0011110110011110010: color_data = Z;
		19'b0011110110011110011: color_data = Z;
		19'b0011110110011110100: color_data = Z;
		19'b0011110110011110101: color_data = Z;
		19'b0011110110011110110: color_data = Z;
		19'b0011110110011110111: color_data = Z;
		19'b0011110110011111000: color_data = Z;
		19'b0011110110011111001: color_data = Z;
		19'b0011110110011111010: color_data = Z;
		19'b0011110110011111011: color_data = Z;
		19'b0011110110011111100: color_data = Z;
		19'b0011110110011111101: color_data = Z;
		19'b0011110110011111110: color_data = Z;
		19'b0011110110011111111: color_data = Z;
		19'b0011110110100000000: color_data = Z;
		19'b0011110110100000001: color_data = Z;
		19'b0011110110100000010: color_data = Z;
		19'b0011110110100000011: color_data = Z;
		19'b0011110110100000100: color_data = Z;
		19'b0011110110100000101: color_data = Z;
		19'b0011110110100000110: color_data = Z;
		19'b0011110110100000111: color_data = Z;
		19'b0011110110100001000: color_data = Z;
		19'b0011110110100001001: color_data = Z;
		19'b0011110110100001010: color_data = Z;
		19'b0011110110100001011: color_data = Z;
		19'b0011110110100001100: color_data = Z;
		19'b0011110110100001101: color_data = Z;
		19'b0011110110100001110: color_data = Z;
		19'b0011110110100001111: color_data = Z;
		19'b0011110110100010000: color_data = Z;
		19'b0011110110100010001: color_data = Z;
		19'b0011110110100010010: color_data = Z;
		19'b0011110110100010011: color_data = Z;
		19'b0011110110100010100: color_data = Z;
		19'b0011110110100010101: color_data = Z;
		19'b0011110110100010110: color_data = Z;
		19'b0011110110100010111: color_data = Z;
		19'b0011110110100011000: color_data = Z;
		19'b0011110110100011001: color_data = Z;
		19'b0011110110100011010: color_data = Z;
		19'b0011110110100011011: color_data = Z;
		19'b0011110110100011100: color_data = Z;
		19'b0011110110100011101: color_data = Z;
		19'b0011110110100011110: color_data = Z;
		19'b0011110110100011111: color_data = Z;
		19'b0011110110100100000: color_data = Z;
		19'b0011110110100100001: color_data = Z;
		19'b0011110110100100010: color_data = Z;
		19'b0011110110100100011: color_data = Z;
		19'b0011110110100100100: color_data = Z;
		19'b0011110110100100101: color_data = Z;
		19'b0011110110100100110: color_data = Z;
		19'b0011110110100100111: color_data = Z;
		19'b0011110110100101000: color_data = Z;
		19'b0011110110100101001: color_data = Z;
		19'b0011110110100101010: color_data = Z;
		19'b0011110110100101011: color_data = Z;
		19'b0011110110100101100: color_data = Z;
		19'b0011110110100101101: color_data = Z;
		19'b0011110110100101110: color_data = Z;
		19'b0011110110100101111: color_data = Z;
		19'b0011110110100110000: color_data = Z;
		19'b0011110110100110001: color_data = Z;
		19'b0011110110100110010: color_data = Z;
		19'b0011110110100110011: color_data = Z;
		19'b0011110110100110100: color_data = Z;
		19'b0011110110100110101: color_data = Z;
		19'b0011110110100110110: color_data = Z;
		19'b0011110110100110111: color_data = Z;
		19'b0011110110100111000: color_data = Z;
		19'b0011110110100111001: color_data = Z;
		19'b0011110110100111010: color_data = Z;
		19'b0011110110100111011: color_data = Z;
		19'b0011110110100111100: color_data = Z;
		19'b0011110110100111101: color_data = Z;
		19'b0011110110100111110: color_data = Z;
		19'b0011110110100111111: color_data = Z;
		19'b0011110110101000000: color_data = Z;
		19'b0011110110101000001: color_data = Z;
		19'b0011110110101000010: color_data = Z;
		19'b0011110110101000011: color_data = Z;
		19'b0011110110101000100: color_data = Z;
		19'b0011110110101000101: color_data = Z;
		19'b0011110110101000110: color_data = Z;
		19'b0011110110101000111: color_data = Z;
		19'b0011110110101001000: color_data = Z;
		19'b0011110110101001001: color_data = Z;
		19'b0011110110101001010: color_data = Z;
		19'b0011110110101001011: color_data = Z;
		19'b0011110110101001100: color_data = Z;
		19'b0011110110101001101: color_data = Z;
		19'b0011110110101001110: color_data = Z;
		19'b0011110110101001111: color_data = Z;
		19'b0011110110101010000: color_data = Z;
		19'b0011110110101010001: color_data = Z;
		19'b0011110110101010010: color_data = Z;
		19'b0011110110101010011: color_data = Z;
		19'b0011110110101010100: color_data = Z;
		19'b0011110110101010101: color_data = Z;
		19'b0011110110101010110: color_data = Z;
		19'b0011110110101010111: color_data = Z;
		19'b0011110110101011000: color_data = Z;
		19'b0011110110101011001: color_data = Z;
		19'b0011110110101011010: color_data = Z;
		19'b0011110110101011011: color_data = Z;
		19'b0011110110101011100: color_data = Z;
		19'b0011110110101011101: color_data = Z;
		19'b0011110110101011110: color_data = Z;
		19'b0011110110101011111: color_data = Z;
		19'b0011110110101100000: color_data = Z;
		19'b0011110110101100001: color_data = Z;
		19'b0011110110101100010: color_data = Z;
		19'b0011110110101100011: color_data = Z;
		19'b0011110110101100100: color_data = Z;
		19'b0011110110101100101: color_data = Z;
		19'b0011110110101100110: color_data = Z;
		19'b0011110110101100111: color_data = Z;
		19'b0011110110101101000: color_data = Z;
		19'b0011110110101101001: color_data = Z;
		19'b0011110110101101010: color_data = Z;
		19'b0011110110101101011: color_data = Z;
		19'b0011110110101101100: color_data = Z;
		19'b0011110110101101101: color_data = Z;
		19'b0011110110101101110: color_data = Z;
		19'b0011110110101101111: color_data = Z;
		19'b0011110110101110000: color_data = Z;
		19'b0011110110101110001: color_data = Z;
		19'b0011110110101110010: color_data = Z;
		19'b0011110110101110011: color_data = Z;
		19'b0011110110101110100: color_data = Z;
		19'b0011110110101110101: color_data = Z;
		19'b0011110110101110110: color_data = Z;
		19'b0011110110101110111: color_data = Z;
		19'b0011110110101111000: color_data = Z;
		19'b0011110110101111001: color_data = Z;
		19'b0011110110101111010: color_data = Z;
		19'b0011110110101111011: color_data = Z;
		19'b0011110110101111100: color_data = Z;
		19'b0011110110101111101: color_data = Z;
		19'b0011110110101111110: color_data = Z;
		19'b0011110110101111111: color_data = Z;
		19'b0011110110110000000: color_data = Z;
		19'b0011110110110000001: color_data = Z;
		19'b0011110110110000010: color_data = Z;
		19'b0011110110110000011: color_data = Z;
		19'b0011110110110000100: color_data = Z;
		19'b0011110110110000101: color_data = Z;
		19'b0011110110110000110: color_data = Z;
		19'b0011110110110000111: color_data = Z;
		19'b0011110110110001000: color_data = Z;
		19'b0011110110110001001: color_data = Z;
		19'b0011110110110001010: color_data = Z;
		19'b0011110110110001011: color_data = Z;
		19'b0011110110110001100: color_data = Z;
		19'b0011110110111000101: color_data = Z;
		19'b0011110110111000110: color_data = Z;
		19'b0011110110111000111: color_data = Z;
		19'b0011110110111001001: color_data = Z;
		19'b0011110110111001010: color_data = Z;
		19'b0011110110111001011: color_data = Z;
		19'b0011110110111011010: color_data = Z;
		19'b0011110110111011011: color_data = Z;
		19'b0011110110111011100: color_data = Z;
		19'b0011110110111011101: color_data = Z;
		19'b0011110110111011110: color_data = Z;
		19'b0011110110111011111: color_data = Z;
		19'b0011110110111100000: color_data = Z;
		19'b0011111000010110001: color_data = Z;
		19'b0011111000010110010: color_data = Z;
		19'b0011111000010110011: color_data = Z;
		19'b0011111000010111000: color_data = Z;
		19'b0011111000010111001: color_data = Z;
		19'b0011111000010111010: color_data = Z;
		19'b0011111000010111011: color_data = Z;
		19'b0011111000010111100: color_data = Z;
		19'b0011111000010111101: color_data = Z;
		19'b0011111000010111110: color_data = Z;
		19'b0011111000010111111: color_data = Z;
		19'b0011111000011000000: color_data = Z;
		19'b0011111000011000001: color_data = Z;
		19'b0011111000011000010: color_data = Z;
		19'b0011111000011000011: color_data = Z;
		19'b0011111000011000100: color_data = Z;
		19'b0011111000011001111: color_data = Z;
		19'b0011111000011010000: color_data = Z;
		19'b0011111000011010001: color_data = Z;
		19'b0011111000011010111: color_data = Z;
		19'b0011111000011011000: color_data = Z;
		19'b0011111000011011001: color_data = Z;
		19'b0011111000011011010: color_data = Z;
		19'b0011111000011011011: color_data = Z;
		19'b0011111000011011100: color_data = Z;
		19'b0011111000011011101: color_data = Z;
		19'b0011111000011011110: color_data = Z;
		19'b0011111000011011111: color_data = Z;
		19'b0011111000011100000: color_data = Z;
		19'b0011111000011100001: color_data = Z;
		19'b0011111000011100010: color_data = Z;
		19'b0011111000011100011: color_data = Z;
		19'b0011111000011100100: color_data = Z;
		19'b0011111000011100101: color_data = Z;
		19'b0011111000011100110: color_data = Z;
		19'b0011111000011100111: color_data = Z;
		19'b0011111000011101000: color_data = Z;
		19'b0011111000011101001: color_data = Z;
		19'b0011111000011101100: color_data = Z;
		19'b0011111000011101101: color_data = Z;
		19'b0011111000011101110: color_data = Z;
		19'b0011111000011101111: color_data = Z;
		19'b0011111000011110000: color_data = Z;
		19'b0011111000011110001: color_data = Z;
		19'b0011111000011110010: color_data = Z;
		19'b0011111000011110011: color_data = Z;
		19'b0011111000011110100: color_data = Z;
		19'b0011111000011110101: color_data = Z;
		19'b0011111000011110110: color_data = Z;
		19'b0011111000011110111: color_data = Z;
		19'b0011111000011111000: color_data = Z;
		19'b0011111000011111001: color_data = Z;
		19'b0011111000011111010: color_data = Z;
		19'b0011111000011111011: color_data = Z;
		19'b0011111000011111100: color_data = Z;
		19'b0011111000011111101: color_data = Z;
		19'b0011111000011111110: color_data = Z;
		19'b0011111000011111111: color_data = Z;
		19'b0011111000100000000: color_data = Z;
		19'b0011111000100000001: color_data = Z;
		19'b0011111000100000010: color_data = Z;
		19'b0011111000100000011: color_data = Z;
		19'b0011111000100000100: color_data = Z;
		19'b0011111000100000101: color_data = Z;
		19'b0011111000100000110: color_data = Z;
		19'b0011111000100000111: color_data = Z;
		19'b0011111000100001000: color_data = Z;
		19'b0011111000100001001: color_data = Z;
		19'b0011111000100001010: color_data = Z;
		19'b0011111000100001011: color_data = Z;
		19'b0011111000100001100: color_data = Z;
		19'b0011111000100001101: color_data = Z;
		19'b0011111000100001110: color_data = Z;
		19'b0011111000100001111: color_data = Z;
		19'b0011111000100010000: color_data = Z;
		19'b0011111000100010001: color_data = Z;
		19'b0011111000100010010: color_data = Z;
		19'b0011111000100010011: color_data = Z;
		19'b0011111000100010100: color_data = Z;
		19'b0011111000100010101: color_data = Z;
		19'b0011111000100010110: color_data = Z;
		19'b0011111000100010111: color_data = Z;
		19'b0011111000100011000: color_data = Z;
		19'b0011111000100011001: color_data = Z;
		19'b0011111000100011010: color_data = Z;
		19'b0011111000100011011: color_data = Z;
		19'b0011111000100011100: color_data = Z;
		19'b0011111000100011101: color_data = Z;
		19'b0011111000100011110: color_data = Z;
		19'b0011111000100011111: color_data = Z;
		19'b0011111000100100000: color_data = Z;
		19'b0011111000100100001: color_data = Z;
		19'b0011111000100100010: color_data = Z;
		19'b0011111000100100011: color_data = Z;
		19'b0011111000100100100: color_data = Z;
		19'b0011111000100100101: color_data = Z;
		19'b0011111000100100110: color_data = Z;
		19'b0011111000100100111: color_data = Z;
		19'b0011111000100101000: color_data = Z;
		19'b0011111000100101001: color_data = Z;
		19'b0011111000100101010: color_data = Z;
		19'b0011111000100101011: color_data = Z;
		19'b0011111000100101100: color_data = Z;
		19'b0011111000100101101: color_data = Z;
		19'b0011111000100101110: color_data = Z;
		19'b0011111000100101111: color_data = Z;
		19'b0011111000100110000: color_data = Z;
		19'b0011111000100110001: color_data = Z;
		19'b0011111000100110010: color_data = Z;
		19'b0011111000100110011: color_data = Z;
		19'b0011111000100110100: color_data = Z;
		19'b0011111000100110101: color_data = Z;
		19'b0011111000100110110: color_data = Z;
		19'b0011111000100110111: color_data = Z;
		19'b0011111000100111000: color_data = Z;
		19'b0011111000100111001: color_data = Z;
		19'b0011111000100111010: color_data = Z;
		19'b0011111000100111011: color_data = Z;
		19'b0011111000100111100: color_data = Z;
		19'b0011111000100111101: color_data = Z;
		19'b0011111000100111110: color_data = Z;
		19'b0011111000100111111: color_data = Z;
		19'b0011111000101000000: color_data = Z;
		19'b0011111000101000001: color_data = Z;
		19'b0011111000101000010: color_data = Z;
		19'b0011111000101000011: color_data = Z;
		19'b0011111000101000100: color_data = Z;
		19'b0011111000101000101: color_data = Z;
		19'b0011111000101000110: color_data = Z;
		19'b0011111000101000111: color_data = Z;
		19'b0011111000101001000: color_data = Z;
		19'b0011111000101001001: color_data = Z;
		19'b0011111000101001010: color_data = Z;
		19'b0011111000101001011: color_data = Z;
		19'b0011111000101001100: color_data = Z;
		19'b0011111000101001101: color_data = Z;
		19'b0011111000101001110: color_data = Z;
		19'b0011111000101001111: color_data = Z;
		19'b0011111000101010000: color_data = Z;
		19'b0011111000101010001: color_data = Z;
		19'b0011111000101010010: color_data = Z;
		19'b0011111000101010011: color_data = Z;
		19'b0011111000101010100: color_data = Z;
		19'b0011111000101010101: color_data = Z;
		19'b0011111000101010110: color_data = Z;
		19'b0011111000101010111: color_data = Z;
		19'b0011111000101011000: color_data = Z;
		19'b0011111000101011001: color_data = Z;
		19'b0011111000101011010: color_data = Z;
		19'b0011111000101011011: color_data = Z;
		19'b0011111000101011100: color_data = Z;
		19'b0011111000101011101: color_data = Z;
		19'b0011111000101011110: color_data = Z;
		19'b0011111000101011111: color_data = Z;
		19'b0011111000101100000: color_data = Z;
		19'b0011111000101100001: color_data = Z;
		19'b0011111000101100010: color_data = Z;
		19'b0011111000101100011: color_data = Z;
		19'b0011111000101100100: color_data = Z;
		19'b0011111000101100101: color_data = Z;
		19'b0011111000101100110: color_data = Z;
		19'b0011111000101100111: color_data = Z;
		19'b0011111000101101000: color_data = Z;
		19'b0011111000101101001: color_data = Z;
		19'b0011111000101101010: color_data = Z;
		19'b0011111000101101011: color_data = Z;
		19'b0011111000101101100: color_data = Z;
		19'b0011111000101101101: color_data = Z;
		19'b0011111000101101110: color_data = Z;
		19'b0011111000101101111: color_data = Z;
		19'b0011111000101110000: color_data = Z;
		19'b0011111000101110001: color_data = Z;
		19'b0011111000101110010: color_data = Z;
		19'b0011111000101110011: color_data = Z;
		19'b0011111000101110100: color_data = Z;
		19'b0011111000101110101: color_data = Z;
		19'b0011111000101110110: color_data = Z;
		19'b0011111000101110111: color_data = Z;
		19'b0011111000101111000: color_data = Z;
		19'b0011111000101111001: color_data = Z;
		19'b0011111000101111010: color_data = Z;
		19'b0011111000101111011: color_data = Z;
		19'b0011111000101111100: color_data = Z;
		19'b0011111000101111101: color_data = Z;
		19'b0011111000101111110: color_data = Z;
		19'b0011111000101111111: color_data = Z;
		19'b0011111000110000000: color_data = Z;
		19'b0011111000110000001: color_data = Z;
		19'b0011111000110000010: color_data = Z;
		19'b0011111000110000011: color_data = Z;
		19'b0011111000110000100: color_data = Z;
		19'b0011111000110000101: color_data = Z;
		19'b0011111000110000110: color_data = Z;
		19'b0011111000110000111: color_data = Z;
		19'b0011111000110001000: color_data = Z;
		19'b0011111000110001001: color_data = Z;
		19'b0011111000110001010: color_data = Z;
		19'b0011111000110001011: color_data = Z;
		19'b0011111000111000110: color_data = Z;
		19'b0011111000111000111: color_data = Z;
		19'b0011111000111001000: color_data = Z;
		19'b0011111000111001001: color_data = Z;
		19'b0011111000111001010: color_data = Z;
		19'b0011111000111001011: color_data = Z;
		19'b0011111000111001100: color_data = Z;
		19'b0011111000111011010: color_data = Z;
		19'b0011111000111011011: color_data = Z;
		19'b0011111000111011110: color_data = Z;
		19'b0011111000111011111: color_data = Z;
		19'b0011111000111100000: color_data = Z;
		19'b0011111010010110000: color_data = Z;
		19'b0011111010010110001: color_data = Z;
		19'b0011111010010110010: color_data = Z;
		19'b0011111010010110011: color_data = Z;
		19'b0011111010010111000: color_data = Z;
		19'b0011111010010111001: color_data = Z;
		19'b0011111010010111010: color_data = Z;
		19'b0011111010010111011: color_data = Z;
		19'b0011111010010111100: color_data = Z;
		19'b0011111010010111101: color_data = Z;
		19'b0011111010010111110: color_data = Z;
		19'b0011111010010111111: color_data = Z;
		19'b0011111010011000000: color_data = Z;
		19'b0011111010011000001: color_data = Z;
		19'b0011111010011000010: color_data = Z;
		19'b0011111010011001101: color_data = Z;
		19'b0011111010011001110: color_data = Z;
		19'b0011111010011001111: color_data = Z;
		19'b0011111010011010110: color_data = Z;
		19'b0011111010011010111: color_data = Z;
		19'b0011111010011011000: color_data = Z;
		19'b0011111010011011001: color_data = Z;
		19'b0011111010011011010: color_data = Z;
		19'b0011111010011011011: color_data = Z;
		19'b0011111010011011100: color_data = Z;
		19'b0011111010011011101: color_data = Z;
		19'b0011111010011011110: color_data = Z;
		19'b0011111010011011111: color_data = Z;
		19'b0011111010011100000: color_data = Z;
		19'b0011111010011100001: color_data = Z;
		19'b0011111010011100010: color_data = Z;
		19'b0011111010011100011: color_data = Z;
		19'b0011111010011100100: color_data = Z;
		19'b0011111010011100101: color_data = Z;
		19'b0011111010011100110: color_data = Z;
		19'b0011111010011100111: color_data = Z;
		19'b0011111010011101000: color_data = Z;
		19'b0011111010011101101: color_data = Z;
		19'b0011111010011101110: color_data = Z;
		19'b0011111010011101111: color_data = Z;
		19'b0011111010011110000: color_data = Z;
		19'b0011111010011110001: color_data = Z;
		19'b0011111010011110010: color_data = Z;
		19'b0011111010011110011: color_data = Z;
		19'b0011111010011110100: color_data = Z;
		19'b0011111010011110101: color_data = Z;
		19'b0011111010011110110: color_data = Z;
		19'b0011111010011110111: color_data = Z;
		19'b0011111010011111000: color_data = Z;
		19'b0011111010011111001: color_data = Z;
		19'b0011111010011111010: color_data = Z;
		19'b0011111010011111011: color_data = Z;
		19'b0011111010011111100: color_data = Z;
		19'b0011111010011111101: color_data = Z;
		19'b0011111010011111110: color_data = Z;
		19'b0011111010011111111: color_data = Z;
		19'b0011111010100000000: color_data = Z;
		19'b0011111010100000001: color_data = Z;
		19'b0011111010100000010: color_data = Z;
		19'b0011111010100000011: color_data = Z;
		19'b0011111010100000100: color_data = Z;
		19'b0011111010100000101: color_data = Z;
		19'b0011111010100000110: color_data = Z;
		19'b0011111010100000111: color_data = Z;
		19'b0011111010100001000: color_data = Z;
		19'b0011111010100001001: color_data = Z;
		19'b0011111010100001010: color_data = Z;
		19'b0011111010100001011: color_data = Z;
		19'b0011111010100001100: color_data = Z;
		19'b0011111010100001101: color_data = Z;
		19'b0011111010100001110: color_data = Z;
		19'b0011111010100001111: color_data = Z;
		19'b0011111010100010000: color_data = Z;
		19'b0011111010100010001: color_data = Z;
		19'b0011111010100010010: color_data = Z;
		19'b0011111010100010011: color_data = Z;
		19'b0011111010100010100: color_data = Z;
		19'b0011111010100010101: color_data = Z;
		19'b0011111010100010110: color_data = Z;
		19'b0011111010100010111: color_data = Z;
		19'b0011111010100011000: color_data = Z;
		19'b0011111010100011001: color_data = Z;
		19'b0011111010100011010: color_data = Z;
		19'b0011111010100011011: color_data = Z;
		19'b0011111010100011100: color_data = Z;
		19'b0011111010100011101: color_data = Z;
		19'b0011111010100011110: color_data = Z;
		19'b0011111010100011111: color_data = Z;
		19'b0011111010100100000: color_data = Z;
		19'b0011111010100100001: color_data = Z;
		19'b0011111010100100010: color_data = Z;
		19'b0011111010100100011: color_data = Z;
		19'b0011111010100100100: color_data = Z;
		19'b0011111010100100101: color_data = Z;
		19'b0011111010100100110: color_data = Z;
		19'b0011111010100100111: color_data = Z;
		19'b0011111010100101000: color_data = Z;
		19'b0011111010100101001: color_data = Z;
		19'b0011111010100101010: color_data = Z;
		19'b0011111010100101011: color_data = Z;
		19'b0011111010100101100: color_data = Z;
		19'b0011111010100101101: color_data = Z;
		19'b0011111010100101110: color_data = Z;
		19'b0011111010100101111: color_data = Z;
		19'b0011111010100110000: color_data = Z;
		19'b0011111010100110001: color_data = Z;
		19'b0011111010100110010: color_data = Z;
		19'b0011111010100110011: color_data = Z;
		19'b0011111010100110100: color_data = Z;
		19'b0011111010100110101: color_data = Z;
		19'b0011111010100110110: color_data = Z;
		19'b0011111010100110111: color_data = Z;
		19'b0011111010100111000: color_data = Z;
		19'b0011111010100111001: color_data = Z;
		19'b0011111010100111010: color_data = Z;
		19'b0011111010100111011: color_data = Z;
		19'b0011111010100111100: color_data = Z;
		19'b0011111010100111101: color_data = Z;
		19'b0011111010100111110: color_data = Z;
		19'b0011111010100111111: color_data = Z;
		19'b0011111010101000000: color_data = Z;
		19'b0011111010101000001: color_data = Z;
		19'b0011111010101000010: color_data = Z;
		19'b0011111010101000011: color_data = Z;
		19'b0011111010101000100: color_data = Z;
		19'b0011111010101000101: color_data = Z;
		19'b0011111010101000110: color_data = Z;
		19'b0011111010101000111: color_data = Z;
		19'b0011111010101001000: color_data = Z;
		19'b0011111010101001001: color_data = Z;
		19'b0011111010101001010: color_data = Z;
		19'b0011111010101001011: color_data = Z;
		19'b0011111010101001100: color_data = Z;
		19'b0011111010101001101: color_data = Z;
		19'b0011111010101001110: color_data = Z;
		19'b0011111010101001111: color_data = Z;
		19'b0011111010101010000: color_data = Z;
		19'b0011111010101010001: color_data = Z;
		19'b0011111010101010010: color_data = Z;
		19'b0011111010101010011: color_data = Z;
		19'b0011111010101010100: color_data = Z;
		19'b0011111010101010101: color_data = Z;
		19'b0011111010101010110: color_data = Z;
		19'b0011111010101010111: color_data = Z;
		19'b0011111010101011000: color_data = Z;
		19'b0011111010101011001: color_data = Z;
		19'b0011111010101011010: color_data = Z;
		19'b0011111010101011011: color_data = Z;
		19'b0011111010101011100: color_data = Z;
		19'b0011111010101011101: color_data = Z;
		19'b0011111010101011110: color_data = Z;
		19'b0011111010101011111: color_data = Z;
		19'b0011111010101100000: color_data = Z;
		19'b0011111010101100001: color_data = Z;
		19'b0011111010101100010: color_data = Z;
		19'b0011111010101100011: color_data = Z;
		19'b0011111010101100100: color_data = Z;
		19'b0011111010101100101: color_data = Z;
		19'b0011111010101100110: color_data = Z;
		19'b0011111010101100111: color_data = Z;
		19'b0011111010101101000: color_data = Z;
		19'b0011111010101101001: color_data = Z;
		19'b0011111010101101010: color_data = Z;
		19'b0011111010101101011: color_data = Z;
		19'b0011111010101101100: color_data = Z;
		19'b0011111010101101101: color_data = Z;
		19'b0011111010101101110: color_data = Z;
		19'b0011111010101101111: color_data = Z;
		19'b0011111010101110000: color_data = Z;
		19'b0011111010101110001: color_data = Z;
		19'b0011111010101110010: color_data = Z;
		19'b0011111010101110011: color_data = Z;
		19'b0011111010101110100: color_data = Z;
		19'b0011111010101110101: color_data = Z;
		19'b0011111010101110110: color_data = Z;
		19'b0011111010101110111: color_data = Z;
		19'b0011111010101111000: color_data = Z;
		19'b0011111010101111001: color_data = Z;
		19'b0011111010101111010: color_data = Z;
		19'b0011111010101111011: color_data = Z;
		19'b0011111010101111100: color_data = Z;
		19'b0011111010101111101: color_data = Z;
		19'b0011111010101111110: color_data = Z;
		19'b0011111010101111111: color_data = Z;
		19'b0011111010110000000: color_data = Z;
		19'b0011111010110000001: color_data = Z;
		19'b0011111010110000010: color_data = Z;
		19'b0011111010110000011: color_data = Z;
		19'b0011111010110000100: color_data = Z;
		19'b0011111010110000101: color_data = Z;
		19'b0011111010110000110: color_data = Z;
		19'b0011111010110000111: color_data = Z;
		19'b0011111010110001000: color_data = Z;
		19'b0011111010110001001: color_data = Z;
		19'b0011111010110001010: color_data = Z;
		19'b0011111010111000111: color_data = Z;
		19'b0011111010111001000: color_data = Z;
		19'b0011111010111001001: color_data = Z;
		19'b0011111010111001010: color_data = Z;
		19'b0011111010111001011: color_data = Z;
		19'b0011111010111001100: color_data = Z;
		19'b0011111010111011010: color_data = Z;
		19'b0011111010111011011: color_data = Z;
		19'b0011111010111011110: color_data = Z;
		19'b0011111010111011111: color_data = Z;
		19'b0011111010111100000: color_data = Z;
		19'b0011111100010101111: color_data = Z;
		19'b0011111100010110000: color_data = Z;
		19'b0011111100010110001: color_data = Z;
		19'b0011111100010110010: color_data = Z;
		19'b0011111100010110111: color_data = Z;
		19'b0011111100010111000: color_data = Z;
		19'b0011111100010111001: color_data = Z;
		19'b0011111100010111010: color_data = Z;
		19'b0011111100010111011: color_data = Z;
		19'b0011111100010111100: color_data = Z;
		19'b0011111100010111101: color_data = Z;
		19'b0011111100010111110: color_data = Z;
		19'b0011111100010111111: color_data = Z;
		19'b0011111100011001100: color_data = Z;
		19'b0011111100011001101: color_data = Z;
		19'b0011111100011010101: color_data = Z;
		19'b0011111100011010110: color_data = Z;
		19'b0011111100011010111: color_data = Z;
		19'b0011111100011011000: color_data = Z;
		19'b0011111100011011001: color_data = Z;
		19'b0011111100011011010: color_data = Z;
		19'b0011111100011011011: color_data = Z;
		19'b0011111100011011100: color_data = Z;
		19'b0011111100011011101: color_data = Z;
		19'b0011111100011011110: color_data = Z;
		19'b0011111100011011111: color_data = Z;
		19'b0011111100011100000: color_data = Z;
		19'b0011111100011100001: color_data = Z;
		19'b0011111100011100010: color_data = Z;
		19'b0011111100011100011: color_data = Z;
		19'b0011111100011100100: color_data = Z;
		19'b0011111100011100101: color_data = Z;
		19'b0011111100011100110: color_data = Z;
		19'b0011111100011100111: color_data = Z;
		19'b0011111100011101000: color_data = Z;
		19'b0011111100011101001: color_data = Z;
		19'b0011111100011101010: color_data = Z;
		19'b0011111100011101011: color_data = Z;
		19'b0011111100011101100: color_data = Z;
		19'b0011111100011101101: color_data = Z;
		19'b0011111100011101110: color_data = Z;
		19'b0011111100011101111: color_data = Z;
		19'b0011111100011110000: color_data = Z;
		19'b0011111100011110001: color_data = Z;
		19'b0011111100011110010: color_data = Z;
		19'b0011111100011110011: color_data = Z;
		19'b0011111100011110100: color_data = Z;
		19'b0011111100011110101: color_data = Z;
		19'b0011111100011110110: color_data = Z;
		19'b0011111100011110111: color_data = Z;
		19'b0011111100011111000: color_data = Z;
		19'b0011111100011111001: color_data = Z;
		19'b0011111100011111010: color_data = Z;
		19'b0011111100011111011: color_data = Z;
		19'b0011111100011111100: color_data = Z;
		19'b0011111100011111101: color_data = Z;
		19'b0011111100011111110: color_data = Z;
		19'b0011111100011111111: color_data = Z;
		19'b0011111100100000000: color_data = Z;
		19'b0011111100100000001: color_data = Z;
		19'b0011111100100000010: color_data = Z;
		19'b0011111100100000011: color_data = Z;
		19'b0011111100100000100: color_data = Z;
		19'b0011111100100000101: color_data = Z;
		19'b0011111100100000110: color_data = Z;
		19'b0011111100100000111: color_data = Z;
		19'b0011111100100001000: color_data = Z;
		19'b0011111100100001001: color_data = Z;
		19'b0011111100100001010: color_data = Z;
		19'b0011111100100001011: color_data = Z;
		19'b0011111100100001100: color_data = Z;
		19'b0011111100100001101: color_data = Z;
		19'b0011111100100001110: color_data = Z;
		19'b0011111100100001111: color_data = Z;
		19'b0011111100100010000: color_data = Z;
		19'b0011111100100010001: color_data = Z;
		19'b0011111100100010010: color_data = Z;
		19'b0011111100100010011: color_data = Z;
		19'b0011111100100010100: color_data = Z;
		19'b0011111100100010101: color_data = Z;
		19'b0011111100100010110: color_data = Z;
		19'b0011111100100010111: color_data = Z;
		19'b0011111100100011000: color_data = Z;
		19'b0011111100100011001: color_data = Z;
		19'b0011111100100011010: color_data = Z;
		19'b0011111100100011011: color_data = Z;
		19'b0011111100100011100: color_data = Z;
		19'b0011111100100011101: color_data = Z;
		19'b0011111100100011110: color_data = Z;
		19'b0011111100100011111: color_data = Z;
		19'b0011111100100100000: color_data = Z;
		19'b0011111100100100001: color_data = Z;
		19'b0011111100100100010: color_data = Z;
		19'b0011111100100100011: color_data = Z;
		19'b0011111100100100100: color_data = Z;
		19'b0011111100100100101: color_data = Z;
		19'b0011111100100100110: color_data = Z;
		19'b0011111100100100111: color_data = Z;
		19'b0011111100100101000: color_data = Z;
		19'b0011111100100101001: color_data = Z;
		19'b0011111100100101010: color_data = Z;
		19'b0011111100100101011: color_data = Z;
		19'b0011111100100101100: color_data = Z;
		19'b0011111100100101101: color_data = Z;
		19'b0011111100100101110: color_data = Z;
		19'b0011111100100101111: color_data = Z;
		19'b0011111100100110000: color_data = Z;
		19'b0011111100100110001: color_data = Z;
		19'b0011111100100110010: color_data = Z;
		19'b0011111100100110011: color_data = Z;
		19'b0011111100100110100: color_data = Z;
		19'b0011111100100110101: color_data = Z;
		19'b0011111100100110110: color_data = Z;
		19'b0011111100100110111: color_data = Z;
		19'b0011111100100111000: color_data = Z;
		19'b0011111100100111001: color_data = Z;
		19'b0011111100100111010: color_data = Z;
		19'b0011111100100111011: color_data = Z;
		19'b0011111100100111100: color_data = Z;
		19'b0011111100100111101: color_data = Z;
		19'b0011111100100111110: color_data = Z;
		19'b0011111100100111111: color_data = Z;
		19'b0011111100101000000: color_data = Z;
		19'b0011111100101000001: color_data = Z;
		19'b0011111100101000010: color_data = Z;
		19'b0011111100101000011: color_data = Z;
		19'b0011111100101000100: color_data = Z;
		19'b0011111100101000101: color_data = Z;
		19'b0011111100101000110: color_data = Z;
		19'b0011111100101000111: color_data = Z;
		19'b0011111100101001000: color_data = Z;
		19'b0011111100101001001: color_data = Z;
		19'b0011111100101001010: color_data = Z;
		19'b0011111100101001011: color_data = Z;
		19'b0011111100101001100: color_data = Z;
		19'b0011111100101001101: color_data = Z;
		19'b0011111100101001110: color_data = Z;
		19'b0011111100101001111: color_data = Z;
		19'b0011111100101010000: color_data = Z;
		19'b0011111100101010001: color_data = Z;
		19'b0011111100101010010: color_data = Z;
		19'b0011111100101010011: color_data = Z;
		19'b0011111100101010100: color_data = Z;
		19'b0011111100101010101: color_data = Z;
		19'b0011111100101010110: color_data = Z;
		19'b0011111100101010111: color_data = Z;
		19'b0011111100101011000: color_data = Z;
		19'b0011111100101011001: color_data = Z;
		19'b0011111100101011010: color_data = Z;
		19'b0011111100101011011: color_data = Z;
		19'b0011111100101011100: color_data = Z;
		19'b0011111100101011101: color_data = Z;
		19'b0011111100101011110: color_data = Z;
		19'b0011111100101011111: color_data = Z;
		19'b0011111100101100000: color_data = Z;
		19'b0011111100101100001: color_data = Z;
		19'b0011111100101100010: color_data = Z;
		19'b0011111100101100011: color_data = Z;
		19'b0011111100101100100: color_data = Z;
		19'b0011111100101100101: color_data = Z;
		19'b0011111100101100110: color_data = Z;
		19'b0011111100101100111: color_data = Z;
		19'b0011111100101101000: color_data = Z;
		19'b0011111100101101001: color_data = Z;
		19'b0011111100101101010: color_data = Z;
		19'b0011111100101101011: color_data = Z;
		19'b0011111100101101100: color_data = Z;
		19'b0011111100101101101: color_data = Z;
		19'b0011111100101101110: color_data = Z;
		19'b0011111100101101111: color_data = Z;
		19'b0011111100101110000: color_data = Z;
		19'b0011111100101110001: color_data = Z;
		19'b0011111100101110010: color_data = Z;
		19'b0011111100101110011: color_data = Z;
		19'b0011111100101110100: color_data = Z;
		19'b0011111100101110101: color_data = Z;
		19'b0011111100101110110: color_data = Z;
		19'b0011111100101110111: color_data = Z;
		19'b0011111100101111000: color_data = Z;
		19'b0011111100101111001: color_data = Z;
		19'b0011111100101111010: color_data = Z;
		19'b0011111100101111011: color_data = Z;
		19'b0011111100101111100: color_data = Z;
		19'b0011111100101111101: color_data = Z;
		19'b0011111100101111110: color_data = Z;
		19'b0011111100101111111: color_data = Z;
		19'b0011111100110000000: color_data = Z;
		19'b0011111100110000001: color_data = Z;
		19'b0011111100110000010: color_data = Z;
		19'b0011111100110000011: color_data = Z;
		19'b0011111100110000100: color_data = Z;
		19'b0011111100110000101: color_data = Z;
		19'b0011111100110000110: color_data = Z;
		19'b0011111100110000111: color_data = Z;
		19'b0011111100110001000: color_data = Z;
		19'b0011111100110001001: color_data = Z;
		19'b0011111100111001000: color_data = Z;
		19'b0011111100111001001: color_data = Z;
		19'b0011111100111001010: color_data = Z;
		19'b0011111100111001011: color_data = Z;
		19'b0011111100111001100: color_data = Z;
		19'b0011111100111001101: color_data = Z;
		19'b0011111100111001110: color_data = Z;
		19'b0011111100111011010: color_data = Z;
		19'b0011111100111011011: color_data = Z;
		19'b0011111100111011110: color_data = Z;
		19'b0011111100111011111: color_data = Z;
		19'b0011111100111100000: color_data = Z;
		19'b0011111100111100001: color_data = Z;
		19'b0011111110010101100: color_data = Z;
		19'b0011111110010101101: color_data = Z;
		19'b0011111110010101110: color_data = Z;
		19'b0011111110010101111: color_data = Z;
		19'b0011111110010110000: color_data = Z;
		19'b0011111110010110001: color_data = Z;
		19'b0011111110010110111: color_data = Z;
		19'b0011111110010111000: color_data = Z;
		19'b0011111110010111001: color_data = Z;
		19'b0011111110010111010: color_data = Z;
		19'b0011111110010111011: color_data = Z;
		19'b0011111110010111100: color_data = Z;
		19'b0011111110010111101: color_data = Z;
		19'b0011111110011001010: color_data = Z;
		19'b0011111110011001011: color_data = Z;
		19'b0011111110011010011: color_data = Z;
		19'b0011111110011010100: color_data = Z;
		19'b0011111110011010101: color_data = Z;
		19'b0011111110011010110: color_data = Z;
		19'b0011111110011010111: color_data = Z;
		19'b0011111110011011000: color_data = Z;
		19'b0011111110011011001: color_data = Z;
		19'b0011111110011011010: color_data = Z;
		19'b0011111110011011011: color_data = Z;
		19'b0011111110011011101: color_data = Z;
		19'b0011111110011011110: color_data = Z;
		19'b0011111110011011111: color_data = Z;
		19'b0011111110011100000: color_data = Z;
		19'b0011111110011100001: color_data = Z;
		19'b0011111110011100010: color_data = Z;
		19'b0011111110011100101: color_data = Z;
		19'b0011111110011100110: color_data = Z;
		19'b0011111110011100111: color_data = Z;
		19'b0011111110011101000: color_data = Z;
		19'b0011111110011101001: color_data = Z;
		19'b0011111110011101010: color_data = Z;
		19'b0011111110011101011: color_data = Z;
		19'b0011111110011101100: color_data = Z;
		19'b0011111110011101101: color_data = Z;
		19'b0011111110011101110: color_data = Z;
		19'b0011111110011101111: color_data = Z;
		19'b0011111110011110000: color_data = Z;
		19'b0011111110011110001: color_data = Z;
		19'b0011111110011110010: color_data = Z;
		19'b0011111110011110011: color_data = Z;
		19'b0011111110011110100: color_data = Z;
		19'b0011111110011110101: color_data = Z;
		19'b0011111110011110110: color_data = Z;
		19'b0011111110011110111: color_data = Z;
		19'b0011111110011111000: color_data = Z;
		19'b0011111110011111001: color_data = Z;
		19'b0011111110011111010: color_data = Z;
		19'b0011111110011111011: color_data = Z;
		19'b0011111110011111100: color_data = Z;
		19'b0011111110011111101: color_data = Z;
		19'b0011111110011111110: color_data = Z;
		19'b0011111110011111111: color_data = Z;
		19'b0011111110100000000: color_data = Z;
		19'b0011111110100000001: color_data = Z;
		19'b0011111110100000010: color_data = Z;
		19'b0011111110100000011: color_data = Z;
		19'b0011111110100000100: color_data = Z;
		19'b0011111110100000101: color_data = Z;
		19'b0011111110100000110: color_data = Z;
		19'b0011111110100000111: color_data = Z;
		19'b0011111110100001000: color_data = Z;
		19'b0011111110100001001: color_data = Z;
		19'b0011111110100001010: color_data = Z;
		19'b0011111110100001011: color_data = Z;
		19'b0011111110100001100: color_data = Z;
		19'b0011111110100001101: color_data = Z;
		19'b0011111110100001110: color_data = Z;
		19'b0011111110100001111: color_data = Z;
		19'b0011111110100010000: color_data = Z;
		19'b0011111110100010001: color_data = Z;
		19'b0011111110100010010: color_data = Z;
		19'b0011111110100010011: color_data = Z;
		19'b0011111110100010100: color_data = Z;
		19'b0011111110100010101: color_data = Z;
		19'b0011111110100010110: color_data = Z;
		19'b0011111110100010111: color_data = Z;
		19'b0011111110100011000: color_data = Z;
		19'b0011111110100011001: color_data = Z;
		19'b0011111110100011010: color_data = Z;
		19'b0011111110100011011: color_data = Z;
		19'b0011111110100011100: color_data = Z;
		19'b0011111110100011101: color_data = Z;
		19'b0011111110100011110: color_data = Z;
		19'b0011111110100011111: color_data = Z;
		19'b0011111110100100000: color_data = Z;
		19'b0011111110100100001: color_data = Z;
		19'b0011111110100100010: color_data = Z;
		19'b0011111110100100011: color_data = Z;
		19'b0011111110100100100: color_data = Z;
		19'b0011111110100100101: color_data = Z;
		19'b0011111110100100110: color_data = Z;
		19'b0011111110100100111: color_data = Z;
		19'b0011111110100101000: color_data = Z;
		19'b0011111110100101001: color_data = Z;
		19'b0011111110100101010: color_data = Z;
		19'b0011111110100101011: color_data = Z;
		19'b0011111110100101100: color_data = Z;
		19'b0011111110100101101: color_data = Z;
		19'b0011111110100101110: color_data = Z;
		19'b0011111110100101111: color_data = Z;
		19'b0011111110100110000: color_data = Z;
		19'b0011111110100110001: color_data = Z;
		19'b0011111110100110010: color_data = Z;
		19'b0011111110100110011: color_data = Z;
		19'b0011111110100110100: color_data = Z;
		19'b0011111110100110101: color_data = Z;
		19'b0011111110100110110: color_data = Z;
		19'b0011111110100110111: color_data = Z;
		19'b0011111110100111000: color_data = Z;
		19'b0011111110100111001: color_data = Z;
		19'b0011111110100111010: color_data = Z;
		19'b0011111110100111011: color_data = Z;
		19'b0011111110100111100: color_data = Z;
		19'b0011111110100111101: color_data = Z;
		19'b0011111110100111110: color_data = Z;
		19'b0011111110100111111: color_data = Z;
		19'b0011111110101000000: color_data = Z;
		19'b0011111110101000001: color_data = Z;
		19'b0011111110101000010: color_data = Z;
		19'b0011111110101000011: color_data = Z;
		19'b0011111110101000100: color_data = Z;
		19'b0011111110101000101: color_data = Z;
		19'b0011111110101000110: color_data = Z;
		19'b0011111110101000111: color_data = Z;
		19'b0011111110101001000: color_data = Z;
		19'b0011111110101001001: color_data = Z;
		19'b0011111110101001010: color_data = Z;
		19'b0011111110101001011: color_data = Z;
		19'b0011111110101001100: color_data = Z;
		19'b0011111110101001101: color_data = Z;
		19'b0011111110101001110: color_data = Z;
		19'b0011111110101001111: color_data = Z;
		19'b0011111110101010000: color_data = Z;
		19'b0011111110101010001: color_data = Z;
		19'b0011111110101010010: color_data = Z;
		19'b0011111110101010011: color_data = Z;
		19'b0011111110101010100: color_data = Z;
		19'b0011111110101010101: color_data = Z;
		19'b0011111110101010110: color_data = Z;
		19'b0011111110101010111: color_data = Z;
		19'b0011111110101011000: color_data = Z;
		19'b0011111110101011001: color_data = Z;
		19'b0011111110101011010: color_data = Z;
		19'b0011111110101011011: color_data = Z;
		19'b0011111110101011100: color_data = Z;
		19'b0011111110101011101: color_data = Z;
		19'b0011111110101011110: color_data = Z;
		19'b0011111110101011111: color_data = Z;
		19'b0011111110101100000: color_data = Z;
		19'b0011111110101100001: color_data = Z;
		19'b0011111110101100010: color_data = Z;
		19'b0011111110101100011: color_data = Z;
		19'b0011111110101100100: color_data = Z;
		19'b0011111110101100101: color_data = Z;
		19'b0011111110101100110: color_data = Z;
		19'b0011111110101100111: color_data = Z;
		19'b0011111110101101000: color_data = Z;
		19'b0011111110101101001: color_data = Z;
		19'b0011111110101101010: color_data = Z;
		19'b0011111110101101011: color_data = Z;
		19'b0011111110101101100: color_data = Z;
		19'b0011111110101101101: color_data = Z;
		19'b0011111110101101110: color_data = Z;
		19'b0011111110101101111: color_data = Z;
		19'b0011111110101110000: color_data = Z;
		19'b0011111110101110001: color_data = Z;
		19'b0011111110101110010: color_data = Z;
		19'b0011111110101110011: color_data = Z;
		19'b0011111110101110100: color_data = Z;
		19'b0011111110101110101: color_data = Z;
		19'b0011111110101110110: color_data = Z;
		19'b0011111110101110111: color_data = Z;
		19'b0011111110101111000: color_data = Z;
		19'b0011111110101111001: color_data = Z;
		19'b0011111110101111010: color_data = Z;
		19'b0011111110101111011: color_data = Z;
		19'b0011111110101111100: color_data = Z;
		19'b0011111110101111101: color_data = Z;
		19'b0011111110101111110: color_data = Z;
		19'b0011111110101111111: color_data = Z;
		19'b0011111110110000000: color_data = Z;
		19'b0011111110110000001: color_data = Z;
		19'b0011111110110000010: color_data = Z;
		19'b0011111110110000011: color_data = Z;
		19'b0011111110110000100: color_data = Z;
		19'b0011111110110000101: color_data = Z;
		19'b0011111110110000110: color_data = Z;
		19'b0011111110110000111: color_data = Z;
		19'b0011111110110001000: color_data = Z;
		19'b0011111110110001001: color_data = Z;
		19'b0011111110111001000: color_data = Z;
		19'b0011111110111001001: color_data = Z;
		19'b0011111110111001010: color_data = Z;
		19'b0011111110111001011: color_data = Z;
		19'b0011111110111001100: color_data = Z;
		19'b0011111110111001101: color_data = Z;
		19'b0011111110111001110: color_data = Z;
		19'b0011111110111001111: color_data = Z;
		19'b0011111110111011010: color_data = Z;
		19'b0011111110111011011: color_data = Z;
		19'b0011111110111011100: color_data = Z;
		19'b0011111110111011111: color_data = Z;
		19'b0011111110111100000: color_data = Z;
		19'b0011111110111100001: color_data = Z;
		19'b0100000000010101011: color_data = Z;
		19'b0100000000010101100: color_data = Z;
		19'b0100000000010101101: color_data = Z;
		19'b0100000000010101110: color_data = Z;
		19'b0100000000010101111: color_data = Z;
		19'b0100000000010110000: color_data = Z;
		19'b0100000000010110110: color_data = Z;
		19'b0100000000010110111: color_data = Z;
		19'b0100000000010111000: color_data = Z;
		19'b0100000000010111001: color_data = Z;
		19'b0100000000010111010: color_data = Z;
		19'b0100000000010111011: color_data = Z;
		19'b0100000000010111100: color_data = Z;
		19'b0100000000011001000: color_data = Z;
		19'b0100000000011001001: color_data = Z;
		19'b0100000000011010001: color_data = Z;
		19'b0100000000011010010: color_data = Z;
		19'b0100000000011010011: color_data = Z;
		19'b0100000000011010100: color_data = Z;
		19'b0100000000011010101: color_data = Z;
		19'b0100000000011010110: color_data = Z;
		19'b0100000000011010111: color_data = Z;
		19'b0100000000011011000: color_data = Z;
		19'b0100000000011011001: color_data = Z;
		19'b0100000000011011010: color_data = Z;
		19'b0100000000011011110: color_data = Z;
		19'b0100000000011011111: color_data = Z;
		19'b0100000000011100101: color_data = Z;
		19'b0100000000011100110: color_data = Z;
		19'b0100000000011100111: color_data = Z;
		19'b0100000000011101000: color_data = Z;
		19'b0100000000011101001: color_data = Z;
		19'b0100000000011101010: color_data = Z;
		19'b0100000000011101011: color_data = Z;
		19'b0100000000011101100: color_data = Z;
		19'b0100000000011101101: color_data = Z;
		19'b0100000000011101110: color_data = Z;
		19'b0100000000011101111: color_data = Z;
		19'b0100000000011110000: color_data = Z;
		19'b0100000000011110001: color_data = Z;
		19'b0100000000011110010: color_data = Z;
		19'b0100000000011110011: color_data = Z;
		19'b0100000000011110100: color_data = Z;
		19'b0100000000011110101: color_data = Z;
		19'b0100000000011110110: color_data = Z;
		19'b0100000000011110111: color_data = Z;
		19'b0100000000011111000: color_data = Z;
		19'b0100000000011111001: color_data = Z;
		19'b0100000000011111010: color_data = Z;
		19'b0100000000011111011: color_data = Z;
		19'b0100000000011111100: color_data = Z;
		19'b0100000000011111101: color_data = Z;
		19'b0100000000011111110: color_data = Z;
		19'b0100000000011111111: color_data = Z;
		19'b0100000000100000000: color_data = Z;
		19'b0100000000100000001: color_data = Z;
		19'b0100000000100000010: color_data = Z;
		19'b0100000000100000011: color_data = Z;
		19'b0100000000100000100: color_data = Z;
		19'b0100000000100000101: color_data = Z;
		19'b0100000000100000110: color_data = Z;
		19'b0100000000100000111: color_data = Z;
		19'b0100000000100001000: color_data = Z;
		19'b0100000000100001001: color_data = Z;
		19'b0100000000100001010: color_data = Z;
		19'b0100000000100001011: color_data = Z;
		19'b0100000000100001100: color_data = Z;
		19'b0100000000100001101: color_data = Z;
		19'b0100000000100001110: color_data = Z;
		19'b0100000000100001111: color_data = Z;
		19'b0100000000100010000: color_data = Z;
		19'b0100000000100010001: color_data = Z;
		19'b0100000000100010010: color_data = Z;
		19'b0100000000100010011: color_data = Z;
		19'b0100000000100010100: color_data = Z;
		19'b0100000000100010101: color_data = Z;
		19'b0100000000100010110: color_data = Z;
		19'b0100000000100010111: color_data = Z;
		19'b0100000000100011000: color_data = Z;
		19'b0100000000100011001: color_data = Z;
		19'b0100000000100011010: color_data = Z;
		19'b0100000000100011011: color_data = Z;
		19'b0100000000100011100: color_data = Z;
		19'b0100000000100011101: color_data = Z;
		19'b0100000000100011110: color_data = Z;
		19'b0100000000100011111: color_data = Z;
		19'b0100000000100100000: color_data = Z;
		19'b0100000000100100001: color_data = Z;
		19'b0100000000100100010: color_data = Z;
		19'b0100000000100100011: color_data = Z;
		19'b0100000000100100100: color_data = Z;
		19'b0100000000100100101: color_data = Z;
		19'b0100000000100100110: color_data = Z;
		19'b0100000000100100111: color_data = Z;
		19'b0100000000100101000: color_data = Z;
		19'b0100000000100101001: color_data = Z;
		19'b0100000000100101010: color_data = Z;
		19'b0100000000100101011: color_data = Z;
		19'b0100000000100101100: color_data = Z;
		19'b0100000000100101101: color_data = Z;
		19'b0100000000100101110: color_data = Z;
		19'b0100000000100101111: color_data = Z;
		19'b0100000000100110000: color_data = Z;
		19'b0100000000100110001: color_data = Z;
		19'b0100000000100110010: color_data = Z;
		19'b0100000000100110011: color_data = Z;
		19'b0100000000100110100: color_data = Z;
		19'b0100000000100110101: color_data = Z;
		19'b0100000000100110110: color_data = Z;
		19'b0100000000100110111: color_data = Z;
		19'b0100000000100111000: color_data = Z;
		19'b0100000000100111001: color_data = Z;
		19'b0100000000100111010: color_data = Z;
		19'b0100000000100111011: color_data = Z;
		19'b0100000000100111100: color_data = Z;
		19'b0100000000100111101: color_data = Z;
		19'b0100000000100111110: color_data = Z;
		19'b0100000000100111111: color_data = Z;
		19'b0100000000101000000: color_data = Z;
		19'b0100000000101000001: color_data = Z;
		19'b0100000000101000010: color_data = Z;
		19'b0100000000101000011: color_data = Z;
		19'b0100000000101000100: color_data = Z;
		19'b0100000000101000101: color_data = Z;
		19'b0100000000101000110: color_data = Z;
		19'b0100000000101000111: color_data = Z;
		19'b0100000000101001000: color_data = Z;
		19'b0100000000101001001: color_data = Z;
		19'b0100000000101001010: color_data = Z;
		19'b0100000000101001011: color_data = Z;
		19'b0100000000101001100: color_data = Z;
		19'b0100000000101001101: color_data = Z;
		19'b0100000000101001110: color_data = Z;
		19'b0100000000101001111: color_data = Z;
		19'b0100000000101010000: color_data = Z;
		19'b0100000000101010001: color_data = Z;
		19'b0100000000101010010: color_data = Z;
		19'b0100000000101010011: color_data = Z;
		19'b0100000000101010100: color_data = Z;
		19'b0100000000101010101: color_data = Z;
		19'b0100000000101010110: color_data = Z;
		19'b0100000000101010111: color_data = Z;
		19'b0100000000101011000: color_data = Z;
		19'b0100000000101011001: color_data = Z;
		19'b0100000000101011010: color_data = Z;
		19'b0100000000101011011: color_data = Z;
		19'b0100000000101011100: color_data = Z;
		19'b0100000000101011101: color_data = Z;
		19'b0100000000101011110: color_data = Z;
		19'b0100000000101011111: color_data = Z;
		19'b0100000000101100000: color_data = Z;
		19'b0100000000101100001: color_data = Z;
		19'b0100000000101100010: color_data = Z;
		19'b0100000000101100011: color_data = Z;
		19'b0100000000101100100: color_data = Z;
		19'b0100000000101100101: color_data = Z;
		19'b0100000000101100110: color_data = Z;
		19'b0100000000101100111: color_data = Z;
		19'b0100000000101101000: color_data = Z;
		19'b0100000000101101001: color_data = Z;
		19'b0100000000101101010: color_data = Z;
		19'b0100000000101101011: color_data = Z;
		19'b0100000000101101100: color_data = Z;
		19'b0100000000101101101: color_data = Z;
		19'b0100000000101101110: color_data = Z;
		19'b0100000000101101111: color_data = Z;
		19'b0100000000101110000: color_data = Z;
		19'b0100000000101110001: color_data = Z;
		19'b0100000000101110010: color_data = Z;
		19'b0100000000101110011: color_data = Z;
		19'b0100000000101110100: color_data = Z;
		19'b0100000000101110101: color_data = Z;
		19'b0100000000101110110: color_data = Z;
		19'b0100000000101110111: color_data = Z;
		19'b0100000000101111000: color_data = Z;
		19'b0100000000101111001: color_data = Z;
		19'b0100000000101111010: color_data = Z;
		19'b0100000000101111011: color_data = Z;
		19'b0100000000101111100: color_data = Z;
		19'b0100000000101111101: color_data = Z;
		19'b0100000000101111110: color_data = Z;
		19'b0100000000101111111: color_data = Z;
		19'b0100000000110000000: color_data = Z;
		19'b0100000000110000001: color_data = Z;
		19'b0100000000110000010: color_data = Z;
		19'b0100000000110000011: color_data = Z;
		19'b0100000000110000100: color_data = Z;
		19'b0100000000110000101: color_data = Z;
		19'b0100000000110000110: color_data = Z;
		19'b0100000000110000111: color_data = Z;
		19'b0100000000111001100: color_data = Z;
		19'b0100000000111001101: color_data = Z;
		19'b0100000000111001110: color_data = Z;
		19'b0100000000111001111: color_data = Z;
		19'b0100000000111010000: color_data = Z;
		19'b0100000000111010010: color_data = Z;
		19'b0100000000111010011: color_data = Z;
		19'b0100000000111011010: color_data = Z;
		19'b0100000000111011011: color_data = Z;
		19'b0100000000111011100: color_data = Z;
		19'b0100000000111100000: color_data = Z;
		19'b0100000000111100001: color_data = Z;
		19'b0100000010010101011: color_data = Z;
		19'b0100000010010101100: color_data = Z;
		19'b0100000010010101101: color_data = Z;
		19'b0100000010010101110: color_data = Z;
		19'b0100000010010101111: color_data = Z;
		19'b0100000010010110101: color_data = Z;
		19'b0100000010010110110: color_data = Z;
		19'b0100000010010110111: color_data = Z;
		19'b0100000010010111000: color_data = Z;
		19'b0100000010010111001: color_data = Z;
		19'b0100000010010111010: color_data = Z;
		19'b0100000010010111011: color_data = Z;
		19'b0100000010010111100: color_data = Z;
		19'b0100000010011001111: color_data = Z;
		19'b0100000010011010000: color_data = Z;
		19'b0100000010011010001: color_data = Z;
		19'b0100000010011010010: color_data = Z;
		19'b0100000010011010011: color_data = Z;
		19'b0100000010011010100: color_data = Z;
		19'b0100000010011010101: color_data = Z;
		19'b0100000010011010110: color_data = Z;
		19'b0100000010011010111: color_data = Z;
		19'b0100000010011011000: color_data = Z;
		19'b0100000010011100110: color_data = Z;
		19'b0100000010011100111: color_data = Z;
		19'b0100000010011101000: color_data = Z;
		19'b0100000010011101001: color_data = Z;
		19'b0100000010011101010: color_data = Z;
		19'b0100000010011101011: color_data = Z;
		19'b0100000010011101100: color_data = Z;
		19'b0100000010011101101: color_data = Z;
		19'b0100000010011101110: color_data = Z;
		19'b0100000010011101111: color_data = Z;
		19'b0100000010011110000: color_data = Z;
		19'b0100000010011110001: color_data = Z;
		19'b0100000010011110010: color_data = Z;
		19'b0100000010011110011: color_data = Z;
		19'b0100000010011110100: color_data = Z;
		19'b0100000010011110101: color_data = Z;
		19'b0100000010011110110: color_data = Z;
		19'b0100000010011110111: color_data = Z;
		19'b0100000010011111000: color_data = Z;
		19'b0100000010011111001: color_data = Z;
		19'b0100000010011111010: color_data = Z;
		19'b0100000010011111011: color_data = Z;
		19'b0100000010011111100: color_data = Z;
		19'b0100000010011111101: color_data = Z;
		19'b0100000010011111110: color_data = Z;
		19'b0100000010011111111: color_data = Z;
		19'b0100000010100000000: color_data = Z;
		19'b0100000010100000001: color_data = Z;
		19'b0100000010100000010: color_data = Z;
		19'b0100000010100000011: color_data = Z;
		19'b0100000010100000100: color_data = Z;
		19'b0100000010100000101: color_data = Z;
		19'b0100000010100000110: color_data = Z;
		19'b0100000010100000111: color_data = Z;
		19'b0100000010100001000: color_data = Z;
		19'b0100000010100001001: color_data = Z;
		19'b0100000010100001010: color_data = Z;
		19'b0100000010100001011: color_data = Z;
		19'b0100000010100001100: color_data = Z;
		19'b0100000010100001101: color_data = Z;
		19'b0100000010100001110: color_data = Z;
		19'b0100000010100001111: color_data = Z;
		19'b0100000010100010000: color_data = Z;
		19'b0100000010100010001: color_data = Z;
		19'b0100000010100010010: color_data = Z;
		19'b0100000010100010011: color_data = Z;
		19'b0100000010100010100: color_data = Z;
		19'b0100000010100010101: color_data = Z;
		19'b0100000010100010110: color_data = Z;
		19'b0100000010100010111: color_data = Z;
		19'b0100000010100011000: color_data = Z;
		19'b0100000010100011001: color_data = Z;
		19'b0100000010100011010: color_data = Z;
		19'b0100000010100011011: color_data = Z;
		19'b0100000010100011100: color_data = Z;
		19'b0100000010100011101: color_data = Z;
		19'b0100000010100011110: color_data = Z;
		19'b0100000010100011111: color_data = Z;
		19'b0100000010100100000: color_data = Z;
		19'b0100000010100100001: color_data = Z;
		19'b0100000010100100010: color_data = Z;
		19'b0100000010100100011: color_data = Z;
		19'b0100000010100100100: color_data = Z;
		19'b0100000010100100101: color_data = Z;
		19'b0100000010100100110: color_data = Z;
		19'b0100000010100100111: color_data = Z;
		19'b0100000010100101000: color_data = Z;
		19'b0100000010100101001: color_data = Z;
		19'b0100000010100101010: color_data = Z;
		19'b0100000010100101011: color_data = Z;
		19'b0100000010100101100: color_data = Z;
		19'b0100000010100101101: color_data = Z;
		19'b0100000010100101110: color_data = Z;
		19'b0100000010100101111: color_data = Z;
		19'b0100000010100110000: color_data = Z;
		19'b0100000010100110001: color_data = Z;
		19'b0100000010100110010: color_data = Z;
		19'b0100000010100110011: color_data = Z;
		19'b0100000010100110100: color_data = Z;
		19'b0100000010100110101: color_data = Z;
		19'b0100000010100110110: color_data = Z;
		19'b0100000010100110111: color_data = Z;
		19'b0100000010100111000: color_data = Z;
		19'b0100000010100111001: color_data = Z;
		19'b0100000010100111010: color_data = Z;
		19'b0100000010100111011: color_data = Z;
		19'b0100000010100111100: color_data = Z;
		19'b0100000010100111101: color_data = Z;
		19'b0100000010100111110: color_data = Z;
		19'b0100000010100111111: color_data = Z;
		19'b0100000010101000000: color_data = Z;
		19'b0100000010101000001: color_data = Z;
		19'b0100000010101000010: color_data = Z;
		19'b0100000010101000011: color_data = Z;
		19'b0100000010101000100: color_data = Z;
		19'b0100000010101000101: color_data = Z;
		19'b0100000010101000110: color_data = Z;
		19'b0100000010101000111: color_data = Z;
		19'b0100000010101001000: color_data = Z;
		19'b0100000010101001001: color_data = Z;
		19'b0100000010101001010: color_data = Z;
		19'b0100000010101001011: color_data = Z;
		19'b0100000010101001100: color_data = Z;
		19'b0100000010101001101: color_data = Z;
		19'b0100000010101001110: color_data = Z;
		19'b0100000010101001111: color_data = Z;
		19'b0100000010101010000: color_data = Z;
		19'b0100000010101010001: color_data = Z;
		19'b0100000010101010010: color_data = Z;
		19'b0100000010101010011: color_data = Z;
		19'b0100000010101010100: color_data = Z;
		19'b0100000010101010101: color_data = Z;
		19'b0100000010101010110: color_data = Z;
		19'b0100000010101010111: color_data = Z;
		19'b0100000010101011000: color_data = Z;
		19'b0100000010101011001: color_data = Z;
		19'b0100000010101011010: color_data = Z;
		19'b0100000010101011011: color_data = Z;
		19'b0100000010101011100: color_data = Z;
		19'b0100000010101011101: color_data = Z;
		19'b0100000010101011110: color_data = Z;
		19'b0100000010101011111: color_data = Z;
		19'b0100000010101100000: color_data = Z;
		19'b0100000010101100001: color_data = Z;
		19'b0100000010101100010: color_data = Z;
		19'b0100000010101100011: color_data = Z;
		19'b0100000010101100100: color_data = Z;
		19'b0100000010101100101: color_data = Z;
		19'b0100000010101100110: color_data = Z;
		19'b0100000010101100111: color_data = Z;
		19'b0100000010101101000: color_data = Z;
		19'b0100000010101101001: color_data = Z;
		19'b0100000010101101010: color_data = Z;
		19'b0100000010101101011: color_data = Z;
		19'b0100000010101101100: color_data = Z;
		19'b0100000010101101101: color_data = Z;
		19'b0100000010101101110: color_data = Z;
		19'b0100000010101101111: color_data = Z;
		19'b0100000010101110000: color_data = Z;
		19'b0100000010101110001: color_data = Z;
		19'b0100000010101110010: color_data = Z;
		19'b0100000010101110011: color_data = Z;
		19'b0100000010101110100: color_data = Z;
		19'b0100000010101110101: color_data = Z;
		19'b0100000010101110110: color_data = Z;
		19'b0100000010101110111: color_data = Z;
		19'b0100000010101111000: color_data = Z;
		19'b0100000010101111001: color_data = Z;
		19'b0100000010101111010: color_data = Z;
		19'b0100000010101111011: color_data = Z;
		19'b0100000010101111100: color_data = Z;
		19'b0100000010101111101: color_data = Z;
		19'b0100000010101111110: color_data = Z;
		19'b0100000010101111111: color_data = Z;
		19'b0100000010110000000: color_data = Z;
		19'b0100000010110000001: color_data = Z;
		19'b0100000010110000010: color_data = Z;
		19'b0100000010110000011: color_data = Z;
		19'b0100000010110000100: color_data = Z;
		19'b0100000010110000101: color_data = Z;
		19'b0100000010110000110: color_data = Z;
		19'b0100000010110000111: color_data = Z;
		19'b0100000010111001100: color_data = Z;
		19'b0100000010111001101: color_data = Z;
		19'b0100000010111001110: color_data = Z;
		19'b0100000010111001111: color_data = Z;
		19'b0100000010111010000: color_data = Z;
		19'b0100000010111010001: color_data = Z;
		19'b0100000010111010010: color_data = Z;
		19'b0100000010111010011: color_data = Z;
		19'b0100000010111011011: color_data = Z;
		19'b0100000010111011100: color_data = Z;
		19'b0100000010111100000: color_data = Z;
		19'b0100000010111100001: color_data = Z;
		19'b0100000010111100010: color_data = Z;
		19'b0100000100010101011: color_data = Z;
		19'b0100000100010101100: color_data = Z;
		19'b0100000100010110100: color_data = Z;
		19'b0100000100010110101: color_data = Z;
		19'b0100000100010110110: color_data = Z;
		19'b0100000100010110111: color_data = Z;
		19'b0100000100010111000: color_data = Z;
		19'b0100000100010111001: color_data = Z;
		19'b0100000100010111010: color_data = Z;
		19'b0100000100010111011: color_data = Z;
		19'b0100000100011001101: color_data = Z;
		19'b0100000100011001110: color_data = Z;
		19'b0100000100011001111: color_data = Z;
		19'b0100000100011010000: color_data = Z;
		19'b0100000100011010001: color_data = Z;
		19'b0100000100011010010: color_data = Z;
		19'b0100000100011010011: color_data = Z;
		19'b0100000100011010100: color_data = Z;
		19'b0100000100011010101: color_data = Z;
		19'b0100000100011010110: color_data = Z;
		19'b0100000100011010111: color_data = Z;
		19'b0100000100011100001: color_data = Z;
		19'b0100000100011100010: color_data = Z;
		19'b0100000100011100011: color_data = Z;
		19'b0100000100011100110: color_data = Z;
		19'b0100000100011100111: color_data = Z;
		19'b0100000100011101000: color_data = Z;
		19'b0100000100011101001: color_data = Z;
		19'b0100000100011101010: color_data = Z;
		19'b0100000100011101011: color_data = Z;
		19'b0100000100011101100: color_data = Z;
		19'b0100000100011101101: color_data = Z;
		19'b0100000100011101110: color_data = Z;
		19'b0100000100011110001: color_data = Z;
		19'b0100000100011110010: color_data = Z;
		19'b0100000100011110011: color_data = Z;
		19'b0100000100011110100: color_data = Z;
		19'b0100000100011110101: color_data = Z;
		19'b0100000100011111000: color_data = Z;
		19'b0100000100011111001: color_data = Z;
		19'b0100000100011111010: color_data = Z;
		19'b0100000100011111011: color_data = Z;
		19'b0100000100011111100: color_data = Z;
		19'b0100000100011111101: color_data = Z;
		19'b0100000100011111110: color_data = Z;
		19'b0100000100011111111: color_data = Z;
		19'b0100000100100000000: color_data = Z;
		19'b0100000100100000001: color_data = Z;
		19'b0100000100100000010: color_data = Z;
		19'b0100000100100000011: color_data = Z;
		19'b0100000100100000100: color_data = Z;
		19'b0100000100100000101: color_data = Z;
		19'b0100000100100000110: color_data = Z;
		19'b0100000100100000111: color_data = Z;
		19'b0100000100100001000: color_data = Z;
		19'b0100000100100001001: color_data = Z;
		19'b0100000100100001010: color_data = Z;
		19'b0100000100100001011: color_data = Z;
		19'b0100000100100001100: color_data = Z;
		19'b0100000100100001101: color_data = Z;
		19'b0100000100100001110: color_data = Z;
		19'b0100000100100001111: color_data = Z;
		19'b0100000100100010000: color_data = Z;
		19'b0100000100100010001: color_data = Z;
		19'b0100000100100010010: color_data = Z;
		19'b0100000100100010011: color_data = Z;
		19'b0100000100100010100: color_data = Z;
		19'b0100000100100010101: color_data = Z;
		19'b0100000100100010110: color_data = Z;
		19'b0100000100100010111: color_data = Z;
		19'b0100000100100011000: color_data = Z;
		19'b0100000100100011001: color_data = Z;
		19'b0100000100100011010: color_data = Z;
		19'b0100000100100011011: color_data = Z;
		19'b0100000100100011100: color_data = Z;
		19'b0100000100100011101: color_data = Z;
		19'b0100000100100011110: color_data = Z;
		19'b0100000100100011111: color_data = Z;
		19'b0100000100100100000: color_data = Z;
		19'b0100000100100100001: color_data = Z;
		19'b0100000100100100010: color_data = Z;
		19'b0100000100100100011: color_data = Z;
		19'b0100000100100100100: color_data = Z;
		19'b0100000100100100101: color_data = Z;
		19'b0100000100100100110: color_data = Z;
		19'b0100000100100100111: color_data = Z;
		19'b0100000100100101000: color_data = Z;
		19'b0100000100100101001: color_data = Z;
		19'b0100000100100101010: color_data = Z;
		19'b0100000100100101011: color_data = Z;
		19'b0100000100100101100: color_data = Z;
		19'b0100000100100101101: color_data = Z;
		19'b0100000100100101110: color_data = Z;
		19'b0100000100100101111: color_data = Z;
		19'b0100000100100110000: color_data = Z;
		19'b0100000100100110001: color_data = Z;
		19'b0100000100100110010: color_data = Z;
		19'b0100000100100110011: color_data = Z;
		19'b0100000100100110100: color_data = Z;
		19'b0100000100100110101: color_data = Z;
		19'b0100000100100110110: color_data = Z;
		19'b0100000100100110111: color_data = Z;
		19'b0100000100100111000: color_data = Z;
		19'b0100000100100111001: color_data = Z;
		19'b0100000100100111010: color_data = Z;
		19'b0100000100100111011: color_data = Z;
		19'b0100000100100111100: color_data = Z;
		19'b0100000100100111101: color_data = Z;
		19'b0100000100100111110: color_data = Z;
		19'b0100000100100111111: color_data = Z;
		19'b0100000100101000000: color_data = Z;
		19'b0100000100101000001: color_data = Z;
		19'b0100000100101000010: color_data = Z;
		19'b0100000100101000011: color_data = Z;
		19'b0100000100101000100: color_data = Z;
		19'b0100000100101000101: color_data = Z;
		19'b0100000100101000110: color_data = Z;
		19'b0100000100101000111: color_data = Z;
		19'b0100000100101001000: color_data = Z;
		19'b0100000100101001001: color_data = Z;
		19'b0100000100101001010: color_data = Z;
		19'b0100000100101001011: color_data = Z;
		19'b0100000100101001100: color_data = Z;
		19'b0100000100101001101: color_data = Z;
		19'b0100000100101001110: color_data = Z;
		19'b0100000100101001111: color_data = Z;
		19'b0100000100101010000: color_data = Z;
		19'b0100000100101010001: color_data = Z;
		19'b0100000100101010010: color_data = Z;
		19'b0100000100101010011: color_data = Z;
		19'b0100000100101010100: color_data = Z;
		19'b0100000100101010101: color_data = Z;
		19'b0100000100101010110: color_data = Z;
		19'b0100000100101010111: color_data = Z;
		19'b0100000100101011000: color_data = Z;
		19'b0100000100101011001: color_data = Z;
		19'b0100000100101011010: color_data = Z;
		19'b0100000100101011011: color_data = Z;
		19'b0100000100101011100: color_data = Z;
		19'b0100000100101011101: color_data = Z;
		19'b0100000100101011110: color_data = Z;
		19'b0100000100101011111: color_data = Z;
		19'b0100000100101100000: color_data = Z;
		19'b0100000100101100001: color_data = Z;
		19'b0100000100101100010: color_data = Z;
		19'b0100000100101100011: color_data = Z;
		19'b0100000100101100100: color_data = Z;
		19'b0100000100101100101: color_data = Z;
		19'b0100000100101100110: color_data = Z;
		19'b0100000100101100111: color_data = Z;
		19'b0100000100101101000: color_data = Z;
		19'b0100000100101101001: color_data = Z;
		19'b0100000100101101010: color_data = Z;
		19'b0100000100101101011: color_data = Z;
		19'b0100000100101101100: color_data = Z;
		19'b0100000100101101101: color_data = Z;
		19'b0100000100101101110: color_data = Z;
		19'b0100000100101101111: color_data = Z;
		19'b0100000100101110000: color_data = Z;
		19'b0100000100101110001: color_data = Z;
		19'b0100000100101110010: color_data = Z;
		19'b0100000100101110011: color_data = Z;
		19'b0100000100101110100: color_data = Z;
		19'b0100000100101110101: color_data = Z;
		19'b0100000100101110110: color_data = Z;
		19'b0100000100101110111: color_data = Z;
		19'b0100000100101111000: color_data = Z;
		19'b0100000100101111001: color_data = Z;
		19'b0100000100101111010: color_data = Z;
		19'b0100000100101111011: color_data = Z;
		19'b0100000100101111100: color_data = Z;
		19'b0100000100101111101: color_data = Z;
		19'b0100000100101111110: color_data = Z;
		19'b0100000100101111111: color_data = Z;
		19'b0100000100110000000: color_data = Z;
		19'b0100000100110000001: color_data = Z;
		19'b0100000100110000010: color_data = Z;
		19'b0100000100110000011: color_data = Z;
		19'b0100000100110000100: color_data = Z;
		19'b0100000100110000101: color_data = Z;
		19'b0100000100110000110: color_data = Z;
		19'b0100000100111001011: color_data = Z;
		19'b0100000100111001100: color_data = Z;
		19'b0100000100111001101: color_data = Z;
		19'b0100000100111001110: color_data = Z;
		19'b0100000100111001111: color_data = Z;
		19'b0100000100111010000: color_data = Z;
		19'b0100000100111010001: color_data = Z;
		19'b0100000100111010011: color_data = Z;
		19'b0100000100111010100: color_data = Z;
		19'b0100000100111011011: color_data = Z;
		19'b0100000100111100000: color_data = Z;
		19'b0100000100111100001: color_data = Z;
		19'b0100000100111100010: color_data = Z;
		19'b0100000110010101011: color_data = Z;
		19'b0100000110010110100: color_data = Z;
		19'b0100000110010110101: color_data = Z;
		19'b0100000110010110110: color_data = Z;
		19'b0100000110010110111: color_data = Z;
		19'b0100000110010111000: color_data = Z;
		19'b0100000110010111001: color_data = Z;
		19'b0100000110010111010: color_data = Z;
		19'b0100000110011001011: color_data = Z;
		19'b0100000110011001100: color_data = Z;
		19'b0100000110011001101: color_data = Z;
		19'b0100000110011001110: color_data = Z;
		19'b0100000110011010010: color_data = Z;
		19'b0100000110011010011: color_data = Z;
		19'b0100000110011010100: color_data = Z;
		19'b0100000110011010101: color_data = Z;
		19'b0100000110011010110: color_data = Z;
		19'b0100000110011011101: color_data = Z;
		19'b0100000110011011110: color_data = Z;
		19'b0100000110011011111: color_data = Z;
		19'b0100000110011100000: color_data = Z;
		19'b0100000110011100001: color_data = Z;
		19'b0100000110011100010: color_data = Z;
		19'b0100000110011100011: color_data = Z;
		19'b0100000110011100100: color_data = Z;
		19'b0100000110011100101: color_data = Z;
		19'b0100000110011111010: color_data = Z;
		19'b0100000110011111011: color_data = Z;
		19'b0100000110011111100: color_data = Z;
		19'b0100000110011111101: color_data = Z;
		19'b0100000110011111110: color_data = Z;
		19'b0100000110011111111: color_data = Z;
		19'b0100000110100000000: color_data = Z;
		19'b0100000110100000001: color_data = Z;
		19'b0100000110100000010: color_data = Z;
		19'b0100000110100000011: color_data = Z;
		19'b0100000110100000100: color_data = Z;
		19'b0100000110100000101: color_data = Z;
		19'b0100000110100000110: color_data = Z;
		19'b0100000110100000111: color_data = Z;
		19'b0100000110100001000: color_data = Z;
		19'b0100000110100001001: color_data = Z;
		19'b0100000110100001010: color_data = Z;
		19'b0100000110100001011: color_data = Z;
		19'b0100000110100001100: color_data = Z;
		19'b0100000110100001101: color_data = Z;
		19'b0100000110100001110: color_data = Z;
		19'b0100000110100001111: color_data = Z;
		19'b0100000110100010000: color_data = Z;
		19'b0100000110100010001: color_data = Z;
		19'b0100000110100010010: color_data = Z;
		19'b0100000110100010011: color_data = Z;
		19'b0100000110100010100: color_data = Z;
		19'b0100000110100010101: color_data = Z;
		19'b0100000110100010110: color_data = Z;
		19'b0100000110100010111: color_data = Z;
		19'b0100000110100011000: color_data = Z;
		19'b0100000110100011001: color_data = Z;
		19'b0100000110100011010: color_data = Z;
		19'b0100000110100011011: color_data = Z;
		19'b0100000110100011100: color_data = Z;
		19'b0100000110100011101: color_data = Z;
		19'b0100000110100011110: color_data = Z;
		19'b0100000110100011111: color_data = Z;
		19'b0100000110100100000: color_data = Z;
		19'b0100000110100100001: color_data = Z;
		19'b0100000110100100010: color_data = Z;
		19'b0100000110100100011: color_data = Z;
		19'b0100000110100100100: color_data = Z;
		19'b0100000110100100101: color_data = Z;
		19'b0100000110100100110: color_data = Z;
		19'b0100000110100100111: color_data = Z;
		19'b0100000110100101000: color_data = Z;
		19'b0100000110100101001: color_data = Z;
		19'b0100000110100101010: color_data = Z;
		19'b0100000110100101011: color_data = Z;
		19'b0100000110100101100: color_data = Z;
		19'b0100000110100101101: color_data = Z;
		19'b0100000110100101110: color_data = Z;
		19'b0100000110100101111: color_data = Z;
		19'b0100000110100110000: color_data = Z;
		19'b0100000110100110001: color_data = Z;
		19'b0100000110100110010: color_data = Z;
		19'b0100000110100110011: color_data = Z;
		19'b0100000110100110100: color_data = Z;
		19'b0100000110100110101: color_data = Z;
		19'b0100000110100110110: color_data = Z;
		19'b0100000110100110111: color_data = Z;
		19'b0100000110100111000: color_data = Z;
		19'b0100000110100111001: color_data = Z;
		19'b0100000110100111010: color_data = Z;
		19'b0100000110100111011: color_data = Z;
		19'b0100000110100111100: color_data = Z;
		19'b0100000110100111101: color_data = Z;
		19'b0100000110100111110: color_data = Z;
		19'b0100000110100111111: color_data = Z;
		19'b0100000110101000000: color_data = Z;
		19'b0100000110101000001: color_data = Z;
		19'b0100000110101000010: color_data = Z;
		19'b0100000110101000011: color_data = Z;
		19'b0100000110101000100: color_data = Z;
		19'b0100000110101000101: color_data = Z;
		19'b0100000110101000110: color_data = Z;
		19'b0100000110101000111: color_data = Z;
		19'b0100000110101001000: color_data = Z;
		19'b0100000110101001001: color_data = Z;
		19'b0100000110101001010: color_data = Z;
		19'b0100000110101001011: color_data = Z;
		19'b0100000110101001100: color_data = Z;
		19'b0100000110101001101: color_data = Z;
		19'b0100000110101001110: color_data = Z;
		19'b0100000110101001111: color_data = Z;
		19'b0100000110101010000: color_data = Z;
		19'b0100000110101010001: color_data = Z;
		19'b0100000110101010010: color_data = Z;
		19'b0100000110101010011: color_data = Z;
		19'b0100000110101010100: color_data = Z;
		19'b0100000110101010101: color_data = Z;
		19'b0100000110101010110: color_data = Z;
		19'b0100000110101010111: color_data = Z;
		19'b0100000110101011000: color_data = Z;
		19'b0100000110101011001: color_data = Z;
		19'b0100000110101011010: color_data = Z;
		19'b0100000110101011011: color_data = Z;
		19'b0100000110101011100: color_data = Z;
		19'b0100000110101011101: color_data = Z;
		19'b0100000110101011110: color_data = Z;
		19'b0100000110101011111: color_data = Z;
		19'b0100000110101100000: color_data = Z;
		19'b0100000110101100001: color_data = Z;
		19'b0100000110101100010: color_data = Z;
		19'b0100000110101100011: color_data = Z;
		19'b0100000110101100100: color_data = Z;
		19'b0100000110101100101: color_data = Z;
		19'b0100000110101100110: color_data = Z;
		19'b0100000110101100111: color_data = Z;
		19'b0100000110101101000: color_data = Z;
		19'b0100000110101101001: color_data = Z;
		19'b0100000110101101010: color_data = Z;
		19'b0100000110101101011: color_data = Z;
		19'b0100000110101101100: color_data = Z;
		19'b0100000110101101101: color_data = Z;
		19'b0100000110101101110: color_data = Z;
		19'b0100000110101101111: color_data = Z;
		19'b0100000110101110000: color_data = Z;
		19'b0100000110101110001: color_data = Z;
		19'b0100000110101110010: color_data = Z;
		19'b0100000110101110011: color_data = Z;
		19'b0100000110101110100: color_data = Z;
		19'b0100000110101110101: color_data = Z;
		19'b0100000110101110110: color_data = Z;
		19'b0100000110101110111: color_data = Z;
		19'b0100000110101111000: color_data = Z;
		19'b0100000110101111001: color_data = Z;
		19'b0100000110101111010: color_data = Z;
		19'b0100000110101111011: color_data = Z;
		19'b0100000110101111100: color_data = Z;
		19'b0100000110101111101: color_data = Z;
		19'b0100000110101111110: color_data = Z;
		19'b0100000110101111111: color_data = Z;
		19'b0100000110110000000: color_data = Z;
		19'b0100000110110000001: color_data = Z;
		19'b0100000110110000010: color_data = Z;
		19'b0100000110110000011: color_data = Z;
		19'b0100000110110000100: color_data = Z;
		19'b0100000110110000101: color_data = Z;
		19'b0100000110110000110: color_data = Z;
		19'b0100000110111001011: color_data = Z;
		19'b0100000110111001100: color_data = Z;
		19'b0100000110111001101: color_data = Z;
		19'b0100000110111001110: color_data = Z;
		19'b0100000110111001111: color_data = Z;
		19'b0100000110111010000: color_data = Z;
		19'b0100000110111010001: color_data = Z;
		19'b0100000110111010011: color_data = Z;
		19'b0100000110111010100: color_data = Z;
		19'b0100000110111100001: color_data = Z;
		19'b0100000110111100010: color_data = Z;
		19'b0100001000010101010: color_data = Z;
		19'b0100001000010101011: color_data = Z;
		19'b0100001000010110101: color_data = Z;
		19'b0100001000010110110: color_data = Z;
		19'b0100001000010110111: color_data = Z;
		19'b0100001000010111000: color_data = Z;
		19'b0100001000010111001: color_data = Z;
		19'b0100001000011001001: color_data = Z;
		19'b0100001000011001010: color_data = Z;
		19'b0100001000011001011: color_data = Z;
		19'b0100001000011001100: color_data = Z;
		19'b0100001000011010000: color_data = Z;
		19'b0100001000011010001: color_data = Z;
		19'b0100001000011010010: color_data = Z;
		19'b0100001000011010011: color_data = Z;
		19'b0100001000011010100: color_data = Z;
		19'b0100001000011010101: color_data = Z;
		19'b0100001000011010110: color_data = Z;
		19'b0100001000011010111: color_data = Z;
		19'b0100001000011011000: color_data = Z;
		19'b0100001000011011001: color_data = Z;
		19'b0100001000011011010: color_data = Z;
		19'b0100001000011011011: color_data = Z;
		19'b0100001000011011100: color_data = Z;
		19'b0100001000011011101: color_data = Z;
		19'b0100001000011011110: color_data = Z;
		19'b0100001000011011111: color_data = Z;
		19'b0100001000011100000: color_data = Z;
		19'b0100001000011100001: color_data = Z;
		19'b0100001000011100010: color_data = Z;
		19'b0100001000011100011: color_data = Z;
		19'b0100001000011100100: color_data = Z;
		19'b0100001000011111010: color_data = Z;
		19'b0100001000011111011: color_data = Z;
		19'b0100001000011111100: color_data = Z;
		19'b0100001000011111101: color_data = Z;
		19'b0100001000011111110: color_data = Z;
		19'b0100001000011111111: color_data = Z;
		19'b0100001000100000000: color_data = Z;
		19'b0100001000100000001: color_data = Z;
		19'b0100001000100000010: color_data = Z;
		19'b0100001000100000011: color_data = Z;
		19'b0100001000100000100: color_data = Z;
		19'b0100001000100000101: color_data = Z;
		19'b0100001000100000110: color_data = Z;
		19'b0100001000100000111: color_data = Z;
		19'b0100001000100001000: color_data = Z;
		19'b0100001000100001001: color_data = Z;
		19'b0100001000100001010: color_data = Z;
		19'b0100001000100001011: color_data = Z;
		19'b0100001000100001100: color_data = Z;
		19'b0100001000100001101: color_data = Z;
		19'b0100001000100001110: color_data = Z;
		19'b0100001000100001111: color_data = Z;
		19'b0100001000100010000: color_data = Z;
		19'b0100001000100010001: color_data = Z;
		19'b0100001000100010010: color_data = Z;
		19'b0100001000100010011: color_data = Z;
		19'b0100001000100010100: color_data = Z;
		19'b0100001000100010101: color_data = Z;
		19'b0100001000100010110: color_data = Z;
		19'b0100001000100010111: color_data = Z;
		19'b0100001000100011000: color_data = Z;
		19'b0100001000100011001: color_data = Z;
		19'b0100001000100011010: color_data = Z;
		19'b0100001000100011011: color_data = Z;
		19'b0100001000100011100: color_data = Z;
		19'b0100001000100011101: color_data = Z;
		19'b0100001000100011110: color_data = Z;
		19'b0100001000100011111: color_data = Z;
		19'b0100001000100100000: color_data = Z;
		19'b0100001000100100001: color_data = Z;
		19'b0100001000100100010: color_data = Z;
		19'b0100001000100100011: color_data = Z;
		19'b0100001000100100100: color_data = Z;
		19'b0100001000100100101: color_data = Z;
		19'b0100001000100100110: color_data = Z;
		19'b0100001000100100111: color_data = Z;
		19'b0100001000100101000: color_data = Z;
		19'b0100001000100101001: color_data = Z;
		19'b0100001000100101010: color_data = Z;
		19'b0100001000100101011: color_data = Z;
		19'b0100001000100101100: color_data = Z;
		19'b0100001000100101101: color_data = Z;
		19'b0100001000100101110: color_data = Z;
		19'b0100001000100101111: color_data = Z;
		19'b0100001000100110000: color_data = Z;
		19'b0100001000100110001: color_data = Z;
		19'b0100001000100110010: color_data = Z;
		19'b0100001000100110011: color_data = Z;
		19'b0100001000100110100: color_data = Z;
		19'b0100001000100110101: color_data = Z;
		19'b0100001000100110110: color_data = Z;
		19'b0100001000100110111: color_data = Z;
		19'b0100001000100111000: color_data = Z;
		19'b0100001000100111001: color_data = Z;
		19'b0100001000100111010: color_data = Z;
		19'b0100001000100111011: color_data = Z;
		19'b0100001000100111100: color_data = Z;
		19'b0100001000100111101: color_data = Z;
		19'b0100001000100111110: color_data = Z;
		19'b0100001000100111111: color_data = Z;
		19'b0100001000101000000: color_data = Z;
		19'b0100001000101000001: color_data = Z;
		19'b0100001000101000010: color_data = Z;
		19'b0100001000101000011: color_data = Z;
		19'b0100001000101000100: color_data = Z;
		19'b0100001000101000101: color_data = Z;
		19'b0100001000101000110: color_data = Z;
		19'b0100001000101000111: color_data = Z;
		19'b0100001000101001000: color_data = Z;
		19'b0100001000101001001: color_data = Z;
		19'b0100001000101001010: color_data = Z;
		19'b0100001000101001011: color_data = Z;
		19'b0100001000101001100: color_data = Z;
		19'b0100001000101001101: color_data = Z;
		19'b0100001000101001110: color_data = Z;
		19'b0100001000101001111: color_data = Z;
		19'b0100001000101010000: color_data = Z;
		19'b0100001000101010001: color_data = Z;
		19'b0100001000101010010: color_data = Z;
		19'b0100001000101010011: color_data = Z;
		19'b0100001000101010100: color_data = Z;
		19'b0100001000101010101: color_data = Z;
		19'b0100001000101010110: color_data = Z;
		19'b0100001000101010111: color_data = Z;
		19'b0100001000101011000: color_data = Z;
		19'b0100001000101011001: color_data = Z;
		19'b0100001000101011010: color_data = Z;
		19'b0100001000101011011: color_data = Z;
		19'b0100001000101011100: color_data = Z;
		19'b0100001000101011101: color_data = Z;
		19'b0100001000101011110: color_data = Z;
		19'b0100001000101011111: color_data = Z;
		19'b0100001000101100000: color_data = Z;
		19'b0100001000101100001: color_data = Z;
		19'b0100001000101100010: color_data = Z;
		19'b0100001000101100011: color_data = Z;
		19'b0100001000101100100: color_data = Z;
		19'b0100001000101100101: color_data = Z;
		19'b0100001000101100110: color_data = Z;
		19'b0100001000101100111: color_data = Z;
		19'b0100001000101101000: color_data = Z;
		19'b0100001000101101001: color_data = Z;
		19'b0100001000101101010: color_data = Z;
		19'b0100001000101101011: color_data = Z;
		19'b0100001000101101100: color_data = Z;
		19'b0100001000101101101: color_data = Z;
		19'b0100001000101101110: color_data = Z;
		19'b0100001000101101111: color_data = Z;
		19'b0100001000101110000: color_data = Z;
		19'b0100001000101110001: color_data = Z;
		19'b0100001000101110010: color_data = Z;
		19'b0100001000101110011: color_data = Z;
		19'b0100001000101110100: color_data = Z;
		19'b0100001000101110101: color_data = Z;
		19'b0100001000101110110: color_data = Z;
		19'b0100001000101110111: color_data = Z;
		19'b0100001000101111000: color_data = Z;
		19'b0100001000101111001: color_data = Z;
		19'b0100001000101111010: color_data = Z;
		19'b0100001000101111011: color_data = Z;
		19'b0100001000101111100: color_data = Z;
		19'b0100001000101111101: color_data = Z;
		19'b0100001000101111110: color_data = Z;
		19'b0100001000101111111: color_data = Z;
		19'b0100001000110000000: color_data = Z;
		19'b0100001000110000001: color_data = Z;
		19'b0100001000110000010: color_data = Z;
		19'b0100001000110000011: color_data = Z;
		19'b0100001000110000100: color_data = Z;
		19'b0100001000110000101: color_data = Z;
		19'b0100001000110000110: color_data = Z;
		19'b0100001000111001100: color_data = Z;
		19'b0100001000111001101: color_data = Z;
		19'b0100001000111001110: color_data = Z;
		19'b0100001000111001111: color_data = Z;
		19'b0100001000111010000: color_data = Z;
		19'b0100001000111010001: color_data = Z;
		19'b0100001000111010011: color_data = Z;
		19'b0100001000111010100: color_data = Z;
		19'b0100001000111010101: color_data = Z;
		19'b0100001000111100001: color_data = Z;
		19'b0100001000111100010: color_data = Z;
		19'b0100001010010101001: color_data = Z;
		19'b0100001010010101010: color_data = Z;
		19'b0100001010010110101: color_data = Z;
		19'b0100001010010110110: color_data = Z;
		19'b0100001010010110111: color_data = Z;
		19'b0100001010010111000: color_data = Z;
		19'b0100001010011001000: color_data = Z;
		19'b0100001010011001001: color_data = Z;
		19'b0100001010011001010: color_data = Z;
		19'b0100001010011001111: color_data = Z;
		19'b0100001010011010000: color_data = Z;
		19'b0100001010011010001: color_data = Z;
		19'b0100001010011010010: color_data = Z;
		19'b0100001010011010011: color_data = Z;
		19'b0100001010011010100: color_data = Z;
		19'b0100001010011010101: color_data = Z;
		19'b0100001010011010110: color_data = Z;
		19'b0100001010011010111: color_data = Z;
		19'b0100001010011011000: color_data = Z;
		19'b0100001010011011001: color_data = Z;
		19'b0100001010011011010: color_data = Z;
		19'b0100001010011011011: color_data = Z;
		19'b0100001010011100000: color_data = Z;
		19'b0100001010011100001: color_data = Z;
		19'b0100001010011111010: color_data = Z;
		19'b0100001010011111011: color_data = Z;
		19'b0100001010011111100: color_data = Z;
		19'b0100001010011111101: color_data = Z;
		19'b0100001010011111110: color_data = Z;
		19'b0100001010011111111: color_data = Z;
		19'b0100001010100000000: color_data = Z;
		19'b0100001010100000001: color_data = Z;
		19'b0100001010100000010: color_data = Z;
		19'b0100001010100000011: color_data = Z;
		19'b0100001010100000100: color_data = Z;
		19'b0100001010100000101: color_data = Z;
		19'b0100001010100000110: color_data = Z;
		19'b0100001010100000111: color_data = Z;
		19'b0100001010100001000: color_data = Z;
		19'b0100001010100001001: color_data = Z;
		19'b0100001010100001010: color_data = Z;
		19'b0100001010100001011: color_data = Z;
		19'b0100001010100001100: color_data = Z;
		19'b0100001010100001101: color_data = Z;
		19'b0100001010100001110: color_data = Z;
		19'b0100001010100001111: color_data = Z;
		19'b0100001010100010000: color_data = Z;
		19'b0100001010100010001: color_data = Z;
		19'b0100001010100010010: color_data = Z;
		19'b0100001010100010011: color_data = Z;
		19'b0100001010100010100: color_data = Z;
		19'b0100001010100010101: color_data = Z;
		19'b0100001010100010110: color_data = Z;
		19'b0100001010100010111: color_data = Z;
		19'b0100001010100011000: color_data = Z;
		19'b0100001010100011001: color_data = Z;
		19'b0100001010100011010: color_data = Z;
		19'b0100001010100011011: color_data = Z;
		19'b0100001010100011100: color_data = Z;
		19'b0100001010100011101: color_data = Z;
		19'b0100001010100011110: color_data = Z;
		19'b0100001010100011111: color_data = Z;
		19'b0100001010100100000: color_data = Z;
		19'b0100001010100100001: color_data = Z;
		19'b0100001010100100010: color_data = Z;
		19'b0100001010100100011: color_data = Z;
		19'b0100001010100100100: color_data = Z;
		19'b0100001010100100101: color_data = Z;
		19'b0100001010100100110: color_data = Z;
		19'b0100001010100100111: color_data = Z;
		19'b0100001010100101000: color_data = Z;
		19'b0100001010100101001: color_data = Z;
		19'b0100001010100101010: color_data = Z;
		19'b0100001010100101011: color_data = Z;
		19'b0100001010100101100: color_data = Z;
		19'b0100001010100101101: color_data = Z;
		19'b0100001010100101110: color_data = Z;
		19'b0100001010100101111: color_data = Z;
		19'b0100001010100110000: color_data = Z;
		19'b0100001010100110001: color_data = Z;
		19'b0100001010100110010: color_data = Z;
		19'b0100001010100110011: color_data = Z;
		19'b0100001010100110100: color_data = Z;
		19'b0100001010100110101: color_data = Z;
		19'b0100001010100110110: color_data = Z;
		19'b0100001010100110111: color_data = Z;
		19'b0100001010100111000: color_data = Z;
		19'b0100001010100111001: color_data = Z;
		19'b0100001010100111010: color_data = Z;
		19'b0100001010100111011: color_data = Z;
		19'b0100001010100111100: color_data = Z;
		19'b0100001010100111101: color_data = Z;
		19'b0100001010100111110: color_data = Z;
		19'b0100001010100111111: color_data = Z;
		19'b0100001010101000000: color_data = Z;
		19'b0100001010101000001: color_data = Z;
		19'b0100001010101000010: color_data = Z;
		19'b0100001010101000011: color_data = Z;
		19'b0100001010101000100: color_data = Z;
		19'b0100001010101000101: color_data = Z;
		19'b0100001010101000110: color_data = Z;
		19'b0100001010101000111: color_data = Z;
		19'b0100001010101001000: color_data = Z;
		19'b0100001010101001001: color_data = Z;
		19'b0100001010101001010: color_data = Z;
		19'b0100001010101001011: color_data = Z;
		19'b0100001010101001100: color_data = Z;
		19'b0100001010101001101: color_data = Z;
		19'b0100001010101001110: color_data = Z;
		19'b0100001010101001111: color_data = Z;
		19'b0100001010101010000: color_data = Z;
		19'b0100001010101010001: color_data = Z;
		19'b0100001010101010010: color_data = Z;
		19'b0100001010101010011: color_data = Z;
		19'b0100001010101010100: color_data = Z;
		19'b0100001010101010101: color_data = Z;
		19'b0100001010101010110: color_data = Z;
		19'b0100001010101010111: color_data = Z;
		19'b0100001010101011000: color_data = Z;
		19'b0100001010101011001: color_data = Z;
		19'b0100001010101011010: color_data = Z;
		19'b0100001010101011011: color_data = Z;
		19'b0100001010101011100: color_data = Z;
		19'b0100001010101011101: color_data = Z;
		19'b0100001010101011110: color_data = Z;
		19'b0100001010101011111: color_data = Z;
		19'b0100001010101100000: color_data = Z;
		19'b0100001010101100001: color_data = Z;
		19'b0100001010101100010: color_data = Z;
		19'b0100001010101100011: color_data = Z;
		19'b0100001010101100100: color_data = Z;
		19'b0100001010101100101: color_data = Z;
		19'b0100001010101100110: color_data = Z;
		19'b0100001010101100111: color_data = Z;
		19'b0100001010101101000: color_data = Z;
		19'b0100001010101101001: color_data = Z;
		19'b0100001010101101010: color_data = Z;
		19'b0100001010101101011: color_data = Z;
		19'b0100001010101101100: color_data = Z;
		19'b0100001010101101101: color_data = Z;
		19'b0100001010101101110: color_data = Z;
		19'b0100001010101101111: color_data = Z;
		19'b0100001010101110000: color_data = Z;
		19'b0100001010101110001: color_data = Z;
		19'b0100001010101110010: color_data = Z;
		19'b0100001010101110011: color_data = Z;
		19'b0100001010101110100: color_data = Z;
		19'b0100001010101110101: color_data = Z;
		19'b0100001010101110110: color_data = Z;
		19'b0100001010101110111: color_data = Z;
		19'b0100001010101111000: color_data = Z;
		19'b0100001010101111001: color_data = Z;
		19'b0100001010101111010: color_data = Z;
		19'b0100001010101111011: color_data = Z;
		19'b0100001010101111100: color_data = Z;
		19'b0100001010101111101: color_data = Z;
		19'b0100001010101111110: color_data = Z;
		19'b0100001010101111111: color_data = Z;
		19'b0100001010110000010: color_data = Z;
		19'b0100001010110000011: color_data = Z;
		19'b0100001010110000100: color_data = Z;
		19'b0100001010110000101: color_data = Z;
		19'b0100001010111001100: color_data = Z;
		19'b0100001010111001101: color_data = Z;
		19'b0100001010111001110: color_data = Z;
		19'b0100001010111001111: color_data = Z;
		19'b0100001010111010000: color_data = Z;
		19'b0100001010111010001: color_data = Z;
		19'b0100001010111010010: color_data = Z;
		19'b0100001010111010011: color_data = Z;
		19'b0100001010111010100: color_data = Z;
		19'b0100001010111010101: color_data = Z;
		19'b0100001010111100001: color_data = Z;
		19'b0100001010111100010: color_data = Z;
		19'b0100001010111100011: color_data = Z;
		19'b0100001100010110100: color_data = Z;
		19'b0100001100010110101: color_data = Z;
		19'b0100001100010110110: color_data = Z;
		19'b0100001100011001000: color_data = Z;
		19'b0100001100011001001: color_data = Z;
		19'b0100001100011001101: color_data = Z;
		19'b0100001100011001110: color_data = Z;
		19'b0100001100011001111: color_data = Z;
		19'b0100001100011010000: color_data = Z;
		19'b0100001100011010001: color_data = Z;
		19'b0100001100011010010: color_data = Z;
		19'b0100001100011010011: color_data = Z;
		19'b0100001100011010100: color_data = Z;
		19'b0100001100011010101: color_data = Z;
		19'b0100001100011010110: color_data = Z;
		19'b0100001100011111011: color_data = Z;
		19'b0100001100011111100: color_data = Z;
		19'b0100001100011111101: color_data = Z;
		19'b0100001100011111110: color_data = Z;
		19'b0100001100011111111: color_data = Z;
		19'b0100001100100000000: color_data = Z;
		19'b0100001100100000001: color_data = Z;
		19'b0100001100100000010: color_data = Z;
		19'b0100001100100000011: color_data = Z;
		19'b0100001100100000100: color_data = Z;
		19'b0100001100100000101: color_data = Z;
		19'b0100001100100000110: color_data = Z;
		19'b0100001100100000111: color_data = Z;
		19'b0100001100100001000: color_data = Z;
		19'b0100001100100001001: color_data = Z;
		19'b0100001100100001010: color_data = Z;
		19'b0100001100100001011: color_data = Z;
		19'b0100001100100001100: color_data = Z;
		19'b0100001100100001101: color_data = Z;
		19'b0100001100100001110: color_data = Z;
		19'b0100001100100001111: color_data = Z;
		19'b0100001100100010000: color_data = Z;
		19'b0100001100100010001: color_data = Z;
		19'b0100001100100010010: color_data = Z;
		19'b0100001100100010011: color_data = Z;
		19'b0100001100100010100: color_data = Z;
		19'b0100001100100010101: color_data = Z;
		19'b0100001100100010110: color_data = Z;
		19'b0100001100100010111: color_data = Z;
		19'b0100001100100011000: color_data = Z;
		19'b0100001100100011001: color_data = Z;
		19'b0100001100100011010: color_data = Z;
		19'b0100001100100011011: color_data = Z;
		19'b0100001100100011100: color_data = Z;
		19'b0100001100100011101: color_data = Z;
		19'b0100001100100011110: color_data = Z;
		19'b0100001100100011111: color_data = Z;
		19'b0100001100100100000: color_data = Z;
		19'b0100001100100100001: color_data = Z;
		19'b0100001100100100010: color_data = Z;
		19'b0100001100100100011: color_data = Z;
		19'b0100001100100100100: color_data = Z;
		19'b0100001100100100101: color_data = Z;
		19'b0100001100100100110: color_data = Z;
		19'b0100001100100100111: color_data = Z;
		19'b0100001100100101000: color_data = Z;
		19'b0100001100100101001: color_data = Z;
		19'b0100001100100101010: color_data = Z;
		19'b0100001100100101011: color_data = Z;
		19'b0100001100100101100: color_data = Z;
		19'b0100001100100101101: color_data = Z;
		19'b0100001100100101110: color_data = Z;
		19'b0100001100100101111: color_data = Z;
		19'b0100001100100110000: color_data = Z;
		19'b0100001100100110001: color_data = Z;
		19'b0100001100100110010: color_data = Z;
		19'b0100001100100110011: color_data = Z;
		19'b0100001100100110100: color_data = Z;
		19'b0100001100100110101: color_data = Z;
		19'b0100001100100110110: color_data = Z;
		19'b0100001100100110111: color_data = Z;
		19'b0100001100100111000: color_data = Z;
		19'b0100001100100111001: color_data = Z;
		19'b0100001100100111010: color_data = Z;
		19'b0100001100100111011: color_data = Z;
		19'b0100001100100111100: color_data = Z;
		19'b0100001100100111101: color_data = Z;
		19'b0100001100100111110: color_data = Z;
		19'b0100001100100111111: color_data = Z;
		19'b0100001100101000000: color_data = Z;
		19'b0100001100101000001: color_data = Z;
		19'b0100001100101000010: color_data = Z;
		19'b0100001100101000011: color_data = Z;
		19'b0100001100101000100: color_data = Z;
		19'b0100001100101000101: color_data = Z;
		19'b0100001100101000110: color_data = Z;
		19'b0100001100101000111: color_data = Z;
		19'b0100001100101001000: color_data = Z;
		19'b0100001100101001001: color_data = Z;
		19'b0100001100101001010: color_data = Z;
		19'b0100001100101001011: color_data = Z;
		19'b0100001100101001100: color_data = Z;
		19'b0100001100101001101: color_data = Z;
		19'b0100001100101001110: color_data = Z;
		19'b0100001100101001111: color_data = Z;
		19'b0100001100101010000: color_data = Z;
		19'b0100001100101010001: color_data = Z;
		19'b0100001100101010010: color_data = Z;
		19'b0100001100101010011: color_data = Z;
		19'b0100001100101010100: color_data = Z;
		19'b0100001100101010101: color_data = Z;
		19'b0100001100101010110: color_data = Z;
		19'b0100001100101010111: color_data = Z;
		19'b0100001100101011000: color_data = Z;
		19'b0100001100101011001: color_data = Z;
		19'b0100001100101011010: color_data = Z;
		19'b0100001100101011011: color_data = Z;
		19'b0100001100101011100: color_data = Z;
		19'b0100001100101011101: color_data = Z;
		19'b0100001100101011110: color_data = Z;
		19'b0100001100101011111: color_data = Z;
		19'b0100001100101100000: color_data = Z;
		19'b0100001100101100001: color_data = Z;
		19'b0100001100101100010: color_data = Z;
		19'b0100001100101100011: color_data = Z;
		19'b0100001100101100100: color_data = Z;
		19'b0100001100101100101: color_data = Z;
		19'b0100001100101100110: color_data = Z;
		19'b0100001100101100111: color_data = Z;
		19'b0100001100101101000: color_data = Z;
		19'b0100001100101101001: color_data = Z;
		19'b0100001100101101010: color_data = Z;
		19'b0100001100101101011: color_data = Z;
		19'b0100001100101101100: color_data = Z;
		19'b0100001100101101101: color_data = Z;
		19'b0100001100101101110: color_data = Z;
		19'b0100001100101101111: color_data = Z;
		19'b0100001100101110000: color_data = Z;
		19'b0100001100101110001: color_data = Z;
		19'b0100001100101110010: color_data = Z;
		19'b0100001100101110011: color_data = Z;
		19'b0100001100101110100: color_data = Z;
		19'b0100001100101110101: color_data = Z;
		19'b0100001100101110110: color_data = Z;
		19'b0100001100101110111: color_data = Z;
		19'b0100001100101111000: color_data = Z;
		19'b0100001100101111001: color_data = Z;
		19'b0100001100101111010: color_data = Z;
		19'b0100001100101111011: color_data = Z;
		19'b0100001100101111100: color_data = Z;
		19'b0100001100101111101: color_data = Z;
		19'b0100001100101111110: color_data = Z;
		19'b0100001100101111111: color_data = Z;
		19'b0100001100110000001: color_data = Z;
		19'b0100001100110000010: color_data = Z;
		19'b0100001100110000011: color_data = Z;
		19'b0100001100110000100: color_data = Z;
		19'b0100001100111001101: color_data = Z;
		19'b0100001100111001110: color_data = Z;
		19'b0100001100111001111: color_data = Z;
		19'b0100001100111010000: color_data = Z;
		19'b0100001100111010001: color_data = Z;
		19'b0100001100111010010: color_data = Z;
		19'b0100001100111010011: color_data = Z;
		19'b0100001100111010100: color_data = Z;
		19'b0100001100111010101: color_data = Z;
		19'b0100001100111010110: color_data = Z;
		19'b0100001100111100011: color_data = Z;
		19'b0100001110010110100: color_data = Z;
		19'b0100001110010110101: color_data = Z;
		19'b0100001110010110110: color_data = Z;
		19'b0100001110011001100: color_data = Z;
		19'b0100001110011001101: color_data = Z;
		19'b0100001110011001110: color_data = Z;
		19'b0100001110011001111: color_data = Z;
		19'b0100001110011010000: color_data = Z;
		19'b0100001110011010001: color_data = Z;
		19'b0100001110011010010: color_data = Z;
		19'b0100001110011010011: color_data = Z;
		19'b0100001110011111011: color_data = Z;
		19'b0100001110011111100: color_data = Z;
		19'b0100001110011111101: color_data = Z;
		19'b0100001110011111110: color_data = Z;
		19'b0100001110011111111: color_data = Z;
		19'b0100001110100000000: color_data = Z;
		19'b0100001110100000001: color_data = Z;
		19'b0100001110100000010: color_data = Z;
		19'b0100001110100000011: color_data = Z;
		19'b0100001110100000100: color_data = Z;
		19'b0100001110100000101: color_data = Z;
		19'b0100001110100000110: color_data = Z;
		19'b0100001110100000111: color_data = Z;
		19'b0100001110100001000: color_data = Z;
		19'b0100001110100001001: color_data = Z;
		19'b0100001110100001010: color_data = Z;
		19'b0100001110100001011: color_data = Z;
		19'b0100001110100001100: color_data = Z;
		19'b0100001110100001101: color_data = Z;
		19'b0100001110100001110: color_data = Z;
		19'b0100001110100001111: color_data = Z;
		19'b0100001110100010000: color_data = Z;
		19'b0100001110100010001: color_data = Z;
		19'b0100001110100010010: color_data = Z;
		19'b0100001110100010011: color_data = Z;
		19'b0100001110100010100: color_data = Z;
		19'b0100001110100010101: color_data = Z;
		19'b0100001110100010110: color_data = Z;
		19'b0100001110100010111: color_data = Z;
		19'b0100001110100011000: color_data = Z;
		19'b0100001110100011001: color_data = Z;
		19'b0100001110100011010: color_data = Z;
		19'b0100001110100011011: color_data = Z;
		19'b0100001110100011100: color_data = Z;
		19'b0100001110100011101: color_data = Z;
		19'b0100001110100011110: color_data = Z;
		19'b0100001110100011111: color_data = Z;
		19'b0100001110100100000: color_data = Z;
		19'b0100001110100100001: color_data = Z;
		19'b0100001110100100010: color_data = Z;
		19'b0100001110100100011: color_data = Z;
		19'b0100001110100100100: color_data = Z;
		19'b0100001110100100101: color_data = Z;
		19'b0100001110100100110: color_data = Z;
		19'b0100001110100100111: color_data = Z;
		19'b0100001110100101000: color_data = Z;
		19'b0100001110100101001: color_data = Z;
		19'b0100001110100101010: color_data = Z;
		19'b0100001110100101011: color_data = Z;
		19'b0100001110100101100: color_data = Z;
		19'b0100001110100101101: color_data = Z;
		19'b0100001110100101110: color_data = Z;
		19'b0100001110100101111: color_data = Z;
		19'b0100001110100110000: color_data = Z;
		19'b0100001110100110001: color_data = Z;
		19'b0100001110100110010: color_data = Z;
		19'b0100001110100110011: color_data = Z;
		19'b0100001110100110100: color_data = Z;
		19'b0100001110100110101: color_data = Z;
		19'b0100001110100110110: color_data = Z;
		19'b0100001110100110111: color_data = Z;
		19'b0100001110100111000: color_data = Z;
		19'b0100001110100111001: color_data = Z;
		19'b0100001110100111010: color_data = Z;
		19'b0100001110100111011: color_data = Z;
		19'b0100001110100111100: color_data = Z;
		19'b0100001110100111101: color_data = Z;
		19'b0100001110100111110: color_data = Z;
		19'b0100001110100111111: color_data = Z;
		19'b0100001110101000000: color_data = Z;
		19'b0100001110101000001: color_data = Z;
		19'b0100001110101000010: color_data = Z;
		19'b0100001110101000011: color_data = Z;
		19'b0100001110101000100: color_data = Z;
		19'b0100001110101000101: color_data = Z;
		19'b0100001110101000110: color_data = Z;
		19'b0100001110101000111: color_data = Z;
		19'b0100001110101001000: color_data = Z;
		19'b0100001110101001001: color_data = Z;
		19'b0100001110101001010: color_data = Z;
		19'b0100001110101001011: color_data = Z;
		19'b0100001110101001100: color_data = Z;
		19'b0100001110101001101: color_data = Z;
		19'b0100001110101001110: color_data = Z;
		19'b0100001110101001111: color_data = Z;
		19'b0100001110101010000: color_data = Z;
		19'b0100001110101010001: color_data = Z;
		19'b0100001110101010010: color_data = Z;
		19'b0100001110101010011: color_data = Z;
		19'b0100001110101010100: color_data = Z;
		19'b0100001110101010101: color_data = Z;
		19'b0100001110101010110: color_data = Z;
		19'b0100001110101010111: color_data = Z;
		19'b0100001110101011000: color_data = Z;
		19'b0100001110101011001: color_data = Z;
		19'b0100001110101011010: color_data = Z;
		19'b0100001110101011011: color_data = Z;
		19'b0100001110101011100: color_data = Z;
		19'b0100001110101011101: color_data = Z;
		19'b0100001110101011110: color_data = Z;
		19'b0100001110101011111: color_data = Z;
		19'b0100001110101100000: color_data = Z;
		19'b0100001110101100001: color_data = Z;
		19'b0100001110101100010: color_data = Z;
		19'b0100001110101100011: color_data = Z;
		19'b0100001110101100100: color_data = Z;
		19'b0100001110101100101: color_data = Z;
		19'b0100001110101100110: color_data = Z;
		19'b0100001110101100111: color_data = Z;
		19'b0100001110101101000: color_data = Z;
		19'b0100001110101101001: color_data = Z;
		19'b0100001110101101010: color_data = Z;
		19'b0100001110101101011: color_data = Z;
		19'b0100001110101101100: color_data = Z;
		19'b0100001110101101101: color_data = Z;
		19'b0100001110101101110: color_data = Z;
		19'b0100001110101101111: color_data = Z;
		19'b0100001110101110000: color_data = Z;
		19'b0100001110101110001: color_data = Z;
		19'b0100001110101110010: color_data = Z;
		19'b0100001110101110011: color_data = Z;
		19'b0100001110101110100: color_data = Z;
		19'b0100001110101110101: color_data = Z;
		19'b0100001110101110110: color_data = Z;
		19'b0100001110101110111: color_data = Z;
		19'b0100001110101111000: color_data = Z;
		19'b0100001110101111001: color_data = Z;
		19'b0100001110101111010: color_data = Z;
		19'b0100001110101111011: color_data = Z;
		19'b0100001110101111100: color_data = Z;
		19'b0100001110101111101: color_data = Z;
		19'b0100001110101111110: color_data = Z;
		19'b0100001110101111111: color_data = Z;
		19'b0100001110110000001: color_data = Z;
		19'b0100001110110000010: color_data = Z;
		19'b0100001110110000011: color_data = Z;
		19'b0100001110110000100: color_data = Z;
		19'b0100001110111001101: color_data = Z;
		19'b0100001110111001110: color_data = Z;
		19'b0100001110111001111: color_data = Z;
		19'b0100001110111010000: color_data = Z;
		19'b0100001110111010001: color_data = Z;
		19'b0100001110111010010: color_data = Z;
		19'b0100001110111010011: color_data = Z;
		19'b0100001110111010100: color_data = Z;
		19'b0100001110111010101: color_data = Z;
		19'b0100001110111010110: color_data = Z;
		19'b0100001110111100000: color_data = Z;
		19'b0100001110111100011: color_data = Z;
		19'b0100010000010110100: color_data = Z;
		19'b0100010000010110101: color_data = Z;
		19'b0100010000011001011: color_data = Z;
		19'b0100010000011001100: color_data = Z;
		19'b0100010000011001101: color_data = Z;
		19'b0100010000011001110: color_data = Z;
		19'b0100010000011001111: color_data = Z;
		19'b0100010000011010000: color_data = Z;
		19'b0100010000011010001: color_data = Z;
		19'b0100010000011111101: color_data = Z;
		19'b0100010000011111110: color_data = Z;
		19'b0100010000011111111: color_data = Z;
		19'b0100010000100000000: color_data = Z;
		19'b0100010000100000001: color_data = Z;
		19'b0100010000100000010: color_data = Z;
		19'b0100010000100000011: color_data = Z;
		19'b0100010000100000100: color_data = Z;
		19'b0100010000100000101: color_data = Z;
		19'b0100010000100000110: color_data = Z;
		19'b0100010000100000111: color_data = Z;
		19'b0100010000100001000: color_data = Z;
		19'b0100010000100001001: color_data = Z;
		19'b0100010000100001010: color_data = Z;
		19'b0100010000100001011: color_data = Z;
		19'b0100010000100001100: color_data = Z;
		19'b0100010000100001101: color_data = Z;
		19'b0100010000100001110: color_data = Z;
		19'b0100010000100001111: color_data = Z;
		19'b0100010000100010000: color_data = Z;
		19'b0100010000100010001: color_data = Z;
		19'b0100010000100010010: color_data = Z;
		19'b0100010000100010011: color_data = Z;
		19'b0100010000100010100: color_data = Z;
		19'b0100010000100010101: color_data = Z;
		19'b0100010000100010110: color_data = Z;
		19'b0100010000100010111: color_data = Z;
		19'b0100010000100011000: color_data = Z;
		19'b0100010000100011001: color_data = Z;
		19'b0100010000100011010: color_data = Z;
		19'b0100010000100011011: color_data = Z;
		19'b0100010000100011100: color_data = Z;
		19'b0100010000100011101: color_data = Z;
		19'b0100010000100011110: color_data = Z;
		19'b0100010000100011111: color_data = Z;
		19'b0100010000100100000: color_data = Z;
		19'b0100010000100100001: color_data = Z;
		19'b0100010000100100010: color_data = Z;
		19'b0100010000100100011: color_data = Z;
		19'b0100010000100100100: color_data = Z;
		19'b0100010000100100101: color_data = Z;
		19'b0100010000100100110: color_data = Z;
		19'b0100010000100100111: color_data = Z;
		19'b0100010000100101000: color_data = Z;
		19'b0100010000100101001: color_data = Z;
		19'b0100010000100101010: color_data = Z;
		19'b0100010000100101011: color_data = Z;
		19'b0100010000100101100: color_data = Z;
		19'b0100010000100101101: color_data = Z;
		19'b0100010000100101110: color_data = Z;
		19'b0100010000100101111: color_data = Z;
		19'b0100010000100110000: color_data = Z;
		19'b0100010000100110001: color_data = Z;
		19'b0100010000100110010: color_data = Z;
		19'b0100010000100110011: color_data = Z;
		19'b0100010000100110100: color_data = Z;
		19'b0100010000100110101: color_data = Z;
		19'b0100010000100110110: color_data = Z;
		19'b0100010000100110111: color_data = Z;
		19'b0100010000100111000: color_data = Z;
		19'b0100010000100111001: color_data = Z;
		19'b0100010000100111010: color_data = Z;
		19'b0100010000100111011: color_data = Z;
		19'b0100010000100111100: color_data = Z;
		19'b0100010000100111101: color_data = Z;
		19'b0100010000100111110: color_data = Z;
		19'b0100010000100111111: color_data = Z;
		19'b0100010000101000000: color_data = Z;
		19'b0100010000101000001: color_data = Z;
		19'b0100010000101000010: color_data = Z;
		19'b0100010000101000011: color_data = Z;
		19'b0100010000101000100: color_data = Z;
		19'b0100010000101000101: color_data = Z;
		19'b0100010000101000110: color_data = Z;
		19'b0100010000101000111: color_data = Z;
		19'b0100010000101001000: color_data = Z;
		19'b0100010000101001001: color_data = Z;
		19'b0100010000101001010: color_data = Z;
		19'b0100010000101001011: color_data = Z;
		19'b0100010000101001100: color_data = Z;
		19'b0100010000101001101: color_data = Z;
		19'b0100010000101001110: color_data = Z;
		19'b0100010000101001111: color_data = Z;
		19'b0100010000101010000: color_data = Z;
		19'b0100010000101010001: color_data = Z;
		19'b0100010000101010010: color_data = Z;
		19'b0100010000101010011: color_data = Z;
		19'b0100010000101010100: color_data = Z;
		19'b0100010000101010101: color_data = Z;
		19'b0100010000101010110: color_data = Z;
		19'b0100010000101010111: color_data = Z;
		19'b0100010000101011000: color_data = Z;
		19'b0100010000101011001: color_data = Z;
		19'b0100010000101011010: color_data = Z;
		19'b0100010000101011011: color_data = Z;
		19'b0100010000101011100: color_data = Z;
		19'b0100010000101011101: color_data = Z;
		19'b0100010000101011110: color_data = Z;
		19'b0100010000101011111: color_data = Z;
		19'b0100010000101100000: color_data = Z;
		19'b0100010000101100001: color_data = Z;
		19'b0100010000101100010: color_data = Z;
		19'b0100010000101100011: color_data = Z;
		19'b0100010000101100100: color_data = Z;
		19'b0100010000101100101: color_data = Z;
		19'b0100010000101100110: color_data = Z;
		19'b0100010000101100111: color_data = Z;
		19'b0100010000101101000: color_data = Z;
		19'b0100010000101101001: color_data = Z;
		19'b0100010000101101010: color_data = Z;
		19'b0100010000101101011: color_data = Z;
		19'b0100010000101101100: color_data = Z;
		19'b0100010000101101101: color_data = Z;
		19'b0100010000101101110: color_data = Z;
		19'b0100010000101101111: color_data = Z;
		19'b0100010000101110000: color_data = Z;
		19'b0100010000101110001: color_data = Z;
		19'b0100010000101110010: color_data = Z;
		19'b0100010000101110011: color_data = Z;
		19'b0100010000101110100: color_data = Z;
		19'b0100010000101110101: color_data = Z;
		19'b0100010000101110110: color_data = Z;
		19'b0100010000101110111: color_data = Z;
		19'b0100010000101111000: color_data = Z;
		19'b0100010000101111001: color_data = Z;
		19'b0100010000101111010: color_data = Z;
		19'b0100010000101111011: color_data = Z;
		19'b0100010000101111100: color_data = Z;
		19'b0100010000101111101: color_data = Z;
		19'b0100010000101111110: color_data = Z;
		19'b0100010000101111111: color_data = Z;
		19'b0100010000110000000: color_data = Z;
		19'b0100010000110000001: color_data = Z;
		19'b0100010000110000010: color_data = Z;
		19'b0100010000110000011: color_data = Z;
		19'b0100010000110000100: color_data = Z;
		19'b0100010000111001101: color_data = Z;
		19'b0100010000111001110: color_data = Z;
		19'b0100010000111001111: color_data = Z;
		19'b0100010000111010000: color_data = Z;
		19'b0100010000111010001: color_data = Z;
		19'b0100010000111010010: color_data = Z;
		19'b0100010000111010011: color_data = Z;
		19'b0100010000111010100: color_data = Z;
		19'b0100010000111010101: color_data = Z;
		19'b0100010000111010110: color_data = Z;
		19'b0100010000111010111: color_data = Z;
		19'b0100010010010110100: color_data = Z;
		19'b0100010010011001011: color_data = Z;
		19'b0100010010011001100: color_data = Z;
		19'b0100010010011001101: color_data = Z;
		19'b0100010010011001110: color_data = Z;
		19'b0100010010011001111: color_data = Z;
		19'b0100010010011010000: color_data = Z;
		19'b0100010010011111110: color_data = Z;
		19'b0100010010011111111: color_data = Z;
		19'b0100010010100000000: color_data = Z;
		19'b0100010010100000001: color_data = Z;
		19'b0100010010100000010: color_data = Z;
		19'b0100010010100000011: color_data = Z;
		19'b0100010010100000100: color_data = Z;
		19'b0100010010100000101: color_data = Z;
		19'b0100010010100000110: color_data = Z;
		19'b0100010010100000111: color_data = Z;
		19'b0100010010100001000: color_data = Z;
		19'b0100010010100001001: color_data = Z;
		19'b0100010010100001010: color_data = Z;
		19'b0100010010100001011: color_data = Z;
		19'b0100010010100001100: color_data = Z;
		19'b0100010010100001101: color_data = Z;
		19'b0100010010100001110: color_data = Z;
		19'b0100010010100001111: color_data = Z;
		19'b0100010010100010000: color_data = Z;
		19'b0100010010100010001: color_data = Z;
		19'b0100010010100010010: color_data = Z;
		19'b0100010010100010011: color_data = Z;
		19'b0100010010100010100: color_data = Z;
		19'b0100010010100010101: color_data = Z;
		19'b0100010010100010110: color_data = Z;
		19'b0100010010100010111: color_data = Z;
		19'b0100010010100011000: color_data = Z;
		19'b0100010010100011001: color_data = Z;
		19'b0100010010100011010: color_data = Z;
		19'b0100010010100011011: color_data = Z;
		19'b0100010010100011100: color_data = Z;
		19'b0100010010100011101: color_data = Z;
		19'b0100010010100011110: color_data = Z;
		19'b0100010010100011111: color_data = Z;
		19'b0100010010100100000: color_data = Z;
		19'b0100010010100100001: color_data = Z;
		19'b0100010010100100010: color_data = Z;
		19'b0100010010100100011: color_data = Z;
		19'b0100010010100100100: color_data = Z;
		19'b0100010010100100101: color_data = Z;
		19'b0100010010100100110: color_data = Z;
		19'b0100010010100100111: color_data = Z;
		19'b0100010010100101000: color_data = Z;
		19'b0100010010100101001: color_data = Z;
		19'b0100010010100101010: color_data = Z;
		19'b0100010010100101011: color_data = Z;
		19'b0100010010100101100: color_data = Z;
		19'b0100010010100101101: color_data = Z;
		19'b0100010010100101110: color_data = Z;
		19'b0100010010100101111: color_data = Z;
		19'b0100010010100110000: color_data = Z;
		19'b0100010010100110001: color_data = Z;
		19'b0100010010100110010: color_data = Z;
		19'b0100010010100110011: color_data = Z;
		19'b0100010010100110100: color_data = Z;
		19'b0100010010100110101: color_data = Z;
		19'b0100010010100110110: color_data = Z;
		19'b0100010010100110111: color_data = Z;
		19'b0100010010100111000: color_data = Z;
		19'b0100010010100111001: color_data = Z;
		19'b0100010010100111010: color_data = Z;
		19'b0100010010100111011: color_data = Z;
		19'b0100010010100111100: color_data = Z;
		19'b0100010010100111101: color_data = Z;
		19'b0100010010100111110: color_data = Z;
		19'b0100010010100111111: color_data = Z;
		19'b0100010010101000000: color_data = Z;
		19'b0100010010101000001: color_data = Z;
		19'b0100010010101000010: color_data = Z;
		19'b0100010010101000011: color_data = Z;
		19'b0100010010101000100: color_data = Z;
		19'b0100010010101000101: color_data = Z;
		19'b0100010010101000110: color_data = Z;
		19'b0100010010101000111: color_data = Z;
		19'b0100010010101001000: color_data = Z;
		19'b0100010010101001001: color_data = Z;
		19'b0100010010101001010: color_data = Z;
		19'b0100010010101001011: color_data = Z;
		19'b0100010010101001100: color_data = Z;
		19'b0100010010101001101: color_data = Z;
		19'b0100010010101001110: color_data = Z;
		19'b0100010010101001111: color_data = Z;
		19'b0100010010101010000: color_data = Z;
		19'b0100010010101010001: color_data = Z;
		19'b0100010010101010010: color_data = Z;
		19'b0100010010101010011: color_data = Z;
		19'b0100010010101010100: color_data = Z;
		19'b0100010010101010101: color_data = Z;
		19'b0100010010101010110: color_data = Z;
		19'b0100010010101010111: color_data = Z;
		19'b0100010010101011000: color_data = Z;
		19'b0100010010101011001: color_data = Z;
		19'b0100010010101011010: color_data = Z;
		19'b0100010010101011011: color_data = Z;
		19'b0100010010101011100: color_data = Z;
		19'b0100010010101011101: color_data = Z;
		19'b0100010010101011110: color_data = Z;
		19'b0100010010101011111: color_data = Z;
		19'b0100010010101100000: color_data = Z;
		19'b0100010010101100001: color_data = Z;
		19'b0100010010101100010: color_data = Z;
		19'b0100010010101100011: color_data = Z;
		19'b0100010010101100100: color_data = Z;
		19'b0100010010101100101: color_data = Z;
		19'b0100010010101100110: color_data = Z;
		19'b0100010010101100111: color_data = Z;
		19'b0100010010101101000: color_data = Z;
		19'b0100010010101101001: color_data = Z;
		19'b0100010010101101010: color_data = Z;
		19'b0100010010101101011: color_data = Z;
		19'b0100010010101101100: color_data = Z;
		19'b0100010010101101101: color_data = Z;
		19'b0100010010101101110: color_data = Z;
		19'b0100010010101101111: color_data = Z;
		19'b0100010010101110000: color_data = Z;
		19'b0100010010101110001: color_data = Z;
		19'b0100010010101110010: color_data = Z;
		19'b0100010010101110011: color_data = Z;
		19'b0100010010101110100: color_data = Z;
		19'b0100010010101110101: color_data = Z;
		19'b0100010010101110110: color_data = Z;
		19'b0100010010101110111: color_data = Z;
		19'b0100010010101111000: color_data = Z;
		19'b0100010010101111001: color_data = Z;
		19'b0100010010101111010: color_data = Z;
		19'b0100010010101111011: color_data = Z;
		19'b0100010010101111100: color_data = Z;
		19'b0100010010101111101: color_data = Z;
		19'b0100010010101111110: color_data = Z;
		19'b0100010010101111111: color_data = Z;
		19'b0100010010110000000: color_data = Z;
		19'b0100010010110000001: color_data = Z;
		19'b0100010010110000010: color_data = Z;
		19'b0100010010110000011: color_data = Z;
		19'b0100010010111001101: color_data = Z;
		19'b0100010010111001110: color_data = Z;
		19'b0100010010111001111: color_data = Z;
		19'b0100010010111010000: color_data = Z;
		19'b0100010010111010001: color_data = Z;
		19'b0100010010111010010: color_data = Z;
		19'b0100010010111010011: color_data = Z;
		19'b0100010010111010100: color_data = Z;
		19'b0100010010111010101: color_data = Z;
		19'b0100010010111010110: color_data = Z;
		19'b0100010010111010111: color_data = Z;
		19'b0100010100011001011: color_data = Z;
		19'b0100010100011001100: color_data = Z;
		19'b0100010100011001101: color_data = Z;
		19'b0100010100100000000: color_data = Z;
		19'b0100010100100000001: color_data = Z;
		19'b0100010100100000010: color_data = Z;
		19'b0100010100100000011: color_data = Z;
		19'b0100010100100000100: color_data = Z;
		19'b0100010100100000101: color_data = Z;
		19'b0100010100100000110: color_data = Z;
		19'b0100010100100000111: color_data = Z;
		19'b0100010100100001000: color_data = Z;
		19'b0100010100100001001: color_data = Z;
		19'b0100010100100001010: color_data = Z;
		19'b0100010100100001011: color_data = Z;
		19'b0100010100100001100: color_data = Z;
		19'b0100010100100001101: color_data = Z;
		19'b0100010100100001110: color_data = Z;
		19'b0100010100100001111: color_data = Z;
		19'b0100010100100010000: color_data = Z;
		19'b0100010100100010001: color_data = Z;
		19'b0100010100100010010: color_data = Z;
		19'b0100010100100010011: color_data = Z;
		19'b0100010100100010100: color_data = Z;
		19'b0100010100100010101: color_data = Z;
		19'b0100010100100010110: color_data = Z;
		19'b0100010100100010111: color_data = Z;
		19'b0100010100100011000: color_data = Z;
		19'b0100010100100011001: color_data = Z;
		19'b0100010100100011010: color_data = Z;
		19'b0100010100100011011: color_data = Z;
		19'b0100010100100011100: color_data = Z;
		19'b0100010100100011101: color_data = Z;
		19'b0100010100100011110: color_data = Z;
		19'b0100010100100011111: color_data = Z;
		19'b0100010100100100000: color_data = Z;
		19'b0100010100100100001: color_data = Z;
		19'b0100010100100100010: color_data = Z;
		19'b0100010100100100011: color_data = Z;
		19'b0100010100100100100: color_data = Z;
		19'b0100010100100100101: color_data = Z;
		19'b0100010100100100110: color_data = Z;
		19'b0100010100100100111: color_data = Z;
		19'b0100010100100101000: color_data = Z;
		19'b0100010100100101001: color_data = Z;
		19'b0100010100100101010: color_data = Z;
		19'b0100010100100101011: color_data = Z;
		19'b0100010100100101100: color_data = Z;
		19'b0100010100100101101: color_data = Z;
		19'b0100010100100101110: color_data = Z;
		19'b0100010100100101111: color_data = Z;
		19'b0100010100100110000: color_data = Z;
		19'b0100010100100110001: color_data = Z;
		19'b0100010100100110010: color_data = Z;
		19'b0100010100100110011: color_data = Z;
		19'b0100010100100110100: color_data = Z;
		19'b0100010100100110101: color_data = Z;
		19'b0100010100100110110: color_data = Z;
		19'b0100010100100110111: color_data = Z;
		19'b0100010100100111000: color_data = Z;
		19'b0100010100100111001: color_data = Z;
		19'b0100010100100111010: color_data = Z;
		19'b0100010100100111011: color_data = Z;
		19'b0100010100100111100: color_data = Z;
		19'b0100010100100111101: color_data = Z;
		19'b0100010100100111110: color_data = Z;
		19'b0100010100100111111: color_data = Z;
		19'b0100010100101000000: color_data = Z;
		19'b0100010100101000001: color_data = Z;
		19'b0100010100101000010: color_data = Z;
		19'b0100010100101000011: color_data = Z;
		19'b0100010100101000100: color_data = Z;
		19'b0100010100101000101: color_data = Z;
		19'b0100010100101000110: color_data = Z;
		19'b0100010100101000111: color_data = Z;
		19'b0100010100101001000: color_data = Z;
		19'b0100010100101001001: color_data = Z;
		19'b0100010100101001010: color_data = Z;
		19'b0100010100101001011: color_data = Z;
		19'b0100010100101001100: color_data = Z;
		19'b0100010100101001101: color_data = Z;
		19'b0100010100101001110: color_data = Z;
		19'b0100010100101001111: color_data = Z;
		19'b0100010100101010000: color_data = Z;
		19'b0100010100101010001: color_data = Z;
		19'b0100010100101010010: color_data = Z;
		19'b0100010100101010011: color_data = Z;
		19'b0100010100101010100: color_data = Z;
		19'b0100010100101010101: color_data = Z;
		19'b0100010100101010110: color_data = Z;
		19'b0100010100101010111: color_data = Z;
		19'b0100010100101011000: color_data = Z;
		19'b0100010100101011001: color_data = Z;
		19'b0100010100101011010: color_data = Z;
		19'b0100010100101011011: color_data = Z;
		19'b0100010100101011100: color_data = Z;
		19'b0100010100101011101: color_data = Z;
		19'b0100010100101011110: color_data = Z;
		19'b0100010100101011111: color_data = Z;
		19'b0100010100101100000: color_data = Z;
		19'b0100010100101100001: color_data = Z;
		19'b0100010100101100010: color_data = Z;
		19'b0100010100101100011: color_data = Z;
		19'b0100010100101100100: color_data = Z;
		19'b0100010100101100101: color_data = Z;
		19'b0100010100101100110: color_data = Z;
		19'b0100010100101100111: color_data = Z;
		19'b0100010100101101000: color_data = Z;
		19'b0100010100101101001: color_data = Z;
		19'b0100010100101101010: color_data = Z;
		19'b0100010100101101011: color_data = Z;
		19'b0100010100101101100: color_data = Z;
		19'b0100010100101101101: color_data = Z;
		19'b0100010100101101110: color_data = Z;
		19'b0100010100101101111: color_data = Z;
		19'b0100010100101110000: color_data = Z;
		19'b0100010100101110001: color_data = Z;
		19'b0100010100101110010: color_data = Z;
		19'b0100010100101110011: color_data = Z;
		19'b0100010100101110100: color_data = Z;
		19'b0100010100101110101: color_data = Z;
		19'b0100010100101110110: color_data = Z;
		19'b0100010100101110111: color_data = Z;
		19'b0100010100101111000: color_data = Z;
		19'b0100010100101111001: color_data = Z;
		19'b0100010100101111010: color_data = Z;
		19'b0100010100101111011: color_data = Z;
		19'b0100010100101111100: color_data = Z;
		19'b0100010100101111101: color_data = Z;
		19'b0100010100101111110: color_data = Z;
		19'b0100010100101111111: color_data = Z;
		19'b0100010100110000000: color_data = Z;
		19'b0100010100110000001: color_data = Z;
		19'b0100010100110000010: color_data = Z;
		19'b0100010100110000011: color_data = Z;
		19'b0100010100111001110: color_data = Z;
		19'b0100010100111001111: color_data = Z;
		19'b0100010100111010000: color_data = Z;
		19'b0100010100111010001: color_data = Z;
		19'b0100010100111010010: color_data = Z;
		19'b0100010100111010011: color_data = Z;
		19'b0100010100111010100: color_data = Z;
		19'b0100010100111010101: color_data = Z;
		19'b0100010100111010110: color_data = Z;
		19'b0100010100111010111: color_data = Z;
		19'b0100010100111011000: color_data = Z;
		19'b0100010110011001000: color_data = Z;
		19'b0100010110011001001: color_data = Z;
		19'b0100010110011001010: color_data = Z;
		19'b0100010110100000000: color_data = Z;
		19'b0100010110100000001: color_data = Z;
		19'b0100010110100000010: color_data = Z;
		19'b0100010110100000011: color_data = Z;
		19'b0100010110100000100: color_data = Z;
		19'b0100010110100000101: color_data = Z;
		19'b0100010110100000110: color_data = Z;
		19'b0100010110100000111: color_data = Z;
		19'b0100010110100001000: color_data = Z;
		19'b0100010110100001001: color_data = Z;
		19'b0100010110100001010: color_data = Z;
		19'b0100010110100001011: color_data = Z;
		19'b0100010110100001100: color_data = Z;
		19'b0100010110100001101: color_data = Z;
		19'b0100010110100001110: color_data = Z;
		19'b0100010110100001111: color_data = Z;
		19'b0100010110100010000: color_data = Z;
		19'b0100010110100010001: color_data = Z;
		19'b0100010110100010010: color_data = Z;
		19'b0100010110100010011: color_data = Z;
		19'b0100010110100010100: color_data = Z;
		19'b0100010110100010101: color_data = Z;
		19'b0100010110100010110: color_data = Z;
		19'b0100010110100010111: color_data = Z;
		19'b0100010110100011000: color_data = Z;
		19'b0100010110100011001: color_data = Z;
		19'b0100010110100011010: color_data = Z;
		19'b0100010110100011011: color_data = Z;
		19'b0100010110100011100: color_data = Z;
		19'b0100010110100011101: color_data = Z;
		19'b0100010110100011110: color_data = Z;
		19'b0100010110100011111: color_data = Z;
		19'b0100010110100100000: color_data = Z;
		19'b0100010110100100001: color_data = Z;
		19'b0100010110100100010: color_data = Z;
		19'b0100010110100100011: color_data = Z;
		19'b0100010110100100100: color_data = Z;
		19'b0100010110100100101: color_data = Z;
		19'b0100010110100100110: color_data = Z;
		19'b0100010110100100111: color_data = Z;
		19'b0100010110100101000: color_data = Z;
		19'b0100010110100101001: color_data = Z;
		19'b0100010110100101010: color_data = Z;
		19'b0100010110100101011: color_data = Z;
		19'b0100010110100101100: color_data = Z;
		19'b0100010110100101101: color_data = Z;
		19'b0100010110100101110: color_data = Z;
		19'b0100010110100101111: color_data = Z;
		19'b0100010110100110000: color_data = Z;
		19'b0100010110100110001: color_data = Z;
		19'b0100010110100110010: color_data = Z;
		19'b0100010110100110011: color_data = Z;
		19'b0100010110100110100: color_data = Z;
		19'b0100010110100110101: color_data = Z;
		19'b0100010110100110110: color_data = Z;
		19'b0100010110100110111: color_data = Z;
		19'b0100010110100111000: color_data = Z;
		19'b0100010110100111001: color_data = Z;
		19'b0100010110100111010: color_data = Z;
		19'b0100010110100111011: color_data = Z;
		19'b0100010110100111100: color_data = Z;
		19'b0100010110100111101: color_data = Z;
		19'b0100010110100111110: color_data = Z;
		19'b0100010110100111111: color_data = Z;
		19'b0100010110101000000: color_data = Z;
		19'b0100010110101000001: color_data = Z;
		19'b0100010110101000010: color_data = Z;
		19'b0100010110101000011: color_data = Z;
		19'b0100010110101000100: color_data = Z;
		19'b0100010110101000101: color_data = Z;
		19'b0100010110101000110: color_data = Z;
		19'b0100010110101000111: color_data = Z;
		19'b0100010110101001000: color_data = Z;
		19'b0100010110101001001: color_data = Z;
		19'b0100010110101001010: color_data = Z;
		19'b0100010110101001011: color_data = Z;
		19'b0100010110101001100: color_data = Z;
		19'b0100010110101001101: color_data = Z;
		19'b0100010110101001110: color_data = Z;
		19'b0100010110101001111: color_data = Z;
		19'b0100010110101010000: color_data = Z;
		19'b0100010110101010001: color_data = Z;
		19'b0100010110101010010: color_data = Z;
		19'b0100010110101010011: color_data = Z;
		19'b0100010110101010100: color_data = Z;
		19'b0100010110101010101: color_data = Z;
		19'b0100010110101010110: color_data = Z;
		19'b0100010110101010111: color_data = Z;
		19'b0100010110101011000: color_data = Z;
		19'b0100010110101011001: color_data = Z;
		19'b0100010110101011010: color_data = Z;
		19'b0100010110101011011: color_data = Z;
		19'b0100010110101011100: color_data = Z;
		19'b0100010110101011101: color_data = Z;
		19'b0100010110101011110: color_data = Z;
		19'b0100010110101011111: color_data = Z;
		19'b0100010110101100000: color_data = Z;
		19'b0100010110101100001: color_data = Z;
		19'b0100010110101100010: color_data = Z;
		19'b0100010110101100011: color_data = Z;
		19'b0100010110101100100: color_data = Z;
		19'b0100010110101100101: color_data = Z;
		19'b0100010110101100110: color_data = Z;
		19'b0100010110101100111: color_data = Z;
		19'b0100010110101101000: color_data = Z;
		19'b0100010110101101001: color_data = Z;
		19'b0100010110101101010: color_data = Z;
		19'b0100010110101101011: color_data = Z;
		19'b0100010110101101100: color_data = Z;
		19'b0100010110101101101: color_data = Z;
		19'b0100010110101101110: color_data = Z;
		19'b0100010110101101111: color_data = Z;
		19'b0100010110101110000: color_data = Z;
		19'b0100010110101110001: color_data = Z;
		19'b0100010110101110010: color_data = Z;
		19'b0100010110101110011: color_data = Z;
		19'b0100010110101110100: color_data = Z;
		19'b0100010110101110101: color_data = Z;
		19'b0100010110101110110: color_data = Z;
		19'b0100010110101110111: color_data = Z;
		19'b0100010110101111000: color_data = Z;
		19'b0100010110101111001: color_data = Z;
		19'b0100010110101111010: color_data = Z;
		19'b0100010110101111011: color_data = Z;
		19'b0100010110101111100: color_data = Z;
		19'b0100010110101111101: color_data = Z;
		19'b0100010110101111110: color_data = Z;
		19'b0100010110101111111: color_data = Z;
		19'b0100010110110000000: color_data = Z;
		19'b0100010110110000001: color_data = Z;
		19'b0100010110110000010: color_data = Z;
		19'b0100010110110000011: color_data = Z;
		19'b0100010110111001110: color_data = Z;
		19'b0100010110111001111: color_data = Z;
		19'b0100010110111010000: color_data = Z;
		19'b0100010110111010001: color_data = Z;
		19'b0100010110111010010: color_data = Z;
		19'b0100010110111010011: color_data = Z;
		19'b0100010110111010100: color_data = Z;
		19'b0100010110111010101: color_data = Z;
		19'b0100010110111010110: color_data = Z;
		19'b0100010110111010111: color_data = Z;
		19'b0100011000011000111: color_data = Z;
		19'b0100011000011001000: color_data = Z;
		19'b0100011000011001001: color_data = Z;
		19'b0100011000100000011: color_data = Z;
		19'b0100011000100000100: color_data = Z;
		19'b0100011000100000101: color_data = Z;
		19'b0100011000100000110: color_data = Z;
		19'b0100011000100000111: color_data = Z;
		19'b0100011000100001000: color_data = Z;
		19'b0100011000100001001: color_data = Z;
		19'b0100011000100001010: color_data = Z;
		19'b0100011000100001011: color_data = Z;
		19'b0100011000100001100: color_data = Z;
		19'b0100011000100001101: color_data = Z;
		19'b0100011000100001110: color_data = Z;
		19'b0100011000100001111: color_data = Z;
		19'b0100011000100010000: color_data = Z;
		19'b0100011000100010001: color_data = Z;
		19'b0100011000100010010: color_data = Z;
		19'b0100011000100010011: color_data = Z;
		19'b0100011000100010100: color_data = Z;
		19'b0100011000100010101: color_data = Z;
		19'b0100011000100010110: color_data = Z;
		19'b0100011000100010111: color_data = Z;
		19'b0100011000100011000: color_data = Z;
		19'b0100011000100011001: color_data = Z;
		19'b0100011000100011010: color_data = Z;
		19'b0100011000100011011: color_data = Z;
		19'b0100011000100011100: color_data = Z;
		19'b0100011000100011101: color_data = Z;
		19'b0100011000100011110: color_data = Z;
		19'b0100011000100011111: color_data = Z;
		19'b0100011000100100000: color_data = Z;
		19'b0100011000100100001: color_data = Z;
		19'b0100011000100100010: color_data = Z;
		19'b0100011000100100011: color_data = Z;
		19'b0100011000100100100: color_data = Z;
		19'b0100011000100100101: color_data = Z;
		19'b0100011000100100110: color_data = Z;
		19'b0100011000100100111: color_data = Z;
		19'b0100011000100101000: color_data = Z;
		19'b0100011000100101001: color_data = Z;
		19'b0100011000100101010: color_data = Z;
		19'b0100011000100101011: color_data = Z;
		19'b0100011000100101100: color_data = Z;
		19'b0100011000100101101: color_data = Z;
		19'b0100011000100101110: color_data = Z;
		19'b0100011000100101111: color_data = Z;
		19'b0100011000100110000: color_data = Z;
		19'b0100011000100110001: color_data = Z;
		19'b0100011000100110010: color_data = Z;
		19'b0100011000100110011: color_data = Z;
		19'b0100011000100110100: color_data = Z;
		19'b0100011000100110101: color_data = Z;
		19'b0100011000100110110: color_data = Z;
		19'b0100011000100110111: color_data = Z;
		19'b0100011000100111000: color_data = Z;
		19'b0100011000100111001: color_data = Z;
		19'b0100011000100111010: color_data = Z;
		19'b0100011000100111011: color_data = Z;
		19'b0100011000100111100: color_data = Z;
		19'b0100011000100111101: color_data = Z;
		19'b0100011000100111110: color_data = Z;
		19'b0100011000100111111: color_data = Z;
		19'b0100011000101000000: color_data = Z;
		19'b0100011000101000001: color_data = Z;
		19'b0100011000101000010: color_data = Z;
		19'b0100011000101000011: color_data = Z;
		19'b0100011000101000100: color_data = Z;
		19'b0100011000101000101: color_data = Z;
		19'b0100011000101000110: color_data = Z;
		19'b0100011000101000111: color_data = Z;
		19'b0100011000101001000: color_data = Z;
		19'b0100011000101001001: color_data = Z;
		19'b0100011000101001010: color_data = Z;
		19'b0100011000101001011: color_data = Z;
		19'b0100011000101001100: color_data = Z;
		19'b0100011000101001101: color_data = Z;
		19'b0100011000101001110: color_data = Z;
		19'b0100011000101001111: color_data = Z;
		19'b0100011000101010000: color_data = Z;
		19'b0100011000101010001: color_data = Z;
		19'b0100011000101010010: color_data = Z;
		19'b0100011000101010011: color_data = Z;
		19'b0100011000101010100: color_data = Z;
		19'b0100011000101010101: color_data = Z;
		19'b0100011000101010110: color_data = Z;
		19'b0100011000101010111: color_data = Z;
		19'b0100011000101011000: color_data = Z;
		19'b0100011000101011001: color_data = Z;
		19'b0100011000101011010: color_data = Z;
		19'b0100011000101011011: color_data = Z;
		19'b0100011000101011100: color_data = Z;
		19'b0100011000101011101: color_data = Z;
		19'b0100011000101011110: color_data = Z;
		19'b0100011000101011111: color_data = Z;
		19'b0100011000101100000: color_data = Z;
		19'b0100011000101100001: color_data = Z;
		19'b0100011000101100010: color_data = Z;
		19'b0100011000101100011: color_data = Z;
		19'b0100011000101100100: color_data = Z;
		19'b0100011000101100101: color_data = Z;
		19'b0100011000101100110: color_data = Z;
		19'b0100011000101100111: color_data = Z;
		19'b0100011000101101000: color_data = Z;
		19'b0100011000101101001: color_data = Z;
		19'b0100011000101101010: color_data = Z;
		19'b0100011000101101011: color_data = Z;
		19'b0100011000101101100: color_data = Z;
		19'b0100011000101101101: color_data = Z;
		19'b0100011000101101110: color_data = Z;
		19'b0100011000101101111: color_data = Z;
		19'b0100011000101110000: color_data = Z;
		19'b0100011000101110001: color_data = Z;
		19'b0100011000101110010: color_data = Z;
		19'b0100011000101110011: color_data = Z;
		19'b0100011000101110100: color_data = Z;
		19'b0100011000101110101: color_data = Z;
		19'b0100011000101110110: color_data = Z;
		19'b0100011000101110111: color_data = Z;
		19'b0100011000101111000: color_data = Z;
		19'b0100011000101111001: color_data = Z;
		19'b0100011000101111010: color_data = Z;
		19'b0100011000101111011: color_data = Z;
		19'b0100011000101111100: color_data = Z;
		19'b0100011000101111101: color_data = Z;
		19'b0100011000101111110: color_data = Z;
		19'b0100011000101111111: color_data = Z;
		19'b0100011000110000000: color_data = Z;
		19'b0100011000110000001: color_data = Z;
		19'b0100011000110000010: color_data = Z;
		19'b0100011000111001110: color_data = Z;
		19'b0100011000111001111: color_data = Z;
		19'b0100011000111010000: color_data = Z;
		19'b0100011000111010001: color_data = Z;
		19'b0100011000111010010: color_data = Z;
		19'b0100011000111010011: color_data = Z;
		19'b0100011000111010100: color_data = Z;
		19'b0100011000111010101: color_data = Z;
		19'b0100011000111010110: color_data = Z;
		19'b0100011000111010111: color_data = Z;
		19'b0100011010100000100: color_data = Z;
		19'b0100011010100000101: color_data = Z;
		19'b0100011010100000110: color_data = Z;
		19'b0100011010100000111: color_data = Z;
		19'b0100011010100001000: color_data = Z;
		19'b0100011010100001001: color_data = Z;
		19'b0100011010100001010: color_data = Z;
		19'b0100011010100001011: color_data = Z;
		19'b0100011010100001100: color_data = Z;
		19'b0100011010100001101: color_data = Z;
		19'b0100011010100001110: color_data = Z;
		19'b0100011010100001111: color_data = Z;
		19'b0100011010100010000: color_data = Z;
		19'b0100011010100010001: color_data = Z;
		19'b0100011010100010010: color_data = Z;
		19'b0100011010100010011: color_data = Z;
		19'b0100011010100010100: color_data = Z;
		19'b0100011010100010101: color_data = Z;
		19'b0100011010100010110: color_data = Z;
		19'b0100011010100010111: color_data = Z;
		19'b0100011010100011000: color_data = Z;
		19'b0100011010100011001: color_data = Z;
		19'b0100011010100011010: color_data = Z;
		19'b0100011010100011011: color_data = Z;
		19'b0100011010100011100: color_data = Z;
		19'b0100011010100011101: color_data = Z;
		19'b0100011010100011110: color_data = Z;
		19'b0100011010100011111: color_data = Z;
		19'b0100011010100100000: color_data = Z;
		19'b0100011010100100001: color_data = Z;
		19'b0100011010100100010: color_data = Z;
		19'b0100011010100100011: color_data = Z;
		19'b0100011010100100100: color_data = Z;
		19'b0100011010100100101: color_data = Z;
		19'b0100011010100100110: color_data = Z;
		19'b0100011010100100111: color_data = Z;
		19'b0100011010100101000: color_data = Z;
		19'b0100011010100101001: color_data = Z;
		19'b0100011010100101010: color_data = Z;
		19'b0100011010100101011: color_data = Z;
		19'b0100011010100101100: color_data = Z;
		19'b0100011010100101101: color_data = Z;
		19'b0100011010100101110: color_data = Z;
		19'b0100011010100101111: color_data = Z;
		19'b0100011010100110000: color_data = Z;
		19'b0100011010100110001: color_data = Z;
		19'b0100011010100110010: color_data = Z;
		19'b0100011010100110011: color_data = Z;
		19'b0100011010100110100: color_data = Z;
		19'b0100011010100110101: color_data = Z;
		19'b0100011010100110110: color_data = Z;
		19'b0100011010100110111: color_data = Z;
		19'b0100011010100111000: color_data = Z;
		19'b0100011010100111001: color_data = Z;
		19'b0100011010100111010: color_data = Z;
		19'b0100011010100111011: color_data = Z;
		19'b0100011010100111100: color_data = Z;
		19'b0100011010100111101: color_data = Z;
		19'b0100011010100111110: color_data = Z;
		19'b0100011010100111111: color_data = Z;
		19'b0100011010101000000: color_data = Z;
		19'b0100011010101000001: color_data = Z;
		19'b0100011010101000010: color_data = Z;
		19'b0100011010101000011: color_data = Z;
		19'b0100011010101000100: color_data = Z;
		19'b0100011010101000101: color_data = Z;
		19'b0100011010101000110: color_data = Z;
		19'b0100011010101000111: color_data = Z;
		19'b0100011010101001000: color_data = Z;
		19'b0100011010101001001: color_data = Z;
		19'b0100011010101001010: color_data = Z;
		19'b0100011010101001011: color_data = Z;
		19'b0100011010101001100: color_data = Z;
		19'b0100011010101001101: color_data = Z;
		19'b0100011010101001110: color_data = Z;
		19'b0100011010101001111: color_data = Z;
		19'b0100011010101010000: color_data = Z;
		19'b0100011010101010001: color_data = Z;
		19'b0100011010101010010: color_data = Z;
		19'b0100011010101010011: color_data = Z;
		19'b0100011010101010100: color_data = Z;
		19'b0100011010101010101: color_data = Z;
		19'b0100011010101010110: color_data = Z;
		19'b0100011010101010111: color_data = Z;
		19'b0100011010101011000: color_data = Z;
		19'b0100011010101011001: color_data = Z;
		19'b0100011010101011010: color_data = Z;
		19'b0100011010101011011: color_data = Z;
		19'b0100011010101011100: color_data = Z;
		19'b0100011010101011101: color_data = Z;
		19'b0100011010101011110: color_data = Z;
		19'b0100011010101011111: color_data = Z;
		19'b0100011010101100000: color_data = Z;
		19'b0100011010101100001: color_data = Z;
		19'b0100011010101100010: color_data = Z;
		19'b0100011010101100011: color_data = Z;
		19'b0100011010101100100: color_data = Z;
		19'b0100011010101100101: color_data = Z;
		19'b0100011010101100110: color_data = Z;
		19'b0100011010101100111: color_data = Z;
		19'b0100011010101101000: color_data = Z;
		19'b0100011010101101001: color_data = Z;
		19'b0100011010101101010: color_data = Z;
		19'b0100011010101101011: color_data = Z;
		19'b0100011010101101100: color_data = Z;
		19'b0100011010101101101: color_data = Z;
		19'b0100011010101101110: color_data = Z;
		19'b0100011010101101111: color_data = Z;
		19'b0100011010101110000: color_data = Z;
		19'b0100011010101110001: color_data = Z;
		19'b0100011010101110010: color_data = Z;
		19'b0100011010101110011: color_data = Z;
		19'b0100011010101110100: color_data = Z;
		19'b0100011010101110101: color_data = Z;
		19'b0100011010101110110: color_data = Z;
		19'b0100011010101110111: color_data = Z;
		19'b0100011010101111000: color_data = Z;
		19'b0100011010101111001: color_data = Z;
		19'b0100011010101111010: color_data = Z;
		19'b0100011010101111011: color_data = Z;
		19'b0100011010101111100: color_data = Z;
		19'b0100011010101111101: color_data = Z;
		19'b0100011010101111110: color_data = Z;
		19'b0100011010101111111: color_data = Z;
		19'b0100011010110000000: color_data = Z;
		19'b0100011010110000001: color_data = Z;
		19'b0100011010110000010: color_data = Z;
		19'b0100011010111001110: color_data = Z;
		19'b0100011010111001111: color_data = Z;
		19'b0100011010111010000: color_data = Z;
		19'b0100011010111010001: color_data = Z;
		19'b0100011010111010010: color_data = Z;
		19'b0100011010111010011: color_data = Z;
		19'b0100011010111010100: color_data = Z;
		19'b0100011010111010101: color_data = Z;
		19'b0100011010111010110: color_data = Z;
		19'b0100011010111010111: color_data = Z;
		19'b0100011010111100000: color_data = Z;
		19'b0100011010111100001: color_data = Z;
		19'b0100011010111100010: color_data = Z;
		19'b0100011100100000101: color_data = Z;
		19'b0100011100100000110: color_data = Z;
		19'b0100011100100000111: color_data = Z;
		19'b0100011100100001000: color_data = Z;
		19'b0100011100100001001: color_data = Z;
		19'b0100011100100001010: color_data = Z;
		19'b0100011100100001011: color_data = Z;
		19'b0100011100100001100: color_data = Z;
		19'b0100011100100001101: color_data = Z;
		19'b0100011100100001110: color_data = Z;
		19'b0100011100100001111: color_data = Z;
		19'b0100011100100010000: color_data = Z;
		19'b0100011100100010001: color_data = Z;
		19'b0100011100100010010: color_data = Z;
		19'b0100011100100010011: color_data = Z;
		19'b0100011100100010100: color_data = Z;
		19'b0100011100100010101: color_data = Z;
		19'b0100011100100010110: color_data = Z;
		19'b0100011100100010111: color_data = Z;
		19'b0100011100100011000: color_data = Z;
		19'b0100011100100011001: color_data = Z;
		19'b0100011100100011010: color_data = Z;
		19'b0100011100100011011: color_data = Z;
		19'b0100011100100011100: color_data = Z;
		19'b0100011100100011101: color_data = Z;
		19'b0100011100100011110: color_data = Z;
		19'b0100011100100011111: color_data = Z;
		19'b0100011100100100000: color_data = Z;
		19'b0100011100100100001: color_data = Z;
		19'b0100011100100100010: color_data = Z;
		19'b0100011100100100011: color_data = Z;
		19'b0100011100100100100: color_data = Z;
		19'b0100011100100100101: color_data = Z;
		19'b0100011100100100110: color_data = Z;
		19'b0100011100100100111: color_data = Z;
		19'b0100011100100101000: color_data = Z;
		19'b0100011100100101001: color_data = Z;
		19'b0100011100100101010: color_data = Z;
		19'b0100011100100101011: color_data = Z;
		19'b0100011100100101100: color_data = Z;
		19'b0100011100100101101: color_data = Z;
		19'b0100011100100101110: color_data = Z;
		19'b0100011100100101111: color_data = Z;
		19'b0100011100100110000: color_data = Z;
		19'b0100011100100110001: color_data = Z;
		19'b0100011100100110010: color_data = Z;
		19'b0100011100100110011: color_data = Z;
		19'b0100011100100110100: color_data = Z;
		19'b0100011100100110101: color_data = Z;
		19'b0100011100100110110: color_data = Z;
		19'b0100011100100110111: color_data = Z;
		19'b0100011100100111000: color_data = Z;
		19'b0100011100100111001: color_data = Z;
		19'b0100011100100111010: color_data = Z;
		19'b0100011100100111011: color_data = Z;
		19'b0100011100100111100: color_data = Z;
		19'b0100011100100111101: color_data = Z;
		19'b0100011100100111110: color_data = Z;
		19'b0100011100100111111: color_data = Z;
		19'b0100011100101000000: color_data = Z;
		19'b0100011100101000001: color_data = Z;
		19'b0100011100101000010: color_data = Z;
		19'b0100011100101000011: color_data = Z;
		19'b0100011100101000100: color_data = Z;
		19'b0100011100101000101: color_data = Z;
		19'b0100011100101000110: color_data = Z;
		19'b0100011100101000111: color_data = Z;
		19'b0100011100101001000: color_data = Z;
		19'b0100011100101001001: color_data = Z;
		19'b0100011100101001010: color_data = Z;
		19'b0100011100101001011: color_data = Z;
		19'b0100011100101001100: color_data = Z;
		19'b0100011100101001101: color_data = Z;
		19'b0100011100101001110: color_data = Z;
		19'b0100011100101001111: color_data = Z;
		19'b0100011100101010000: color_data = Z;
		19'b0100011100101010001: color_data = Z;
		19'b0100011100101010010: color_data = Z;
		19'b0100011100101010011: color_data = Z;
		19'b0100011100101010100: color_data = Z;
		19'b0100011100101010101: color_data = Z;
		19'b0100011100101010110: color_data = Z;
		19'b0100011100101010111: color_data = Z;
		19'b0100011100101011000: color_data = Z;
		19'b0100011100101011001: color_data = Z;
		19'b0100011100101011010: color_data = Z;
		19'b0100011100101011011: color_data = Z;
		19'b0100011100101011100: color_data = Z;
		19'b0100011100101011101: color_data = Z;
		19'b0100011100101011110: color_data = Z;
		19'b0100011100101011111: color_data = Z;
		19'b0100011100101100000: color_data = Z;
		19'b0100011100101100001: color_data = Z;
		19'b0100011100101100010: color_data = Z;
		19'b0100011100101100011: color_data = Z;
		19'b0100011100101100100: color_data = Z;
		19'b0100011100101100101: color_data = Z;
		19'b0100011100101100110: color_data = Z;
		19'b0100011100101100111: color_data = Z;
		19'b0100011100101101000: color_data = Z;
		19'b0100011100101101001: color_data = Z;
		19'b0100011100101101010: color_data = Z;
		19'b0100011100101101011: color_data = Z;
		19'b0100011100101101100: color_data = Z;
		19'b0100011100101101101: color_data = Z;
		19'b0100011100101101110: color_data = Z;
		19'b0100011100101101111: color_data = Z;
		19'b0100011100101110000: color_data = Z;
		19'b0100011100101110001: color_data = Z;
		19'b0100011100101110010: color_data = Z;
		19'b0100011100101110011: color_data = Z;
		19'b0100011100101110100: color_data = Z;
		19'b0100011100101110101: color_data = Z;
		19'b0100011100101110110: color_data = Z;
		19'b0100011100101110111: color_data = Z;
		19'b0100011100101111000: color_data = Z;
		19'b0100011100101111001: color_data = Z;
		19'b0100011100101111010: color_data = Z;
		19'b0100011100101111011: color_data = Z;
		19'b0100011100101111100: color_data = Z;
		19'b0100011100101111101: color_data = Z;
		19'b0100011100101111110: color_data = Z;
		19'b0100011100101111111: color_data = Z;
		19'b0100011100110000000: color_data = Z;
		19'b0100011100110000001: color_data = Z;
		19'b0100011100110000010: color_data = Z;
		19'b0100011100111001110: color_data = Z;
		19'b0100011100111001111: color_data = Z;
		19'b0100011100111010000: color_data = Z;
		19'b0100011100111010001: color_data = Z;
		19'b0100011100111010010: color_data = Z;
		19'b0100011100111010011: color_data = Z;
		19'b0100011100111010100: color_data = Z;
		19'b0100011100111010101: color_data = Z;
		19'b0100011100111010110: color_data = Z;
		19'b0100011100111010111: color_data = Z;
		19'b0100011100111011111: color_data = Z;
		19'b0100011100111100000: color_data = Z;
		19'b0100011100111100001: color_data = Z;
		19'b0100011100111100010: color_data = Z;
		19'b0100011110100000110: color_data = Z;
		19'b0100011110100000111: color_data = Z;
		19'b0100011110100001000: color_data = Z;
		19'b0100011110100001001: color_data = Z;
		19'b0100011110100001010: color_data = Z;
		19'b0100011110100001011: color_data = Z;
		19'b0100011110100001100: color_data = Z;
		19'b0100011110100001101: color_data = Z;
		19'b0100011110100001110: color_data = Z;
		19'b0100011110100001111: color_data = Z;
		19'b0100011110100010000: color_data = Z;
		19'b0100011110100010001: color_data = Z;
		19'b0100011110100010010: color_data = Z;
		19'b0100011110100010011: color_data = Z;
		19'b0100011110100010100: color_data = Z;
		19'b0100011110100010101: color_data = Z;
		19'b0100011110100010110: color_data = Z;
		19'b0100011110100010111: color_data = Z;
		19'b0100011110100011000: color_data = Z;
		19'b0100011110100011001: color_data = Z;
		19'b0100011110100011010: color_data = Z;
		19'b0100011110100011011: color_data = Z;
		19'b0100011110100011100: color_data = Z;
		19'b0100011110100011101: color_data = Z;
		19'b0100011110100011110: color_data = Z;
		19'b0100011110100011111: color_data = Z;
		19'b0100011110100100000: color_data = Z;
		19'b0100011110100100001: color_data = Z;
		19'b0100011110100100010: color_data = Z;
		19'b0100011110100100011: color_data = Z;
		19'b0100011110100100100: color_data = Z;
		19'b0100011110100100101: color_data = Z;
		19'b0100011110100100110: color_data = Z;
		19'b0100011110100100111: color_data = Z;
		19'b0100011110100101000: color_data = Z;
		19'b0100011110100101001: color_data = Z;
		19'b0100011110100101010: color_data = Z;
		19'b0100011110100101011: color_data = Z;
		19'b0100011110100101100: color_data = Z;
		19'b0100011110100101101: color_data = Z;
		19'b0100011110100101110: color_data = Z;
		19'b0100011110100101111: color_data = Z;
		19'b0100011110100110000: color_data = Z;
		19'b0100011110100110001: color_data = Z;
		19'b0100011110100110010: color_data = Z;
		19'b0100011110100110011: color_data = Z;
		19'b0100011110100110100: color_data = Z;
		19'b0100011110100110101: color_data = Z;
		19'b0100011110100110110: color_data = Z;
		19'b0100011110100110111: color_data = Z;
		19'b0100011110100111000: color_data = Z;
		19'b0100011110100111001: color_data = Z;
		19'b0100011110100111010: color_data = Z;
		19'b0100011110100111011: color_data = Z;
		19'b0100011110100111100: color_data = Z;
		19'b0100011110100111101: color_data = Z;
		19'b0100011110100111110: color_data = Z;
		19'b0100011110100111111: color_data = Z;
		19'b0100011110101000000: color_data = Z;
		19'b0100011110101000001: color_data = Z;
		19'b0100011110101000010: color_data = Z;
		19'b0100011110101000011: color_data = Z;
		19'b0100011110101000100: color_data = Z;
		19'b0100011110101000101: color_data = Z;
		19'b0100011110101000110: color_data = Z;
		19'b0100011110101000111: color_data = Z;
		19'b0100011110101001000: color_data = Z;
		19'b0100011110101001001: color_data = Z;
		19'b0100011110101001010: color_data = Z;
		19'b0100011110101001011: color_data = Z;
		19'b0100011110101001100: color_data = Z;
		19'b0100011110101001101: color_data = Z;
		19'b0100011110101001110: color_data = Z;
		19'b0100011110101001111: color_data = Z;
		19'b0100011110101010000: color_data = Z;
		19'b0100011110101010001: color_data = Z;
		19'b0100011110101010010: color_data = Z;
		19'b0100011110101010011: color_data = Z;
		19'b0100011110101010100: color_data = Z;
		19'b0100011110101010101: color_data = Z;
		19'b0100011110101010110: color_data = Z;
		19'b0100011110101010111: color_data = Z;
		19'b0100011110101011000: color_data = Z;
		19'b0100011110101011001: color_data = Z;
		19'b0100011110101011010: color_data = Z;
		19'b0100011110101011011: color_data = Z;
		19'b0100011110101011100: color_data = Z;
		19'b0100011110101011101: color_data = Z;
		19'b0100011110101011110: color_data = Z;
		19'b0100011110101011111: color_data = Z;
		19'b0100011110101100000: color_data = Z;
		19'b0100011110101100001: color_data = Z;
		19'b0100011110101100010: color_data = Z;
		19'b0100011110101100011: color_data = Z;
		19'b0100011110101100100: color_data = Z;
		19'b0100011110101100101: color_data = Z;
		19'b0100011110101100110: color_data = Z;
		19'b0100011110101100111: color_data = Z;
		19'b0100011110101101000: color_data = Z;
		19'b0100011110101101001: color_data = Z;
		19'b0100011110101101010: color_data = Z;
		19'b0100011110101101011: color_data = Z;
		19'b0100011110101101100: color_data = Z;
		19'b0100011110101101101: color_data = Z;
		19'b0100011110101101110: color_data = Z;
		19'b0100011110101101111: color_data = Z;
		19'b0100011110101110000: color_data = Z;
		19'b0100011110101110001: color_data = Z;
		19'b0100011110101110010: color_data = Z;
		19'b0100011110101110011: color_data = Z;
		19'b0100011110101110100: color_data = Z;
		19'b0100011110101110101: color_data = Z;
		19'b0100011110101110110: color_data = Z;
		19'b0100011110101110111: color_data = Z;
		19'b0100011110101111000: color_data = Z;
		19'b0100011110101111001: color_data = Z;
		19'b0100011110101111010: color_data = Z;
		19'b0100011110101111011: color_data = Z;
		19'b0100011110101111100: color_data = Z;
		19'b0100011110101111101: color_data = Z;
		19'b0100011110101111110: color_data = Z;
		19'b0100011110101111111: color_data = Z;
		19'b0100011110110000000: color_data = Z;
		19'b0100011110110000001: color_data = Z;
		19'b0100011110111001110: color_data = Z;
		19'b0100011110111001111: color_data = Z;
		19'b0100011110111010000: color_data = Z;
		19'b0100011110111010001: color_data = Z;
		19'b0100011110111010010: color_data = Z;
		19'b0100011110111010011: color_data = Z;
		19'b0100011110111010100: color_data = Z;
		19'b0100011110111010101: color_data = Z;
		19'b0100011110111010110: color_data = Z;
		19'b0100011110111011111: color_data = Z;
		19'b0100011110111100000: color_data = Z;
		19'b0100011110111100010: color_data = Z;
		19'b0100100000100000110: color_data = Z;
		19'b0100100000100000111: color_data = Z;
		19'b0100100000100001000: color_data = Z;
		19'b0100100000100001101: color_data = Z;
		19'b0100100000100001110: color_data = Z;
		19'b0100100000100001111: color_data = Z;
		19'b0100100000100010000: color_data = Z;
		19'b0100100000100010001: color_data = Z;
		19'b0100100000100010010: color_data = Z;
		19'b0100100000100010011: color_data = Z;
		19'b0100100000100010100: color_data = Z;
		19'b0100100000100010101: color_data = Z;
		19'b0100100000100010110: color_data = Z;
		19'b0100100000100010111: color_data = Z;
		19'b0100100000100011000: color_data = Z;
		19'b0100100000100011001: color_data = Z;
		19'b0100100000100011010: color_data = Z;
		19'b0100100000100011011: color_data = Z;
		19'b0100100000100011100: color_data = Z;
		19'b0100100000100011101: color_data = Z;
		19'b0100100000100011110: color_data = Z;
		19'b0100100000100011111: color_data = Z;
		19'b0100100000100100000: color_data = Z;
		19'b0100100000100100001: color_data = Z;
		19'b0100100000100100010: color_data = Z;
		19'b0100100000100100011: color_data = Z;
		19'b0100100000100100100: color_data = Z;
		19'b0100100000100100101: color_data = Z;
		19'b0100100000100100110: color_data = Z;
		19'b0100100000100100111: color_data = Z;
		19'b0100100000100101000: color_data = Z;
		19'b0100100000100101001: color_data = Z;
		19'b0100100000100101010: color_data = Z;
		19'b0100100000100101011: color_data = Z;
		19'b0100100000100101100: color_data = Z;
		19'b0100100000100101101: color_data = Z;
		19'b0100100000100101110: color_data = Z;
		19'b0100100000100101111: color_data = Z;
		19'b0100100000100110000: color_data = Z;
		19'b0100100000100110001: color_data = Z;
		19'b0100100000100110010: color_data = Z;
		19'b0100100000100110011: color_data = Z;
		19'b0100100000100110100: color_data = Z;
		19'b0100100000100110101: color_data = Z;
		19'b0100100000100110110: color_data = Z;
		19'b0100100000100110111: color_data = Z;
		19'b0100100000100111000: color_data = Z;
		19'b0100100000100111001: color_data = Z;
		19'b0100100000100111010: color_data = Z;
		19'b0100100000100111011: color_data = Z;
		19'b0100100000100111100: color_data = Z;
		19'b0100100000100111101: color_data = Z;
		19'b0100100000100111110: color_data = Z;
		19'b0100100000100111111: color_data = Z;
		19'b0100100000101000000: color_data = Z;
		19'b0100100000101000001: color_data = Z;
		19'b0100100000101000010: color_data = Z;
		19'b0100100000101000011: color_data = Z;
		19'b0100100000101000100: color_data = Z;
		19'b0100100000101000101: color_data = Z;
		19'b0100100000101000110: color_data = Z;
		19'b0100100000101000111: color_data = Z;
		19'b0100100000101001000: color_data = Z;
		19'b0100100000101001001: color_data = Z;
		19'b0100100000101001010: color_data = Z;
		19'b0100100000101001011: color_data = Z;
		19'b0100100000101001100: color_data = Z;
		19'b0100100000101001101: color_data = Z;
		19'b0100100000101001110: color_data = Z;
		19'b0100100000101001111: color_data = Z;
		19'b0100100000101010000: color_data = Z;
		19'b0100100000101010001: color_data = Z;
		19'b0100100000101010010: color_data = Z;
		19'b0100100000101010011: color_data = Z;
		19'b0100100000101010100: color_data = Z;
		19'b0100100000101010101: color_data = Z;
		19'b0100100000101010110: color_data = Z;
		19'b0100100000101010111: color_data = Z;
		19'b0100100000101011000: color_data = Z;
		19'b0100100000101011001: color_data = Z;
		19'b0100100000101011010: color_data = Z;
		19'b0100100000101011011: color_data = Z;
		19'b0100100000101011100: color_data = Z;
		19'b0100100000101011101: color_data = Z;
		19'b0100100000101011110: color_data = Z;
		19'b0100100000101011111: color_data = Z;
		19'b0100100000101100000: color_data = Z;
		19'b0100100000101100001: color_data = Z;
		19'b0100100000101100010: color_data = Z;
		19'b0100100000101100011: color_data = Z;
		19'b0100100000101100100: color_data = Z;
		19'b0100100000101100101: color_data = Z;
		19'b0100100000101100110: color_data = Z;
		19'b0100100000101100111: color_data = Z;
		19'b0100100000101101000: color_data = Z;
		19'b0100100000101101001: color_data = Z;
		19'b0100100000101101010: color_data = Z;
		19'b0100100000101101011: color_data = Z;
		19'b0100100000101101100: color_data = Z;
		19'b0100100000101101101: color_data = Z;
		19'b0100100000101101110: color_data = Z;
		19'b0100100000101101111: color_data = Z;
		19'b0100100000101110000: color_data = Z;
		19'b0100100000101110001: color_data = Z;
		19'b0100100000101110010: color_data = Z;
		19'b0100100000101110011: color_data = Z;
		19'b0100100000101110100: color_data = Z;
		19'b0100100000101110101: color_data = Z;
		19'b0100100000101110110: color_data = Z;
		19'b0100100000101110111: color_data = Z;
		19'b0100100000101111000: color_data = Z;
		19'b0100100000101111001: color_data = Z;
		19'b0100100000101111010: color_data = Z;
		19'b0100100000101111011: color_data = Z;
		19'b0100100000101111100: color_data = Z;
		19'b0100100000101111101: color_data = Z;
		19'b0100100000101111110: color_data = Z;
		19'b0100100000101111111: color_data = Z;
		19'b0100100000110000000: color_data = Z;
		19'b0100100000110000001: color_data = Z;
		19'b0100100000111001110: color_data = Z;
		19'b0100100000111001111: color_data = Z;
		19'b0100100000111010000: color_data = Z;
		19'b0100100000111010001: color_data = Z;
		19'b0100100000111010010: color_data = Z;
		19'b0100100000111010011: color_data = Z;
		19'b0100100000111010100: color_data = Z;
		19'b0100100000111010101: color_data = Z;
		19'b0100100000111010110: color_data = Z;
		19'b0100100000111010111: color_data = Z;
		19'b0100100000111100000: color_data = Z;
		19'b0100100000111100001: color_data = Z;
		19'b0100100000111100010: color_data = Z;
		19'b0100100010100001111: color_data = Z;
		19'b0100100010100010000: color_data = Z;
		19'b0100100010100010001: color_data = Z;
		19'b0100100010100010010: color_data = Z;
		19'b0100100010100010011: color_data = Z;
		19'b0100100010100010100: color_data = Z;
		19'b0100100010100010101: color_data = Z;
		19'b0100100010100010110: color_data = Z;
		19'b0100100010100010111: color_data = Z;
		19'b0100100010100011000: color_data = Z;
		19'b0100100010100011001: color_data = Z;
		19'b0100100010100011010: color_data = Z;
		19'b0100100010100011011: color_data = Z;
		19'b0100100010100011100: color_data = Z;
		19'b0100100010100011101: color_data = Z;
		19'b0100100010100011110: color_data = Z;
		19'b0100100010100011111: color_data = Z;
		19'b0100100010100100000: color_data = Z;
		19'b0100100010100100001: color_data = Z;
		19'b0100100010100100010: color_data = Z;
		19'b0100100010100100011: color_data = Z;
		19'b0100100010100100100: color_data = Z;
		19'b0100100010100100101: color_data = Z;
		19'b0100100010100100110: color_data = Z;
		19'b0100100010100100111: color_data = Z;
		19'b0100100010100101000: color_data = Z;
		19'b0100100010100101001: color_data = Z;
		19'b0100100010100101010: color_data = Z;
		19'b0100100010100101011: color_data = Z;
		19'b0100100010100101100: color_data = Z;
		19'b0100100010100101101: color_data = Z;
		19'b0100100010100101110: color_data = Z;
		19'b0100100010100101111: color_data = Z;
		19'b0100100010100110000: color_data = Z;
		19'b0100100010100110001: color_data = Z;
		19'b0100100010100110010: color_data = Z;
		19'b0100100010100110011: color_data = Z;
		19'b0100100010100110100: color_data = Z;
		19'b0100100010100110101: color_data = Z;
		19'b0100100010100110110: color_data = Z;
		19'b0100100010100110111: color_data = Z;
		19'b0100100010100111000: color_data = Z;
		19'b0100100010100111001: color_data = Z;
		19'b0100100010100111010: color_data = Z;
		19'b0100100010100111011: color_data = Z;
		19'b0100100010100111100: color_data = Z;
		19'b0100100010100111101: color_data = Z;
		19'b0100100010100111110: color_data = Z;
		19'b0100100010100111111: color_data = Z;
		19'b0100100010101000000: color_data = Z;
		19'b0100100010101000001: color_data = Z;
		19'b0100100010101000010: color_data = Z;
		19'b0100100010101000011: color_data = Z;
		19'b0100100010101000100: color_data = Z;
		19'b0100100010101000101: color_data = Z;
		19'b0100100010101000110: color_data = Z;
		19'b0100100010101000111: color_data = Z;
		19'b0100100010101001000: color_data = Z;
		19'b0100100010101001001: color_data = Z;
		19'b0100100010101001010: color_data = Z;
		19'b0100100010101001011: color_data = Z;
		19'b0100100010101001100: color_data = Z;
		19'b0100100010101001101: color_data = Z;
		19'b0100100010101001110: color_data = Z;
		19'b0100100010101001111: color_data = Z;
		19'b0100100010101010000: color_data = Z;
		19'b0100100010101010001: color_data = Z;
		19'b0100100010101010010: color_data = Z;
		19'b0100100010101010011: color_data = Z;
		19'b0100100010101010100: color_data = Z;
		19'b0100100010101010101: color_data = Z;
		19'b0100100010101010110: color_data = Z;
		19'b0100100010101010111: color_data = Z;
		19'b0100100010101011000: color_data = Z;
		19'b0100100010101011001: color_data = Z;
		19'b0100100010101011010: color_data = Z;
		19'b0100100010101011011: color_data = Z;
		19'b0100100010101011100: color_data = Z;
		19'b0100100010101011101: color_data = Z;
		19'b0100100010101011110: color_data = Z;
		19'b0100100010101011111: color_data = Z;
		19'b0100100010101100000: color_data = Z;
		19'b0100100010101100001: color_data = Z;
		19'b0100100010101100010: color_data = Z;
		19'b0100100010101100011: color_data = Z;
		19'b0100100010101100100: color_data = Z;
		19'b0100100010101100101: color_data = Z;
		19'b0100100010101100110: color_data = Z;
		19'b0100100010101100111: color_data = Z;
		19'b0100100010101101000: color_data = Z;
		19'b0100100010101101001: color_data = Z;
		19'b0100100010101101010: color_data = Z;
		19'b0100100010101101011: color_data = Z;
		19'b0100100010101101100: color_data = Z;
		19'b0100100010101101101: color_data = Z;
		19'b0100100010101101110: color_data = Z;
		19'b0100100010101101111: color_data = Z;
		19'b0100100010101110000: color_data = Z;
		19'b0100100010101110001: color_data = Z;
		19'b0100100010101110010: color_data = Z;
		19'b0100100010101110011: color_data = Z;
		19'b0100100010101110100: color_data = Z;
		19'b0100100010101110101: color_data = Z;
		19'b0100100010101110110: color_data = Z;
		19'b0100100010101110111: color_data = Z;
		19'b0100100010101111000: color_data = Z;
		19'b0100100010101111001: color_data = Z;
		19'b0100100010101111010: color_data = Z;
		19'b0100100010101111011: color_data = Z;
		19'b0100100010101111100: color_data = Z;
		19'b0100100010101111101: color_data = Z;
		19'b0100100010101111110: color_data = Z;
		19'b0100100010101111111: color_data = Z;
		19'b0100100010110000000: color_data = Z;
		19'b0100100010110000001: color_data = Z;
		19'b0100100010111001110: color_data = Z;
		19'b0100100010111001111: color_data = Z;
		19'b0100100010111010000: color_data = Z;
		19'b0100100010111010001: color_data = Z;
		19'b0100100010111010010: color_data = Z;
		19'b0100100010111010011: color_data = Z;
		19'b0100100010111010100: color_data = Z;
		19'b0100100010111010101: color_data = Z;
		19'b0100100010111010110: color_data = Z;
		19'b0100100010111010111: color_data = Z;
		19'b0100100010111100000: color_data = Z;
		19'b0100100010111100001: color_data = Z;
		19'b0100100010111100010: color_data = Z;
		19'b0100100100100010001: color_data = Z;
		19'b0100100100100010010: color_data = Z;
		19'b0100100100100010011: color_data = Z;
		19'b0100100100100010100: color_data = Z;
		19'b0100100100100010101: color_data = Z;
		19'b0100100100100010110: color_data = Z;
		19'b0100100100100010111: color_data = Z;
		19'b0100100100100011000: color_data = Z;
		19'b0100100100100011001: color_data = Z;
		19'b0100100100100011010: color_data = Z;
		19'b0100100100100011011: color_data = Z;
		19'b0100100100100011100: color_data = Z;
		19'b0100100100100011101: color_data = Z;
		19'b0100100100100011110: color_data = Z;
		19'b0100100100100011111: color_data = Z;
		19'b0100100100100100000: color_data = Z;
		19'b0100100100100100001: color_data = Z;
		19'b0100100100100100010: color_data = Z;
		19'b0100100100100100011: color_data = Z;
		19'b0100100100100100100: color_data = Z;
		19'b0100100100100100101: color_data = Z;
		19'b0100100100100100110: color_data = Z;
		19'b0100100100100100111: color_data = Z;
		19'b0100100100100101000: color_data = Z;
		19'b0100100100100101001: color_data = Z;
		19'b0100100100100101010: color_data = Z;
		19'b0100100100100101011: color_data = Z;
		19'b0100100100100101100: color_data = Z;
		19'b0100100100100101101: color_data = Z;
		19'b0100100100100101110: color_data = Z;
		19'b0100100100100101111: color_data = Z;
		19'b0100100100100110000: color_data = Z;
		19'b0100100100100110001: color_data = Z;
		19'b0100100100100110010: color_data = Z;
		19'b0100100100100110011: color_data = Z;
		19'b0100100100100110100: color_data = Z;
		19'b0100100100100110101: color_data = Z;
		19'b0100100100100110110: color_data = Z;
		19'b0100100100100110111: color_data = Z;
		19'b0100100100100111000: color_data = Z;
		19'b0100100100100111001: color_data = Z;
		19'b0100100100100111010: color_data = Z;
		19'b0100100100100111011: color_data = Z;
		19'b0100100100100111100: color_data = Z;
		19'b0100100100100111101: color_data = Z;
		19'b0100100100100111110: color_data = Z;
		19'b0100100100100111111: color_data = Z;
		19'b0100100100101000000: color_data = Z;
		19'b0100100100101000001: color_data = Z;
		19'b0100100100101000010: color_data = Z;
		19'b0100100100101000011: color_data = Z;
		19'b0100100100101000100: color_data = Z;
		19'b0100100100101000101: color_data = Z;
		19'b0100100100101000110: color_data = Z;
		19'b0100100100101000111: color_data = Z;
		19'b0100100100101001000: color_data = Z;
		19'b0100100100101001001: color_data = Z;
		19'b0100100100101001010: color_data = Z;
		19'b0100100100101001011: color_data = Z;
		19'b0100100100101001100: color_data = Z;
		19'b0100100100101001101: color_data = Z;
		19'b0100100100101001110: color_data = Z;
		19'b0100100100101001111: color_data = Z;
		19'b0100100100101010000: color_data = Z;
		19'b0100100100101010001: color_data = Z;
		19'b0100100100101010010: color_data = Z;
		19'b0100100100101010011: color_data = Z;
		19'b0100100100101010100: color_data = Z;
		19'b0100100100101010101: color_data = Z;
		19'b0100100100101010110: color_data = Z;
		19'b0100100100101010111: color_data = Z;
		19'b0100100100101011000: color_data = Z;
		19'b0100100100101011001: color_data = Z;
		19'b0100100100101011010: color_data = Z;
		19'b0100100100101011011: color_data = Z;
		19'b0100100100101011100: color_data = Z;
		19'b0100100100101011101: color_data = Z;
		19'b0100100100101011110: color_data = Z;
		19'b0100100100101011111: color_data = Z;
		19'b0100100100101100000: color_data = Z;
		19'b0100100100101100001: color_data = Z;
		19'b0100100100101100010: color_data = Z;
		19'b0100100100101100011: color_data = Z;
		19'b0100100100101100100: color_data = Z;
		19'b0100100100101100101: color_data = Z;
		19'b0100100100101100110: color_data = Z;
		19'b0100100100101100111: color_data = Z;
		19'b0100100100101101000: color_data = Z;
		19'b0100100100101101001: color_data = Z;
		19'b0100100100101101010: color_data = Z;
		19'b0100100100101101011: color_data = Z;
		19'b0100100100101101100: color_data = Z;
		19'b0100100100101101101: color_data = Z;
		19'b0100100100101101110: color_data = Z;
		19'b0100100100101101111: color_data = Z;
		19'b0100100100101110000: color_data = Z;
		19'b0100100100101110001: color_data = Z;
		19'b0100100100101110010: color_data = Z;
		19'b0100100100101110011: color_data = Z;
		19'b0100100100101110100: color_data = Z;
		19'b0100100100101110101: color_data = Z;
		19'b0100100100101110110: color_data = Z;
		19'b0100100100101110111: color_data = Z;
		19'b0100100100101111000: color_data = Z;
		19'b0100100100101111001: color_data = Z;
		19'b0100100100101111010: color_data = Z;
		19'b0100100100101111011: color_data = Z;
		19'b0100100100101111100: color_data = Z;
		19'b0100100100101111101: color_data = Z;
		19'b0100100100101111110: color_data = Z;
		19'b0100100100101111111: color_data = Z;
		19'b0100100100110000000: color_data = Z;
		19'b0100100100110000001: color_data = Z;
		19'b0100100100111001110: color_data = Z;
		19'b0100100100111001111: color_data = Z;
		19'b0100100100111010000: color_data = Z;
		19'b0100100100111010001: color_data = Z;
		19'b0100100100111010010: color_data = Z;
		19'b0100100100111010011: color_data = Z;
		19'b0100100100111010100: color_data = Z;
		19'b0100100100111010101: color_data = Z;
		19'b0100100100111010110: color_data = Z;
		19'b0100100100111010111: color_data = Z;
		19'b0100100100111100000: color_data = Z;
		19'b0100100100111100001: color_data = Z;
		19'b0100100100111100010: color_data = Z;
		19'b0100100110100010010: color_data = Z;
		19'b0100100110100010011: color_data = Z;
		19'b0100100110100010100: color_data = Z;
		19'b0100100110100010101: color_data = Z;
		19'b0100100110100010110: color_data = Z;
		19'b0100100110100010111: color_data = Z;
		19'b0100100110100011000: color_data = Z;
		19'b0100100110100011001: color_data = Z;
		19'b0100100110100011010: color_data = Z;
		19'b0100100110100011011: color_data = Z;
		19'b0100100110100011100: color_data = Z;
		19'b0100100110100011101: color_data = Z;
		19'b0100100110100011110: color_data = Z;
		19'b0100100110100011111: color_data = Z;
		19'b0100100110100100000: color_data = Z;
		19'b0100100110100100001: color_data = Z;
		19'b0100100110100100010: color_data = Z;
		19'b0100100110100100011: color_data = Z;
		19'b0100100110100100100: color_data = Z;
		19'b0100100110100100101: color_data = Z;
		19'b0100100110100100110: color_data = Z;
		19'b0100100110100100111: color_data = Z;
		19'b0100100110100101000: color_data = Z;
		19'b0100100110100101001: color_data = Z;
		19'b0100100110100101010: color_data = Z;
		19'b0100100110100101011: color_data = Z;
		19'b0100100110100101100: color_data = Z;
		19'b0100100110100101101: color_data = Z;
		19'b0100100110100101110: color_data = Z;
		19'b0100100110100101111: color_data = Z;
		19'b0100100110100110000: color_data = Z;
		19'b0100100110100110001: color_data = Z;
		19'b0100100110100110010: color_data = Z;
		19'b0100100110100110011: color_data = Z;
		19'b0100100110100110100: color_data = Z;
		19'b0100100110100110101: color_data = Z;
		19'b0100100110100110110: color_data = Z;
		19'b0100100110100110111: color_data = Z;
		19'b0100100110100111000: color_data = Z;
		19'b0100100110100111001: color_data = Z;
		19'b0100100110100111010: color_data = Z;
		19'b0100100110100111011: color_data = Z;
		19'b0100100110100111100: color_data = Z;
		19'b0100100110100111101: color_data = Z;
		19'b0100100110100111110: color_data = Z;
		19'b0100100110100111111: color_data = Z;
		19'b0100100110101000000: color_data = Z;
		19'b0100100110101000001: color_data = Z;
		19'b0100100110101000010: color_data = Z;
		19'b0100100110101000011: color_data = Z;
		19'b0100100110101000100: color_data = Z;
		19'b0100100110101000101: color_data = Z;
		19'b0100100110101000110: color_data = Z;
		19'b0100100110101000111: color_data = Z;
		19'b0100100110101001000: color_data = Z;
		19'b0100100110101001001: color_data = Z;
		19'b0100100110101001010: color_data = Z;
		19'b0100100110101001011: color_data = Z;
		19'b0100100110101001100: color_data = Z;
		19'b0100100110101001101: color_data = Z;
		19'b0100100110101001110: color_data = Z;
		19'b0100100110101001111: color_data = Z;
		19'b0100100110101010000: color_data = Z;
		19'b0100100110101010001: color_data = Z;
		19'b0100100110101010010: color_data = Z;
		19'b0100100110101010011: color_data = Z;
		19'b0100100110101010100: color_data = Z;
		19'b0100100110101010101: color_data = Z;
		19'b0100100110101010110: color_data = Z;
		19'b0100100110101010111: color_data = Z;
		19'b0100100110101011000: color_data = Z;
		19'b0100100110101011001: color_data = Z;
		19'b0100100110101011010: color_data = Z;
		19'b0100100110101011011: color_data = Z;
		19'b0100100110101011100: color_data = Z;
		19'b0100100110101011101: color_data = Z;
		19'b0100100110101011110: color_data = Z;
		19'b0100100110101011111: color_data = Z;
		19'b0100100110101100000: color_data = Z;
		19'b0100100110101100001: color_data = Z;
		19'b0100100110101100010: color_data = Z;
		19'b0100100110101100011: color_data = Z;
		19'b0100100110101100100: color_data = Z;
		19'b0100100110101100101: color_data = Z;
		19'b0100100110101100110: color_data = Z;
		19'b0100100110101100111: color_data = Z;
		19'b0100100110101101000: color_data = Z;
		19'b0100100110101101001: color_data = Z;
		19'b0100100110101101010: color_data = Z;
		19'b0100100110101101011: color_data = Z;
		19'b0100100110101101100: color_data = Z;
		19'b0100100110101101101: color_data = Z;
		19'b0100100110101101110: color_data = Z;
		19'b0100100110101101111: color_data = Z;
		19'b0100100110101110000: color_data = Z;
		19'b0100100110101110001: color_data = Z;
		19'b0100100110101110010: color_data = Z;
		19'b0100100110101110011: color_data = Z;
		19'b0100100110101110100: color_data = Z;
		19'b0100100110101110101: color_data = Z;
		19'b0100100110101110110: color_data = Z;
		19'b0100100110101110111: color_data = Z;
		19'b0100100110101111000: color_data = Z;
		19'b0100100110101111001: color_data = Z;
		19'b0100100110101111010: color_data = Z;
		19'b0100100110101111011: color_data = Z;
		19'b0100100110101111100: color_data = Z;
		19'b0100100110101111101: color_data = Z;
		19'b0100100110101111110: color_data = Z;
		19'b0100100110101111111: color_data = Z;
		19'b0100100110110000000: color_data = Z;
		19'b0100100110110000001: color_data = Z;
		19'b0100100110111001110: color_data = Z;
		19'b0100100110111001111: color_data = Z;
		19'b0100100110111010000: color_data = Z;
		19'b0100100110111010001: color_data = Z;
		19'b0100100110111010010: color_data = Z;
		19'b0100100110111010011: color_data = Z;
		19'b0100100110111010100: color_data = Z;
		19'b0100100110111010101: color_data = Z;
		19'b0100100110111010110: color_data = Z;
		19'b0100100110111010111: color_data = Z;
		19'b0100100110111100000: color_data = Z;
		19'b0100100110111100001: color_data = Z;
		19'b0100100110111100010: color_data = Z;
		19'b0100101000100010010: color_data = Z;
		19'b0100101000100010101: color_data = Z;
		19'b0100101000100010110: color_data = Z;
		19'b0100101000100010111: color_data = Z;
		19'b0100101000100011000: color_data = Z;
		19'b0100101000100011001: color_data = Z;
		19'b0100101000100011010: color_data = Z;
		19'b0100101000100011011: color_data = Z;
		19'b0100101000100011100: color_data = Z;
		19'b0100101000100011101: color_data = Z;
		19'b0100101000100011110: color_data = Z;
		19'b0100101000100011111: color_data = Z;
		19'b0100101000100100000: color_data = Z;
		19'b0100101000100100001: color_data = Z;
		19'b0100101000100100010: color_data = Z;
		19'b0100101000100100011: color_data = Z;
		19'b0100101000100100100: color_data = Z;
		19'b0100101000100100101: color_data = Z;
		19'b0100101000100100110: color_data = Z;
		19'b0100101000100100111: color_data = Z;
		19'b0100101000100101000: color_data = Z;
		19'b0100101000100101001: color_data = Z;
		19'b0100101000100101010: color_data = Z;
		19'b0100101000100101011: color_data = Z;
		19'b0100101000100101100: color_data = Z;
		19'b0100101000100101101: color_data = Z;
		19'b0100101000100101110: color_data = Z;
		19'b0100101000100101111: color_data = Z;
		19'b0100101000100110000: color_data = Z;
		19'b0100101000100110001: color_data = Z;
		19'b0100101000100110010: color_data = Z;
		19'b0100101000100110011: color_data = Z;
		19'b0100101000100110100: color_data = Z;
		19'b0100101000100110101: color_data = Z;
		19'b0100101000100110110: color_data = Z;
		19'b0100101000100110111: color_data = Z;
		19'b0100101000100111000: color_data = Z;
		19'b0100101000100111001: color_data = Z;
		19'b0100101000100111010: color_data = Z;
		19'b0100101000100111011: color_data = Z;
		19'b0100101000100111100: color_data = Z;
		19'b0100101000100111101: color_data = Z;
		19'b0100101000100111110: color_data = Z;
		19'b0100101000100111111: color_data = Z;
		19'b0100101000101000000: color_data = Z;
		19'b0100101000101000001: color_data = Z;
		19'b0100101000101000010: color_data = Z;
		19'b0100101000101000011: color_data = Z;
		19'b0100101000101000100: color_data = Z;
		19'b0100101000101000101: color_data = Z;
		19'b0100101000101000110: color_data = Z;
		19'b0100101000101000111: color_data = Z;
		19'b0100101000101001000: color_data = Z;
		19'b0100101000101001001: color_data = Z;
		19'b0100101000101001010: color_data = Z;
		19'b0100101000101001011: color_data = Z;
		19'b0100101000101001100: color_data = Z;
		19'b0100101000101001101: color_data = Z;
		19'b0100101000101001110: color_data = Z;
		19'b0100101000101001111: color_data = Z;
		19'b0100101000101010000: color_data = Z;
		19'b0100101000101010001: color_data = Z;
		19'b0100101000101010010: color_data = Z;
		19'b0100101000101010011: color_data = Z;
		19'b0100101000101010100: color_data = Z;
		19'b0100101000101010101: color_data = Z;
		19'b0100101000101010110: color_data = Z;
		19'b0100101000101010111: color_data = Z;
		19'b0100101000101011000: color_data = Z;
		19'b0100101000101011001: color_data = Z;
		19'b0100101000101011010: color_data = Z;
		19'b0100101000101011011: color_data = Z;
		19'b0100101000101011100: color_data = Z;
		19'b0100101000101011101: color_data = Z;
		19'b0100101000101011110: color_data = Z;
		19'b0100101000101011111: color_data = Z;
		19'b0100101000101100000: color_data = Z;
		19'b0100101000101100001: color_data = Z;
		19'b0100101000101100010: color_data = Z;
		19'b0100101000101100011: color_data = Z;
		19'b0100101000101100100: color_data = Z;
		19'b0100101000101100101: color_data = Z;
		19'b0100101000101100110: color_data = Z;
		19'b0100101000101100111: color_data = Z;
		19'b0100101000101101000: color_data = Z;
		19'b0100101000101101001: color_data = Z;
		19'b0100101000101101010: color_data = Z;
		19'b0100101000101101011: color_data = Z;
		19'b0100101000101101100: color_data = Z;
		19'b0100101000101101101: color_data = Z;
		19'b0100101000101101110: color_data = Z;
		19'b0100101000101101111: color_data = Z;
		19'b0100101000101110000: color_data = Z;
		19'b0100101000101110001: color_data = Z;
		19'b0100101000101110010: color_data = Z;
		19'b0100101000101110011: color_data = Z;
		19'b0100101000101110100: color_data = Z;
		19'b0100101000101110101: color_data = Z;
		19'b0100101000101110110: color_data = Z;
		19'b0100101000101110111: color_data = Z;
		19'b0100101000101111000: color_data = Z;
		19'b0100101000101111001: color_data = Z;
		19'b0100101000101111010: color_data = Z;
		19'b0100101000101111011: color_data = Z;
		19'b0100101000101111100: color_data = Z;
		19'b0100101000101111101: color_data = Z;
		19'b0100101000101111110: color_data = Z;
		19'b0100101000101111111: color_data = Z;
		19'b0100101000110000000: color_data = Z;
		19'b0100101000111001110: color_data = Z;
		19'b0100101000111001111: color_data = Z;
		19'b0100101000111010000: color_data = Z;
		19'b0100101000111010001: color_data = Z;
		19'b0100101000111010010: color_data = Z;
		19'b0100101000111010011: color_data = Z;
		19'b0100101000111010100: color_data = Z;
		19'b0100101000111010101: color_data = Z;
		19'b0100101000111010110: color_data = Z;
		19'b0100101000111010111: color_data = Z;
		19'b0100101000111011000: color_data = Z;
		19'b0100101000111011001: color_data = Z;
		19'b0100101000111011010: color_data = Z;
		19'b0100101000111011011: color_data = Z;
		19'b0100101000111100001: color_data = Z;
		19'b0100101000111100010: color_data = Z;
		19'b0100101010100001111: color_data = Z;
		19'b0100101010100010000: color_data = Z;
		19'b0100101010100010001: color_data = Z;
		19'b0100101010100010010: color_data = Z;
		19'b0100101010100010011: color_data = Z;
		19'b0100101010100010100: color_data = Z;
		19'b0100101010100010101: color_data = Z;
		19'b0100101010100010110: color_data = Z;
		19'b0100101010100010111: color_data = Z;
		19'b0100101010100011000: color_data = Z;
		19'b0100101010100011001: color_data = Z;
		19'b0100101010100011010: color_data = Z;
		19'b0100101010100011011: color_data = Z;
		19'b0100101010100011100: color_data = Z;
		19'b0100101010100011101: color_data = Z;
		19'b0100101010100100001: color_data = Z;
		19'b0100101010100100010: color_data = Z;
		19'b0100101010100100011: color_data = Z;
		19'b0100101010100100100: color_data = Z;
		19'b0100101010100100101: color_data = Z;
		19'b0100101010100100110: color_data = Z;
		19'b0100101010100100111: color_data = Z;
		19'b0100101010100101000: color_data = Z;
		19'b0100101010100101001: color_data = Z;
		19'b0100101010100101010: color_data = Z;
		19'b0100101010100101011: color_data = Z;
		19'b0100101010100101100: color_data = Z;
		19'b0100101010100101101: color_data = Z;
		19'b0100101010100101110: color_data = Z;
		19'b0100101010100101111: color_data = Z;
		19'b0100101010100110000: color_data = Z;
		19'b0100101010100110001: color_data = Z;
		19'b0100101010100110010: color_data = Z;
		19'b0100101010100110011: color_data = Z;
		19'b0100101010100110100: color_data = Z;
		19'b0100101010100110101: color_data = Z;
		19'b0100101010100110110: color_data = Z;
		19'b0100101010100110111: color_data = Z;
		19'b0100101010100111000: color_data = Z;
		19'b0100101010100111001: color_data = Z;
		19'b0100101010100111010: color_data = Z;
		19'b0100101010100111011: color_data = Z;
		19'b0100101010100111100: color_data = Z;
		19'b0100101010100111101: color_data = Z;
		19'b0100101010100111110: color_data = Z;
		19'b0100101010100111111: color_data = Z;
		19'b0100101010101000000: color_data = Z;
		19'b0100101010101000001: color_data = Z;
		19'b0100101010101000010: color_data = Z;
		19'b0100101010101000011: color_data = Z;
		19'b0100101010101000100: color_data = Z;
		19'b0100101010101000101: color_data = Z;
		19'b0100101010101000110: color_data = Z;
		19'b0100101010101000111: color_data = Z;
		19'b0100101010101001000: color_data = Z;
		19'b0100101010101001001: color_data = Z;
		19'b0100101010101001010: color_data = Z;
		19'b0100101010101001011: color_data = Z;
		19'b0100101010101001100: color_data = Z;
		19'b0100101010101001101: color_data = Z;
		19'b0100101010101001110: color_data = Z;
		19'b0100101010101001111: color_data = Z;
		19'b0100101010101010000: color_data = Z;
		19'b0100101010101010001: color_data = Z;
		19'b0100101010101010010: color_data = Z;
		19'b0100101010101010011: color_data = Z;
		19'b0100101010101010100: color_data = Z;
		19'b0100101010101010101: color_data = Z;
		19'b0100101010101010110: color_data = Z;
		19'b0100101010101010111: color_data = Z;
		19'b0100101010101011000: color_data = Z;
		19'b0100101010101011001: color_data = Z;
		19'b0100101010101011010: color_data = Z;
		19'b0100101010101011011: color_data = Z;
		19'b0100101010101011100: color_data = Z;
		19'b0100101010101011101: color_data = Z;
		19'b0100101010101011110: color_data = Z;
		19'b0100101010101011111: color_data = Z;
		19'b0100101010101100000: color_data = Z;
		19'b0100101010101100001: color_data = Z;
		19'b0100101010101100010: color_data = Z;
		19'b0100101010101100011: color_data = Z;
		19'b0100101010101100100: color_data = Z;
		19'b0100101010101100101: color_data = Z;
		19'b0100101010101100110: color_data = Z;
		19'b0100101010101100111: color_data = Z;
		19'b0100101010101101000: color_data = Z;
		19'b0100101010101101001: color_data = Z;
		19'b0100101010101101010: color_data = Z;
		19'b0100101010101101011: color_data = Z;
		19'b0100101010101101100: color_data = Z;
		19'b0100101010101101101: color_data = Z;
		19'b0100101010101101110: color_data = Z;
		19'b0100101010101101111: color_data = Z;
		19'b0100101010101110000: color_data = Z;
		19'b0100101010101110001: color_data = Z;
		19'b0100101010101110010: color_data = Z;
		19'b0100101010101110011: color_data = Z;
		19'b0100101010101110100: color_data = Z;
		19'b0100101010101110101: color_data = Z;
		19'b0100101010101110110: color_data = Z;
		19'b0100101010101110111: color_data = Z;
		19'b0100101010101111000: color_data = Z;
		19'b0100101010101111001: color_data = Z;
		19'b0100101010101111010: color_data = Z;
		19'b0100101010101111011: color_data = Z;
		19'b0100101010101111100: color_data = Z;
		19'b0100101010101111101: color_data = Z;
		19'b0100101010101111110: color_data = Z;
		19'b0100101010101111111: color_data = Z;
		19'b0100101010110000000: color_data = Z;
		19'b0100101010111001110: color_data = Z;
		19'b0100101010111001111: color_data = Z;
		19'b0100101010111010000: color_data = Z;
		19'b0100101010111010001: color_data = Z;
		19'b0100101010111010010: color_data = Z;
		19'b0100101010111010011: color_data = Z;
		19'b0100101010111010100: color_data = Z;
		19'b0100101010111010101: color_data = Z;
		19'b0100101010111010110: color_data = Z;
		19'b0100101010111010111: color_data = Z;
		19'b0100101010111011000: color_data = Z;
		19'b0100101010111011001: color_data = Z;
		19'b0100101010111011010: color_data = Z;
		19'b0100101010111011011: color_data = Z;
		19'b0100101010111100010: color_data = Z;
		19'b0100101100100001111: color_data = Z;
		19'b0100101100100010000: color_data = Z;
		19'b0100101100100010001: color_data = Z;
		19'b0100101100100010010: color_data = Z;
		19'b0100101100100010011: color_data = Z;
		19'b0100101100100010100: color_data = Z;
		19'b0100101100100010101: color_data = Z;
		19'b0100101100100010110: color_data = Z;
		19'b0100101100100010111: color_data = Z;
		19'b0100101100100011000: color_data = Z;
		19'b0100101100100011001: color_data = Z;
		19'b0100101100100011010: color_data = Z;
		19'b0100101100100011011: color_data = Z;
		19'b0100101100100011100: color_data = Z;
		19'b0100101100100100011: color_data = Z;
		19'b0100101100100100100: color_data = Z;
		19'b0100101100100100101: color_data = Z;
		19'b0100101100100100110: color_data = Z;
		19'b0100101100100100111: color_data = Z;
		19'b0100101100100101000: color_data = Z;
		19'b0100101100100101001: color_data = Z;
		19'b0100101100100101010: color_data = Z;
		19'b0100101100100101011: color_data = Z;
		19'b0100101100100101100: color_data = Z;
		19'b0100101100100101101: color_data = Z;
		19'b0100101100100101110: color_data = Z;
		19'b0100101100100101111: color_data = Z;
		19'b0100101100100110000: color_data = Z;
		19'b0100101100100110001: color_data = Z;
		19'b0100101100100110010: color_data = Z;
		19'b0100101100100110011: color_data = Z;
		19'b0100101100100110100: color_data = Z;
		19'b0100101100100110101: color_data = Z;
		19'b0100101100100110110: color_data = Z;
		19'b0100101100100110111: color_data = Z;
		19'b0100101100100111000: color_data = Z;
		19'b0100101100100111001: color_data = Z;
		19'b0100101100100111010: color_data = Z;
		19'b0100101100100111011: color_data = Z;
		19'b0100101100100111100: color_data = Z;
		19'b0100101100100111101: color_data = Z;
		19'b0100101100100111110: color_data = Z;
		19'b0100101100100111111: color_data = Z;
		19'b0100101100101000000: color_data = Z;
		19'b0100101100101000001: color_data = Z;
		19'b0100101100101000010: color_data = Z;
		19'b0100101100101000011: color_data = Z;
		19'b0100101100101000100: color_data = Z;
		19'b0100101100101000101: color_data = Z;
		19'b0100101100101000110: color_data = Z;
		19'b0100101100101000111: color_data = Z;
		19'b0100101100101001000: color_data = Z;
		19'b0100101100101001001: color_data = Z;
		19'b0100101100101001010: color_data = Z;
		19'b0100101100101001011: color_data = Z;
		19'b0100101100101001100: color_data = Z;
		19'b0100101100101001101: color_data = Z;
		19'b0100101100101001110: color_data = Z;
		19'b0100101100101001111: color_data = Z;
		19'b0100101100101010000: color_data = Z;
		19'b0100101100101010001: color_data = Z;
		19'b0100101100101010010: color_data = Z;
		19'b0100101100101010011: color_data = Z;
		19'b0100101100101010100: color_data = Z;
		19'b0100101100101010101: color_data = Z;
		19'b0100101100101010110: color_data = Z;
		19'b0100101100101010111: color_data = Z;
		19'b0100101100101011000: color_data = Z;
		19'b0100101100101011001: color_data = Z;
		19'b0100101100101011010: color_data = Z;
		19'b0100101100101011011: color_data = Z;
		19'b0100101100101011100: color_data = Z;
		19'b0100101100101011101: color_data = Z;
		19'b0100101100101011110: color_data = Z;
		19'b0100101100101011111: color_data = Z;
		19'b0100101100101100000: color_data = Z;
		19'b0100101100101100001: color_data = Z;
		19'b0100101100101100010: color_data = Z;
		19'b0100101100101100011: color_data = Z;
		19'b0100101100101100100: color_data = Z;
		19'b0100101100101100101: color_data = Z;
		19'b0100101100101100110: color_data = Z;
		19'b0100101100101100111: color_data = Z;
		19'b0100101100101101000: color_data = Z;
		19'b0100101100101101001: color_data = Z;
		19'b0100101100101101010: color_data = Z;
		19'b0100101100101101011: color_data = Z;
		19'b0100101100101101100: color_data = Z;
		19'b0100101100101101101: color_data = Z;
		19'b0100101100101101110: color_data = Z;
		19'b0100101100101101111: color_data = Z;
		19'b0100101100101110000: color_data = Z;
		19'b0100101100101110001: color_data = Z;
		19'b0100101100101110010: color_data = Z;
		19'b0100101100101110011: color_data = Z;
		19'b0100101100101110100: color_data = Z;
		19'b0100101100101110101: color_data = Z;
		19'b0100101100101110110: color_data = Z;
		19'b0100101100101110111: color_data = Z;
		19'b0100101100101111000: color_data = Z;
		19'b0100101100101111001: color_data = Z;
		19'b0100101100101111010: color_data = Z;
		19'b0100101100101111011: color_data = Z;
		19'b0100101100101111100: color_data = Z;
		19'b0100101100101111101: color_data = Z;
		19'b0100101100101111110: color_data = Z;
		19'b0100101100101111111: color_data = Z;
		19'b0100101100110000000: color_data = Z;
		19'b0100101100111001110: color_data = Z;
		19'b0100101100111001111: color_data = Z;
		19'b0100101100111010000: color_data = Z;
		19'b0100101100111010001: color_data = Z;
		19'b0100101100111010010: color_data = Z;
		19'b0100101100111010011: color_data = Z;
		19'b0100101100111010100: color_data = Z;
		19'b0100101100111010101: color_data = Z;
		19'b0100101100111010110: color_data = Z;
		19'b0100101100111010111: color_data = Z;
		19'b0100101100111011000: color_data = Z;
		19'b0100101100111011001: color_data = Z;
		19'b0100101100111011010: color_data = Z;
		19'b0100101100111011011: color_data = Z;
		19'b0100101100111011100: color_data = Z;
		19'b0100101110100010000: color_data = Z;
		19'b0100101110100010001: color_data = Z;
		19'b0100101110100010010: color_data = Z;
		19'b0100101110100010011: color_data = Z;
		19'b0100101110100010100: color_data = Z;
		19'b0100101110100010101: color_data = Z;
		19'b0100101110100010110: color_data = Z;
		19'b0100101110100010111: color_data = Z;
		19'b0100101110100011000: color_data = Z;
		19'b0100101110100011001: color_data = Z;
		19'b0100101110100011010: color_data = Z;
		19'b0100101110100011011: color_data = Z;
		19'b0100101110100100100: color_data = Z;
		19'b0100101110100100101: color_data = Z;
		19'b0100101110100100110: color_data = Z;
		19'b0100101110100100111: color_data = Z;
		19'b0100101110100101000: color_data = Z;
		19'b0100101110100101001: color_data = Z;
		19'b0100101110100101010: color_data = Z;
		19'b0100101110100101011: color_data = Z;
		19'b0100101110100101100: color_data = Z;
		19'b0100101110100101101: color_data = Z;
		19'b0100101110100101110: color_data = Z;
		19'b0100101110100101111: color_data = Z;
		19'b0100101110100110000: color_data = Z;
		19'b0100101110100110001: color_data = Z;
		19'b0100101110100110010: color_data = Z;
		19'b0100101110100110011: color_data = Z;
		19'b0100101110100110100: color_data = Z;
		19'b0100101110100110101: color_data = Z;
		19'b0100101110100110110: color_data = Z;
		19'b0100101110100110111: color_data = Z;
		19'b0100101110100111000: color_data = Z;
		19'b0100101110100111001: color_data = Z;
		19'b0100101110100111010: color_data = Z;
		19'b0100101110100111011: color_data = Z;
		19'b0100101110100111100: color_data = Z;
		19'b0100101110100111101: color_data = Z;
		19'b0100101110100111110: color_data = Z;
		19'b0100101110100111111: color_data = Z;
		19'b0100101110101000000: color_data = Z;
		19'b0100101110101000001: color_data = Z;
		19'b0100101110101000010: color_data = Z;
		19'b0100101110101000011: color_data = Z;
		19'b0100101110101000100: color_data = Z;
		19'b0100101110101000101: color_data = Z;
		19'b0100101110101000110: color_data = Z;
		19'b0100101110101000111: color_data = Z;
		19'b0100101110101001000: color_data = Z;
		19'b0100101110101001001: color_data = Z;
		19'b0100101110101001010: color_data = Z;
		19'b0100101110101001011: color_data = Z;
		19'b0100101110101001100: color_data = Z;
		19'b0100101110101001101: color_data = Z;
		19'b0100101110101001110: color_data = Z;
		19'b0100101110101001111: color_data = Z;
		19'b0100101110101010000: color_data = Z;
		19'b0100101110101010001: color_data = Z;
		19'b0100101110101010010: color_data = Z;
		19'b0100101110101010011: color_data = Z;
		19'b0100101110101010100: color_data = Z;
		19'b0100101110101010101: color_data = Z;
		19'b0100101110101010110: color_data = Z;
		19'b0100101110101010111: color_data = Z;
		19'b0100101110101011000: color_data = Z;
		19'b0100101110101011001: color_data = Z;
		19'b0100101110101011010: color_data = Z;
		19'b0100101110101011011: color_data = Z;
		19'b0100101110101011100: color_data = Z;
		19'b0100101110101011101: color_data = Z;
		19'b0100101110101011110: color_data = Z;
		19'b0100101110101011111: color_data = Z;
		19'b0100101110101100000: color_data = Z;
		19'b0100101110101100001: color_data = Z;
		19'b0100101110101100010: color_data = Z;
		19'b0100101110101100011: color_data = Z;
		19'b0100101110101100100: color_data = Z;
		19'b0100101110101100101: color_data = Z;
		19'b0100101110101100110: color_data = Z;
		19'b0100101110101100111: color_data = Z;
		19'b0100101110101101000: color_data = Z;
		19'b0100101110101101001: color_data = Z;
		19'b0100101110101101010: color_data = Z;
		19'b0100101110101101011: color_data = Z;
		19'b0100101110101101100: color_data = Z;
		19'b0100101110101101101: color_data = Z;
		19'b0100101110101101110: color_data = Z;
		19'b0100101110101101111: color_data = Z;
		19'b0100101110101110000: color_data = Z;
		19'b0100101110101110001: color_data = Z;
		19'b0100101110101110010: color_data = Z;
		19'b0100101110101110011: color_data = Z;
		19'b0100101110101110100: color_data = Z;
		19'b0100101110101110101: color_data = Z;
		19'b0100101110101110110: color_data = Z;
		19'b0100101110101110111: color_data = Z;
		19'b0100101110101111000: color_data = Z;
		19'b0100101110101111001: color_data = Z;
		19'b0100101110101111010: color_data = Z;
		19'b0100101110101111011: color_data = Z;
		19'b0100101110101111100: color_data = Z;
		19'b0100101110101111101: color_data = Z;
		19'b0100101110101111110: color_data = Z;
		19'b0100101110101111111: color_data = Z;
		19'b0100101110110000000: color_data = Z;
		19'b0100101110111001110: color_data = Z;
		19'b0100101110111001111: color_data = Z;
		19'b0100101110111010000: color_data = Z;
		19'b0100101110111010001: color_data = Z;
		19'b0100101110111010010: color_data = Z;
		19'b0100101110111010011: color_data = Z;
		19'b0100101110111010100: color_data = Z;
		19'b0100101110111010101: color_data = Z;
		19'b0100101110111010110: color_data = Z;
		19'b0100101110111010111: color_data = Z;
		19'b0100101110111011000: color_data = Z;
		19'b0100101110111011001: color_data = Z;
		19'b0100101110111011010: color_data = Z;
		19'b0100101110111011011: color_data = Z;
		19'b0100101110111011100: color_data = Z;
		19'b0100110000100010001: color_data = Z;
		19'b0100110000100010010: color_data = Z;
		19'b0100110000100010011: color_data = Z;
		19'b0100110000100010100: color_data = Z;
		19'b0100110000100010101: color_data = Z;
		19'b0100110000100010110: color_data = Z;
		19'b0100110000100010111: color_data = Z;
		19'b0100110000100011000: color_data = Z;
		19'b0100110000100011001: color_data = Z;
		19'b0100110000100011010: color_data = Z;
		19'b0100110000100011011: color_data = Z;
		19'b0100110000100011100: color_data = Z;
		19'b0100110000100100100: color_data = Z;
		19'b0100110000100100101: color_data = Z;
		19'b0100110000100100110: color_data = Z;
		19'b0100110000100100111: color_data = Z;
		19'b0100110000100101000: color_data = Z;
		19'b0100110000100101001: color_data = Z;
		19'b0100110000100101010: color_data = Z;
		19'b0100110000100101011: color_data = Z;
		19'b0100110000100101100: color_data = Z;
		19'b0100110000100101101: color_data = Z;
		19'b0100110000100101110: color_data = Z;
		19'b0100110000100101111: color_data = Z;
		19'b0100110000100110000: color_data = Z;
		19'b0100110000100110001: color_data = Z;
		19'b0100110000100110010: color_data = Z;
		19'b0100110000100110011: color_data = Z;
		19'b0100110000100110100: color_data = Z;
		19'b0100110000100110101: color_data = Z;
		19'b0100110000100110110: color_data = Z;
		19'b0100110000100110111: color_data = Z;
		19'b0100110000100111000: color_data = Z;
		19'b0100110000100111001: color_data = Z;
		19'b0100110000100111010: color_data = Z;
		19'b0100110000100111011: color_data = Z;
		19'b0100110000100111100: color_data = Z;
		19'b0100110000100111101: color_data = Z;
		19'b0100110000100111110: color_data = Z;
		19'b0100110000100111111: color_data = Z;
		19'b0100110000101000000: color_data = Z;
		19'b0100110000101000001: color_data = Z;
		19'b0100110000101000010: color_data = Z;
		19'b0100110000101000011: color_data = Z;
		19'b0100110000101000100: color_data = Z;
		19'b0100110000101000101: color_data = Z;
		19'b0100110000101000110: color_data = Z;
		19'b0100110000101000111: color_data = Z;
		19'b0100110000101001000: color_data = Z;
		19'b0100110000101001001: color_data = Z;
		19'b0100110000101001010: color_data = Z;
		19'b0100110000101001011: color_data = Z;
		19'b0100110000101001100: color_data = Z;
		19'b0100110000101001101: color_data = Z;
		19'b0100110000101001110: color_data = Z;
		19'b0100110000101001111: color_data = Z;
		19'b0100110000101010000: color_data = Z;
		19'b0100110000101010001: color_data = Z;
		19'b0100110000101010010: color_data = Z;
		19'b0100110000101010011: color_data = Z;
		19'b0100110000101010100: color_data = Z;
		19'b0100110000101010101: color_data = Z;
		19'b0100110000101010110: color_data = Z;
		19'b0100110000101010111: color_data = Z;
		19'b0100110000101011000: color_data = Z;
		19'b0100110000101011001: color_data = Z;
		19'b0100110000101011010: color_data = Z;
		19'b0100110000101011011: color_data = Z;
		19'b0100110000101011100: color_data = Z;
		19'b0100110000101011101: color_data = Z;
		19'b0100110000101011110: color_data = Z;
		19'b0100110000101011111: color_data = Z;
		19'b0100110000101100000: color_data = Z;
		19'b0100110000101100001: color_data = Z;
		19'b0100110000101100010: color_data = Z;
		19'b0100110000101100011: color_data = Z;
		19'b0100110000101100100: color_data = Z;
		19'b0100110000101100101: color_data = Z;
		19'b0100110000101100110: color_data = Z;
		19'b0100110000101100111: color_data = Z;
		19'b0100110000101101000: color_data = Z;
		19'b0100110000101101001: color_data = Z;
		19'b0100110000101101010: color_data = Z;
		19'b0100110000101101011: color_data = Z;
		19'b0100110000101101100: color_data = Z;
		19'b0100110000101101101: color_data = Z;
		19'b0100110000101101110: color_data = Z;
		19'b0100110000101101111: color_data = Z;
		19'b0100110000101110000: color_data = Z;
		19'b0100110000101110001: color_data = Z;
		19'b0100110000101110010: color_data = Z;
		19'b0100110000101110011: color_data = Z;
		19'b0100110000101110100: color_data = Z;
		19'b0100110000101110101: color_data = Z;
		19'b0100110000101110110: color_data = Z;
		19'b0100110000101110111: color_data = Z;
		19'b0100110000101111000: color_data = Z;
		19'b0100110000101111001: color_data = Z;
		19'b0100110000101111010: color_data = Z;
		19'b0100110000101111011: color_data = Z;
		19'b0100110000101111100: color_data = Z;
		19'b0100110000101111101: color_data = Z;
		19'b0100110000101111110: color_data = Z;
		19'b0100110000101111111: color_data = Z;
		19'b0100110000110000000: color_data = Z;
		19'b0100110000111001110: color_data = Z;
		19'b0100110000111001111: color_data = Z;
		19'b0100110000111010000: color_data = Z;
		19'b0100110000111010001: color_data = Z;
		19'b0100110000111010010: color_data = Z;
		19'b0100110000111010011: color_data = Z;
		19'b0100110000111010100: color_data = Z;
		19'b0100110000111010101: color_data = Z;
		19'b0100110000111010110: color_data = Z;
		19'b0100110000111010111: color_data = Z;
		19'b0100110000111011000: color_data = Z;
		19'b0100110000111011001: color_data = Z;
		19'b0100110000111011010: color_data = Z;
		19'b0100110000111011011: color_data = Z;
		19'b0100110000111011100: color_data = Z;
		19'b0100110000111011101: color_data = Z;
		19'b0100110010100010010: color_data = Z;
		19'b0100110010100010011: color_data = Z;
		19'b0100110010100010100: color_data = Z;
		19'b0100110010100010101: color_data = Z;
		19'b0100110010100010110: color_data = Z;
		19'b0100110010100010111: color_data = Z;
		19'b0100110010100011000: color_data = Z;
		19'b0100110010100011001: color_data = Z;
		19'b0100110010100011010: color_data = Z;
		19'b0100110010100011011: color_data = Z;
		19'b0100110010100011100: color_data = Z;
		19'b0100110010100100110: color_data = Z;
		19'b0100110010100100111: color_data = Z;
		19'b0100110010100101000: color_data = Z;
		19'b0100110010100101001: color_data = Z;
		19'b0100110010100101010: color_data = Z;
		19'b0100110010100101011: color_data = Z;
		19'b0100110010100101100: color_data = Z;
		19'b0100110010100101101: color_data = Z;
		19'b0100110010100101110: color_data = Z;
		19'b0100110010100101111: color_data = Z;
		19'b0100110010100110000: color_data = Z;
		19'b0100110010100110001: color_data = Z;
		19'b0100110010100110010: color_data = Z;
		19'b0100110010100110011: color_data = Z;
		19'b0100110010100110100: color_data = Z;
		19'b0100110010100110101: color_data = Z;
		19'b0100110010100110110: color_data = Z;
		19'b0100110010100110111: color_data = Z;
		19'b0100110010100111000: color_data = Z;
		19'b0100110010100111001: color_data = Z;
		19'b0100110010100111010: color_data = Z;
		19'b0100110010100111011: color_data = Z;
		19'b0100110010100111100: color_data = Z;
		19'b0100110010100111101: color_data = Z;
		19'b0100110010100111110: color_data = Z;
		19'b0100110010100111111: color_data = Z;
		19'b0100110010101000000: color_data = Z;
		19'b0100110010101000001: color_data = Z;
		19'b0100110010101000010: color_data = Z;
		19'b0100110010101000011: color_data = Z;
		19'b0100110010101000100: color_data = Z;
		19'b0100110010101000101: color_data = Z;
		19'b0100110010101000110: color_data = Z;
		19'b0100110010101000111: color_data = Z;
		19'b0100110010101001000: color_data = Z;
		19'b0100110010101001001: color_data = Z;
		19'b0100110010101001010: color_data = Z;
		19'b0100110010101001011: color_data = Z;
		19'b0100110010101001100: color_data = Z;
		19'b0100110010101001101: color_data = Z;
		19'b0100110010101001110: color_data = Z;
		19'b0100110010101001111: color_data = Z;
		19'b0100110010101010000: color_data = Z;
		19'b0100110010101010001: color_data = Z;
		19'b0100110010101010010: color_data = Z;
		19'b0100110010101010011: color_data = Z;
		19'b0100110010101010100: color_data = Z;
		19'b0100110010101010101: color_data = Z;
		19'b0100110010101010110: color_data = Z;
		19'b0100110010101010111: color_data = Z;
		19'b0100110010101011000: color_data = Z;
		19'b0100110010101011001: color_data = Z;
		19'b0100110010101011010: color_data = Z;
		19'b0100110010101011011: color_data = Z;
		19'b0100110010101011100: color_data = Z;
		19'b0100110010101011101: color_data = Z;
		19'b0100110010101011110: color_data = Z;
		19'b0100110010101011111: color_data = Z;
		19'b0100110010101100000: color_data = Z;
		19'b0100110010101100001: color_data = Z;
		19'b0100110010101100010: color_data = Z;
		19'b0100110010101100011: color_data = Z;
		19'b0100110010101100100: color_data = Z;
		19'b0100110010101100101: color_data = Z;
		19'b0100110010101100110: color_data = Z;
		19'b0100110010101100111: color_data = Z;
		19'b0100110010101101000: color_data = Z;
		19'b0100110010101101001: color_data = Z;
		19'b0100110010101101010: color_data = Z;
		19'b0100110010101101011: color_data = Z;
		19'b0100110010101101100: color_data = Z;
		19'b0100110010101101101: color_data = Z;
		19'b0100110010101101110: color_data = Z;
		19'b0100110010101101111: color_data = Z;
		19'b0100110010101110000: color_data = Z;
		19'b0100110010101110001: color_data = Z;
		19'b0100110010101110010: color_data = Z;
		19'b0100110010101110011: color_data = Z;
		19'b0100110010101110100: color_data = Z;
		19'b0100110010101110101: color_data = Z;
		19'b0100110010101110110: color_data = Z;
		19'b0100110010101110111: color_data = Z;
		19'b0100110010101111000: color_data = Z;
		19'b0100110010101111001: color_data = Z;
		19'b0100110010101111010: color_data = Z;
		19'b0100110010101111011: color_data = Z;
		19'b0100110010101111100: color_data = Z;
		19'b0100110010101111101: color_data = Z;
		19'b0100110010101111110: color_data = Z;
		19'b0100110010101111111: color_data = Z;
		19'b0100110010110000000: color_data = Z;
		19'b0100110010111001110: color_data = Z;
		19'b0100110010111001111: color_data = Z;
		19'b0100110010111010000: color_data = Z;
		19'b0100110010111010001: color_data = Z;
		19'b0100110010111010010: color_data = Z;
		19'b0100110010111010011: color_data = Z;
		19'b0100110010111010100: color_data = Z;
		19'b0100110010111010101: color_data = Z;
		19'b0100110010111010110: color_data = Z;
		19'b0100110010111010111: color_data = Z;
		19'b0100110010111011000: color_data = Z;
		19'b0100110010111011001: color_data = Z;
		19'b0100110010111011010: color_data = Z;
		19'b0100110010111011011: color_data = Z;
		19'b0100110010111011100: color_data = Z;
		19'b0100110010111011101: color_data = Z;
		19'b0100110100100010011: color_data = Z;
		19'b0100110100100010100: color_data = Z;
		19'b0100110100100010101: color_data = Z;
		19'b0100110100100010110: color_data = Z;
		19'b0100110100100010111: color_data = Z;
		19'b0100110100100011000: color_data = Z;
		19'b0100110100100011001: color_data = Z;
		19'b0100110100100011010: color_data = Z;
		19'b0100110100100011011: color_data = Z;
		19'b0100110100100011110: color_data = Z;
		19'b0100110100100011111: color_data = Z;
		19'b0100110100100100110: color_data = Z;
		19'b0100110100100100111: color_data = Z;
		19'b0100110100100101000: color_data = Z;
		19'b0100110100100101001: color_data = Z;
		19'b0100110100100101010: color_data = Z;
		19'b0100110100100101011: color_data = Z;
		19'b0100110100100101100: color_data = Z;
		19'b0100110100100101101: color_data = Z;
		19'b0100110100100101110: color_data = Z;
		19'b0100110100100101111: color_data = Z;
		19'b0100110100100110000: color_data = Z;
		19'b0100110100100110001: color_data = Z;
		19'b0100110100100110010: color_data = Z;
		19'b0100110100100110011: color_data = Z;
		19'b0100110100100110100: color_data = Z;
		19'b0100110100100110101: color_data = Z;
		19'b0100110100100110110: color_data = Z;
		19'b0100110100100110111: color_data = Z;
		19'b0100110100100111000: color_data = Z;
		19'b0100110100100111001: color_data = Z;
		19'b0100110100100111010: color_data = Z;
		19'b0100110100100111011: color_data = Z;
		19'b0100110100100111100: color_data = Z;
		19'b0100110100100111101: color_data = Z;
		19'b0100110100100111110: color_data = Z;
		19'b0100110100100111111: color_data = Z;
		19'b0100110100101000000: color_data = Z;
		19'b0100110100101000001: color_data = Z;
		19'b0100110100101000010: color_data = Z;
		19'b0100110100101000011: color_data = Z;
		19'b0100110100101000100: color_data = Z;
		19'b0100110100101000101: color_data = Z;
		19'b0100110100101000110: color_data = Z;
		19'b0100110100101000111: color_data = Z;
		19'b0100110100101001000: color_data = Z;
		19'b0100110100101001001: color_data = Z;
		19'b0100110100101001010: color_data = Z;
		19'b0100110100101001011: color_data = Z;
		19'b0100110100101001100: color_data = Z;
		19'b0100110100101001101: color_data = Z;
		19'b0100110100101001110: color_data = Z;
		19'b0100110100101001111: color_data = Z;
		19'b0100110100101010000: color_data = Z;
		19'b0100110100101010001: color_data = Z;
		19'b0100110100101010010: color_data = Z;
		19'b0100110100101010011: color_data = Z;
		19'b0100110100101010100: color_data = Z;
		19'b0100110100101010101: color_data = Z;
		19'b0100110100101010110: color_data = Z;
		19'b0100110100101010111: color_data = Z;
		19'b0100110100101011000: color_data = Z;
		19'b0100110100101011001: color_data = Z;
		19'b0100110100101011010: color_data = Z;
		19'b0100110100101011011: color_data = Z;
		19'b0100110100101011100: color_data = Z;
		19'b0100110100101011101: color_data = Z;
		19'b0100110100101011110: color_data = Z;
		19'b0100110100101011111: color_data = Z;
		19'b0100110100101100000: color_data = Z;
		19'b0100110100101100001: color_data = Z;
		19'b0100110100101100010: color_data = Z;
		19'b0100110100101100011: color_data = Z;
		19'b0100110100101100100: color_data = Z;
		19'b0100110100101100101: color_data = Z;
		19'b0100110100101100110: color_data = Z;
		19'b0100110100101100111: color_data = Z;
		19'b0100110100101101000: color_data = Z;
		19'b0100110100101101001: color_data = Z;
		19'b0100110100101101010: color_data = Z;
		19'b0100110100101101011: color_data = Z;
		19'b0100110100101101100: color_data = Z;
		19'b0100110100101101101: color_data = Z;
		19'b0100110100101101110: color_data = Z;
		19'b0100110100101101111: color_data = Z;
		19'b0100110100101110000: color_data = Z;
		19'b0100110100101110001: color_data = Z;
		19'b0100110100101110010: color_data = Z;
		19'b0100110100101110011: color_data = Z;
		19'b0100110100101110100: color_data = Z;
		19'b0100110100101110101: color_data = Z;
		19'b0100110100101110110: color_data = Z;
		19'b0100110100101110111: color_data = Z;
		19'b0100110100101111000: color_data = Z;
		19'b0100110100101111001: color_data = Z;
		19'b0100110100101111010: color_data = Z;
		19'b0100110100101111011: color_data = Z;
		19'b0100110100101111100: color_data = Z;
		19'b0100110100101111101: color_data = Z;
		19'b0100110100101111110: color_data = Z;
		19'b0100110100101111111: color_data = Z;
		19'b0100110100110000000: color_data = Z;
		19'b0100110100111001110: color_data = Z;
		19'b0100110100111001111: color_data = Z;
		19'b0100110100111010000: color_data = Z;
		19'b0100110100111010001: color_data = Z;
		19'b0100110100111010010: color_data = Z;
		19'b0100110100111010011: color_data = Z;
		19'b0100110100111010100: color_data = Z;
		19'b0100110100111010101: color_data = Z;
		19'b0100110100111010110: color_data = Z;
		19'b0100110100111010111: color_data = Z;
		19'b0100110100111011000: color_data = Z;
		19'b0100110100111011001: color_data = Z;
		19'b0100110100111011010: color_data = Z;
		19'b0100110100111011011: color_data = Z;
		19'b0100110100111011100: color_data = Z;
		19'b0100110100111011101: color_data = Z;
		19'b0100110100111011110: color_data = Z;
		19'b0100110100111011111: color_data = Z;
		19'b0100110110100010100: color_data = Z;
		19'b0100110110100010101: color_data = Z;
		19'b0100110110100010110: color_data = Z;
		19'b0100110110100010111: color_data = Z;
		19'b0100110110100011000: color_data = Z;
		19'b0100110110100011001: color_data = Z;
		19'b0100110110100011110: color_data = Z;
		19'b0100110110100011111: color_data = Z;
		19'b0100110110100100111: color_data = Z;
		19'b0100110110100101000: color_data = Z;
		19'b0100110110100101001: color_data = Z;
		19'b0100110110100101010: color_data = Z;
		19'b0100110110100101011: color_data = Z;
		19'b0100110110100101100: color_data = Z;
		19'b0100110110100101101: color_data = Z;
		19'b0100110110100101110: color_data = Z;
		19'b0100110110100101111: color_data = Z;
		19'b0100110110100110000: color_data = Z;
		19'b0100110110100110001: color_data = Z;
		19'b0100110110100110010: color_data = Z;
		19'b0100110110100110011: color_data = Z;
		19'b0100110110100110100: color_data = Z;
		19'b0100110110100110101: color_data = Z;
		19'b0100110110100110110: color_data = Z;
		19'b0100110110100110111: color_data = Z;
		19'b0100110110100111000: color_data = Z;
		19'b0100110110100111001: color_data = Z;
		19'b0100110110100111010: color_data = Z;
		19'b0100110110100111011: color_data = Z;
		19'b0100110110100111100: color_data = Z;
		19'b0100110110100111101: color_data = Z;
		19'b0100110110100111110: color_data = Z;
		19'b0100110110100111111: color_data = Z;
		19'b0100110110101000000: color_data = Z;
		19'b0100110110101000001: color_data = Z;
		19'b0100110110101000010: color_data = Z;
		19'b0100110110101000011: color_data = Z;
		19'b0100110110101000100: color_data = Z;
		19'b0100110110101000101: color_data = Z;
		19'b0100110110101000110: color_data = Z;
		19'b0100110110101000111: color_data = Z;
		19'b0100110110101001000: color_data = Z;
		19'b0100110110101001001: color_data = Z;
		19'b0100110110101001010: color_data = Z;
		19'b0100110110101001011: color_data = Z;
		19'b0100110110101001100: color_data = Z;
		19'b0100110110101001101: color_data = Z;
		19'b0100110110101001110: color_data = Z;
		19'b0100110110101001111: color_data = Z;
		19'b0100110110101010000: color_data = Z;
		19'b0100110110101010001: color_data = Z;
		19'b0100110110101010010: color_data = Z;
		19'b0100110110101010011: color_data = Z;
		19'b0100110110101010100: color_data = Z;
		19'b0100110110101010101: color_data = Z;
		19'b0100110110101010110: color_data = Z;
		19'b0100110110101010111: color_data = Z;
		19'b0100110110101011000: color_data = Z;
		19'b0100110110101011001: color_data = Z;
		19'b0100110110101011010: color_data = Z;
		19'b0100110110101011011: color_data = Z;
		19'b0100110110101011100: color_data = Z;
		19'b0100110110101011101: color_data = Z;
		19'b0100110110101011110: color_data = Z;
		19'b0100110110101011111: color_data = Z;
		19'b0100110110101100000: color_data = Z;
		19'b0100110110101100001: color_data = Z;
		19'b0100110110101100010: color_data = Z;
		19'b0100110110101100011: color_data = Z;
		19'b0100110110101100100: color_data = Z;
		19'b0100110110101100101: color_data = Z;
		19'b0100110110101100110: color_data = Z;
		19'b0100110110101100111: color_data = Z;
		19'b0100110110101101000: color_data = Z;
		19'b0100110110101101001: color_data = Z;
		19'b0100110110101101010: color_data = Z;
		19'b0100110110101101011: color_data = Z;
		19'b0100110110101101100: color_data = Z;
		19'b0100110110101101101: color_data = Z;
		19'b0100110110101101110: color_data = Z;
		19'b0100110110101101111: color_data = Z;
		19'b0100110110101110000: color_data = Z;
		19'b0100110110101110001: color_data = Z;
		19'b0100110110101110010: color_data = Z;
		19'b0100110110101110011: color_data = Z;
		19'b0100110110101110100: color_data = Z;
		19'b0100110110101110101: color_data = Z;
		19'b0100110110101110110: color_data = Z;
		19'b0100110110101110111: color_data = Z;
		19'b0100110110101111000: color_data = Z;
		19'b0100110110101111001: color_data = Z;
		19'b0100110110101111010: color_data = Z;
		19'b0100110110101111011: color_data = Z;
		19'b0100110110101111100: color_data = Z;
		19'b0100110110101111101: color_data = Z;
		19'b0100110110101111110: color_data = Z;
		19'b0100110110101111111: color_data = Z;
		19'b0100110110110000000: color_data = Z;
		19'b0100110110111001110: color_data = Z;
		19'b0100110110111001111: color_data = Z;
		19'b0100110110111010000: color_data = Z;
		19'b0100110110111010001: color_data = Z;
		19'b0100110110111010010: color_data = Z;
		19'b0100110110111010011: color_data = Z;
		19'b0100110110111010100: color_data = Z;
		19'b0100110110111010101: color_data = Z;
		19'b0100110110111010110: color_data = Z;
		19'b0100110110111010111: color_data = Z;
		19'b0100110110111011000: color_data = Z;
		19'b0100110110111011001: color_data = Z;
		19'b0100110110111011010: color_data = Z;
		19'b0100110110111011011: color_data = Z;
		19'b0100110110111011100: color_data = Z;
		19'b0100110110111011101: color_data = Z;
		19'b0100110110111011110: color_data = Z;
		19'b0100110110111011111: color_data = Z;
		19'b0100111000100010110: color_data = Z;
		19'b0100111000100010111: color_data = Z;
		19'b0100111000100011000: color_data = Z;
		19'b0100111000100011001: color_data = Z;
		19'b0100111000100011010: color_data = Z;
		19'b0100111000100011110: color_data = Z;
		19'b0100111000100011111: color_data = Z;
		19'b0100111000100101001: color_data = Z;
		19'b0100111000100101010: color_data = Z;
		19'b0100111000100101011: color_data = Z;
		19'b0100111000100101100: color_data = Z;
		19'b0100111000100101101: color_data = Z;
		19'b0100111000100101110: color_data = Z;
		19'b0100111000100101111: color_data = Z;
		19'b0100111000100110000: color_data = Z;
		19'b0100111000100110001: color_data = Z;
		19'b0100111000100110010: color_data = Z;
		19'b0100111000100110011: color_data = Z;
		19'b0100111000100110100: color_data = Z;
		19'b0100111000100110101: color_data = Z;
		19'b0100111000100110110: color_data = Z;
		19'b0100111000100110111: color_data = Z;
		19'b0100111000100111000: color_data = Z;
		19'b0100111000100111001: color_data = Z;
		19'b0100111000100111010: color_data = Z;
		19'b0100111000100111011: color_data = Z;
		19'b0100111000100111100: color_data = Z;
		19'b0100111000100111101: color_data = Z;
		19'b0100111000100111110: color_data = Z;
		19'b0100111000100111111: color_data = Z;
		19'b0100111000101000000: color_data = Z;
		19'b0100111000101000001: color_data = Z;
		19'b0100111000101000010: color_data = Z;
		19'b0100111000101000011: color_data = Z;
		19'b0100111000101000100: color_data = Z;
		19'b0100111000101000101: color_data = Z;
		19'b0100111000101000110: color_data = Z;
		19'b0100111000101000111: color_data = Z;
		19'b0100111000101001000: color_data = Z;
		19'b0100111000101001001: color_data = Z;
		19'b0100111000101001010: color_data = Z;
		19'b0100111000101001011: color_data = Z;
		19'b0100111000101001100: color_data = Z;
		19'b0100111000101001101: color_data = Z;
		19'b0100111000101001110: color_data = Z;
		19'b0100111000101001111: color_data = Z;
		19'b0100111000101010000: color_data = Z;
		19'b0100111000101010001: color_data = Z;
		19'b0100111000101010010: color_data = Z;
		19'b0100111000101010011: color_data = Z;
		19'b0100111000101010100: color_data = Z;
		19'b0100111000101010101: color_data = Z;
		19'b0100111000101010110: color_data = Z;
		19'b0100111000101010111: color_data = Z;
		19'b0100111000101011000: color_data = Z;
		19'b0100111000101011001: color_data = Z;
		19'b0100111000101011010: color_data = Z;
		19'b0100111000101011011: color_data = Z;
		19'b0100111000101011100: color_data = Z;
		19'b0100111000101011101: color_data = Z;
		19'b0100111000101011110: color_data = Z;
		19'b0100111000101011111: color_data = Z;
		19'b0100111000101100000: color_data = Z;
		19'b0100111000101100001: color_data = Z;
		19'b0100111000101100010: color_data = Z;
		19'b0100111000101100011: color_data = Z;
		19'b0100111000101100100: color_data = Z;
		19'b0100111000101100101: color_data = Z;
		19'b0100111000101100110: color_data = Z;
		19'b0100111000101100111: color_data = Z;
		19'b0100111000101101000: color_data = Z;
		19'b0100111000101101001: color_data = Z;
		19'b0100111000101101010: color_data = Z;
		19'b0100111000101101011: color_data = Z;
		19'b0100111000101101100: color_data = Z;
		19'b0100111000101101101: color_data = Z;
		19'b0100111000101101110: color_data = Z;
		19'b0100111000101101111: color_data = Z;
		19'b0100111000101110000: color_data = Z;
		19'b0100111000101110001: color_data = Z;
		19'b0100111000101110010: color_data = Z;
		19'b0100111000101110011: color_data = Z;
		19'b0100111000101110100: color_data = Z;
		19'b0100111000101110101: color_data = Z;
		19'b0100111000101110110: color_data = Z;
		19'b0100111000101110111: color_data = Z;
		19'b0100111000101111000: color_data = Z;
		19'b0100111000101111001: color_data = Z;
		19'b0100111000101111010: color_data = Z;
		19'b0100111000101111011: color_data = Z;
		19'b0100111000101111100: color_data = Z;
		19'b0100111000101111101: color_data = Z;
		19'b0100111000101111110: color_data = Z;
		19'b0100111000101111111: color_data = Z;
		19'b0100111000110000000: color_data = Z;
		19'b0100111000111001110: color_data = Z;
		19'b0100111000111001111: color_data = Z;
		19'b0100111000111010000: color_data = Z;
		19'b0100111000111010001: color_data = Z;
		19'b0100111000111010010: color_data = Z;
		19'b0100111000111010011: color_data = Z;
		19'b0100111000111010100: color_data = Z;
		19'b0100111000111010101: color_data = Z;
		19'b0100111000111010110: color_data = Z;
		19'b0100111000111010111: color_data = Z;
		19'b0100111000111011000: color_data = Z;
		19'b0100111000111011001: color_data = Z;
		19'b0100111000111011010: color_data = Z;
		19'b0100111000111011011: color_data = Z;
		19'b0100111000111011100: color_data = Z;
		19'b0100111000111011101: color_data = Z;
		19'b0100111000111011110: color_data = Z;
		19'b0100111000111011111: color_data = Z;
		19'b0100111000111100000: color_data = Z;
		19'b0100111000111100001: color_data = Z;
		19'b0100111010100010111: color_data = Z;
		19'b0100111010100011000: color_data = Z;
		19'b0100111010100011001: color_data = Z;
		19'b0100111010100011010: color_data = Z;
		19'b0100111010100011011: color_data = Z;
		19'b0100111010100011100: color_data = Z;
		19'b0100111010100011101: color_data = Z;
		19'b0100111010100011110: color_data = Z;
		19'b0100111010100011111: color_data = Z;
		19'b0100111010100100000: color_data = Z;
		19'b0100111010100101001: color_data = Z;
		19'b0100111010100101010: color_data = Z;
		19'b0100111010100101011: color_data = Z;
		19'b0100111010100101100: color_data = Z;
		19'b0100111010100101101: color_data = Z;
		19'b0100111010100101110: color_data = Z;
		19'b0100111010100101111: color_data = Z;
		19'b0100111010100110000: color_data = Z;
		19'b0100111010100110001: color_data = Z;
		19'b0100111010100110010: color_data = Z;
		19'b0100111010100110011: color_data = Z;
		19'b0100111010100110100: color_data = Z;
		19'b0100111010100110101: color_data = Z;
		19'b0100111010100110110: color_data = Z;
		19'b0100111010100110111: color_data = Z;
		19'b0100111010100111000: color_data = Z;
		19'b0100111010100111001: color_data = Z;
		19'b0100111010100111010: color_data = Z;
		19'b0100111010100111011: color_data = Z;
		19'b0100111010100111100: color_data = Z;
		19'b0100111010100111101: color_data = Z;
		19'b0100111010100111110: color_data = Z;
		19'b0100111010100111111: color_data = Z;
		19'b0100111010101000000: color_data = Z;
		19'b0100111010101000001: color_data = Z;
		19'b0100111010101000010: color_data = Z;
		19'b0100111010101000011: color_data = Z;
		19'b0100111010101000100: color_data = Z;
		19'b0100111010101000101: color_data = Z;
		19'b0100111010101000110: color_data = Z;
		19'b0100111010101000111: color_data = Z;
		19'b0100111010101001000: color_data = Z;
		19'b0100111010101001001: color_data = Z;
		19'b0100111010101001010: color_data = Z;
		19'b0100111010101001011: color_data = Z;
		19'b0100111010101001100: color_data = Z;
		19'b0100111010101001101: color_data = Z;
		19'b0100111010101001110: color_data = Z;
		19'b0100111010101001111: color_data = Z;
		19'b0100111010101010000: color_data = Z;
		19'b0100111010101010001: color_data = Z;
		19'b0100111010101010010: color_data = Z;
		19'b0100111010101010011: color_data = Z;
		19'b0100111010101010100: color_data = Z;
		19'b0100111010101010101: color_data = Z;
		19'b0100111010101010110: color_data = Z;
		19'b0100111010101010111: color_data = Z;
		19'b0100111010101011000: color_data = Z;
		19'b0100111010101011001: color_data = Z;
		19'b0100111010101011010: color_data = Z;
		19'b0100111010101011011: color_data = Z;
		19'b0100111010101011100: color_data = Z;
		19'b0100111010101011101: color_data = Z;
		19'b0100111010101011110: color_data = Z;
		19'b0100111010101011111: color_data = Z;
		19'b0100111010101100000: color_data = Z;
		19'b0100111010101100001: color_data = Z;
		19'b0100111010101100010: color_data = Z;
		19'b0100111010101100011: color_data = Z;
		19'b0100111010101100100: color_data = Z;
		19'b0100111010101100101: color_data = Z;
		19'b0100111010101100110: color_data = Z;
		19'b0100111010101100111: color_data = Z;
		19'b0100111010101101000: color_data = Z;
		19'b0100111010101101001: color_data = Z;
		19'b0100111010101101010: color_data = Z;
		19'b0100111010101101011: color_data = Z;
		19'b0100111010101101100: color_data = Z;
		19'b0100111010101101101: color_data = Z;
		19'b0100111010101101110: color_data = Z;
		19'b0100111010101101111: color_data = Z;
		19'b0100111010101110000: color_data = Z;
		19'b0100111010101110001: color_data = Z;
		19'b0100111010101110010: color_data = Z;
		19'b0100111010101110011: color_data = Z;
		19'b0100111010101110100: color_data = Z;
		19'b0100111010101110101: color_data = Z;
		19'b0100111010101110110: color_data = Z;
		19'b0100111010101110111: color_data = Z;
		19'b0100111010101111000: color_data = Z;
		19'b0100111010101111001: color_data = Z;
		19'b0100111010101111010: color_data = Z;
		19'b0100111010101111011: color_data = Z;
		19'b0100111010101111100: color_data = Z;
		19'b0100111010101111101: color_data = Z;
		19'b0100111010101111110: color_data = Z;
		19'b0100111010101111111: color_data = Z;
		19'b0100111010110000000: color_data = Z;
		19'b0100111010111001110: color_data = Z;
		19'b0100111010111001111: color_data = Z;
		19'b0100111010111010000: color_data = Z;
		19'b0100111010111010001: color_data = Z;
		19'b0100111010111010010: color_data = Z;
		19'b0100111010111010011: color_data = Z;
		19'b0100111010111010100: color_data = Z;
		19'b0100111010111010101: color_data = Z;
		19'b0100111010111010110: color_data = Z;
		19'b0100111010111010111: color_data = Z;
		19'b0100111010111011000: color_data = Z;
		19'b0100111010111011001: color_data = Z;
		19'b0100111010111011010: color_data = Z;
		19'b0100111010111011011: color_data = Z;
		19'b0100111010111011100: color_data = Z;
		19'b0100111010111011101: color_data = Z;
		19'b0100111010111011110: color_data = Z;
		19'b0100111010111011111: color_data = Z;
		19'b0100111010111100000: color_data = Z;
		19'b0100111100100011000: color_data = Z;
		19'b0100111100100011001: color_data = Z;
		19'b0100111100100011010: color_data = Z;
		19'b0100111100100011011: color_data = Z;
		19'b0100111100100011100: color_data = Z;
		19'b0100111100100011101: color_data = Z;
		19'b0100111100100011110: color_data = Z;
		19'b0100111100100011111: color_data = Z;
		19'b0100111100100100000: color_data = Z;
		19'b0100111100100101001: color_data = Z;
		19'b0100111100100101010: color_data = Z;
		19'b0100111100100101011: color_data = Z;
		19'b0100111100100101100: color_data = Z;
		19'b0100111100100101101: color_data = Z;
		19'b0100111100100101110: color_data = Z;
		19'b0100111100100101111: color_data = Z;
		19'b0100111100100110000: color_data = Z;
		19'b0100111100100110001: color_data = Z;
		19'b0100111100100110010: color_data = Z;
		19'b0100111100100110011: color_data = Z;
		19'b0100111100100110100: color_data = Z;
		19'b0100111100100110101: color_data = Z;
		19'b0100111100100110110: color_data = Z;
		19'b0100111100100110111: color_data = Z;
		19'b0100111100100111000: color_data = Z;
		19'b0100111100100111001: color_data = Z;
		19'b0100111100100111010: color_data = Z;
		19'b0100111100100111011: color_data = Z;
		19'b0100111100100111100: color_data = Z;
		19'b0100111100100111101: color_data = Z;
		19'b0100111100100111110: color_data = Z;
		19'b0100111100100111111: color_data = Z;
		19'b0100111100101000000: color_data = Z;
		19'b0100111100101000001: color_data = Z;
		19'b0100111100101000010: color_data = Z;
		19'b0100111100101000011: color_data = Z;
		19'b0100111100101000100: color_data = Z;
		19'b0100111100101000101: color_data = Z;
		19'b0100111100101000110: color_data = Z;
		19'b0100111100101000111: color_data = Z;
		19'b0100111100101001000: color_data = Z;
		19'b0100111100101001001: color_data = Z;
		19'b0100111100101001010: color_data = Z;
		19'b0100111100101001011: color_data = Z;
		19'b0100111100101001100: color_data = Z;
		19'b0100111100101001101: color_data = Z;
		19'b0100111100101001110: color_data = Z;
		19'b0100111100101001111: color_data = Z;
		19'b0100111100101010000: color_data = Z;
		19'b0100111100101010001: color_data = Z;
		19'b0100111100101010010: color_data = Z;
		19'b0100111100101010011: color_data = Z;
		19'b0100111100101010100: color_data = Z;
		19'b0100111100101010101: color_data = Z;
		19'b0100111100101010110: color_data = Z;
		19'b0100111100101010111: color_data = Z;
		19'b0100111100101011000: color_data = Z;
		19'b0100111100101011001: color_data = Z;
		19'b0100111100101011010: color_data = Z;
		19'b0100111100101011011: color_data = Z;
		19'b0100111100101011100: color_data = Z;
		19'b0100111100101011101: color_data = Z;
		19'b0100111100101011110: color_data = Z;
		19'b0100111100101011111: color_data = Z;
		19'b0100111100101100000: color_data = Z;
		19'b0100111100101100001: color_data = Z;
		19'b0100111100101100010: color_data = Z;
		19'b0100111100101100011: color_data = Z;
		19'b0100111100101100100: color_data = Z;
		19'b0100111100101100101: color_data = Z;
		19'b0100111100101100110: color_data = Z;
		19'b0100111100101100111: color_data = Z;
		19'b0100111100101101000: color_data = Z;
		19'b0100111100101101001: color_data = Z;
		19'b0100111100101101010: color_data = Z;
		19'b0100111100101101011: color_data = Z;
		19'b0100111100101101100: color_data = Z;
		19'b0100111100101101101: color_data = Z;
		19'b0100111100101101110: color_data = Z;
		19'b0100111100101101111: color_data = Z;
		19'b0100111100101110000: color_data = Z;
		19'b0100111100101110001: color_data = Z;
		19'b0100111100101110010: color_data = Z;
		19'b0100111100101110011: color_data = Z;
		19'b0100111100101110100: color_data = Z;
		19'b0100111100101110101: color_data = Z;
		19'b0100111100101110110: color_data = Z;
		19'b0100111100101110111: color_data = Z;
		19'b0100111100101111000: color_data = Z;
		19'b0100111100101111001: color_data = Z;
		19'b0100111100101111010: color_data = Z;
		19'b0100111100101111011: color_data = Z;
		19'b0100111100101111100: color_data = Z;
		19'b0100111100101111101: color_data = Z;
		19'b0100111100101111110: color_data = Z;
		19'b0100111100101111111: color_data = Z;
		19'b0100111100110000000: color_data = Z;
		19'b0100111100111001110: color_data = Z;
		19'b0100111100111001111: color_data = Z;
		19'b0100111100111010000: color_data = Z;
		19'b0100111100111010001: color_data = Z;
		19'b0100111100111010010: color_data = Z;
		19'b0100111100111010011: color_data = Z;
		19'b0100111100111010100: color_data = Z;
		19'b0100111100111010101: color_data = Z;
		19'b0100111100111010110: color_data = Z;
		19'b0100111100111010111: color_data = Z;
		19'b0100111100111011000: color_data = Z;
		19'b0100111100111011001: color_data = Z;
		19'b0100111100111011010: color_data = Z;
		19'b0100111100111011011: color_data = Z;
		19'b0100111100111011100: color_data = Z;
		19'b0100111100111011101: color_data = Z;
		19'b0100111100111011110: color_data = Z;
		19'b0100111100111011111: color_data = Z;
		19'b0100111110100011010: color_data = Z;
		19'b0100111110100011011: color_data = Z;
		19'b0100111110100011100: color_data = Z;
		19'b0100111110100011101: color_data = Z;
		19'b0100111110100011110: color_data = Z;
		19'b0100111110100011111: color_data = Z;
		19'b0100111110100100000: color_data = Z;
		19'b0100111110100101001: color_data = Z;
		19'b0100111110100101010: color_data = Z;
		19'b0100111110100101011: color_data = Z;
		19'b0100111110100101100: color_data = Z;
		19'b0100111110100101101: color_data = Z;
		19'b0100111110100101110: color_data = Z;
		19'b0100111110100101111: color_data = Z;
		19'b0100111110100110000: color_data = Z;
		19'b0100111110100110001: color_data = Z;
		19'b0100111110100110010: color_data = Z;
		19'b0100111110100110011: color_data = Z;
		19'b0100111110100110100: color_data = Z;
		19'b0100111110100110101: color_data = Z;
		19'b0100111110100110110: color_data = Z;
		19'b0100111110100110111: color_data = Z;
		19'b0100111110100111000: color_data = Z;
		19'b0100111110100111001: color_data = Z;
		19'b0100111110100111010: color_data = Z;
		19'b0100111110100111011: color_data = Z;
		19'b0100111110100111100: color_data = Z;
		19'b0100111110100111101: color_data = Z;
		19'b0100111110100111110: color_data = Z;
		19'b0100111110100111111: color_data = Z;
		19'b0100111110101000000: color_data = Z;
		19'b0100111110101000001: color_data = Z;
		19'b0100111110101000010: color_data = Z;
		19'b0100111110101000011: color_data = Z;
		19'b0100111110101000100: color_data = Z;
		19'b0100111110101000101: color_data = Z;
		19'b0100111110101000110: color_data = Z;
		19'b0100111110101000111: color_data = Z;
		19'b0100111110101001000: color_data = Z;
		19'b0100111110101001001: color_data = Z;
		19'b0100111110101001010: color_data = Z;
		19'b0100111110101001011: color_data = Z;
		19'b0100111110101001100: color_data = Z;
		19'b0100111110101001101: color_data = Z;
		19'b0100111110101001110: color_data = Z;
		19'b0100111110101001111: color_data = Z;
		19'b0100111110101010000: color_data = Z;
		19'b0100111110101010001: color_data = Z;
		19'b0100111110101010010: color_data = Z;
		19'b0100111110101010011: color_data = Z;
		19'b0100111110101010100: color_data = Z;
		19'b0100111110101010101: color_data = Z;
		19'b0100111110101010110: color_data = Z;
		19'b0100111110101010111: color_data = Z;
		19'b0100111110101011000: color_data = Z;
		19'b0100111110101011001: color_data = Z;
		19'b0100111110101011010: color_data = Z;
		19'b0100111110101011011: color_data = Z;
		19'b0100111110101011100: color_data = Z;
		19'b0100111110101011101: color_data = Z;
		19'b0100111110101011110: color_data = Z;
		19'b0100111110101011111: color_data = Z;
		19'b0100111110101100000: color_data = Z;
		19'b0100111110101100001: color_data = Z;
		19'b0100111110101100010: color_data = Z;
		19'b0100111110101100011: color_data = Z;
		19'b0100111110101100100: color_data = Z;
		19'b0100111110101100101: color_data = Z;
		19'b0100111110101100110: color_data = Z;
		19'b0100111110101100111: color_data = Z;
		19'b0100111110101101000: color_data = Z;
		19'b0100111110101101001: color_data = Z;
		19'b0100111110101101010: color_data = Z;
		19'b0100111110101101011: color_data = Z;
		19'b0100111110101101100: color_data = Z;
		19'b0100111110101101101: color_data = Z;
		19'b0100111110101101110: color_data = Z;
		19'b0100111110101101111: color_data = Z;
		19'b0100111110101110000: color_data = Z;
		19'b0100111110101110001: color_data = Z;
		19'b0100111110101110010: color_data = Z;
		19'b0100111110101110011: color_data = Z;
		19'b0100111110101110100: color_data = Z;
		19'b0100111110101110101: color_data = Z;
		19'b0100111110101110110: color_data = Z;
		19'b0100111110101110111: color_data = Z;
		19'b0100111110101111000: color_data = Z;
		19'b0100111110101111001: color_data = Z;
		19'b0100111110101111010: color_data = Z;
		19'b0100111110101111011: color_data = Z;
		19'b0100111110101111100: color_data = Z;
		19'b0100111110101111101: color_data = Z;
		19'b0100111110101111110: color_data = Z;
		19'b0100111110101111111: color_data = Z;
		19'b0100111110110000000: color_data = Z;
		19'b0100111110111001110: color_data = Z;
		19'b0100111110111001111: color_data = Z;
		19'b0100111110111010000: color_data = Z;
		19'b0100111110111010001: color_data = Z;
		19'b0100111110111010010: color_data = Z;
		19'b0100111110111010011: color_data = Z;
		19'b0100111110111010100: color_data = Z;
		19'b0100111110111010101: color_data = Z;
		19'b0100111110111010110: color_data = Z;
		19'b0100111110111010111: color_data = Z;
		19'b0100111110111011000: color_data = Z;
		19'b0100111110111011001: color_data = Z;
		19'b0100111110111011010: color_data = Z;
		19'b0100111110111011011: color_data = Z;
		19'b0100111110111011100: color_data = Z;
		19'b0100111110111011101: color_data = Z;
		19'b0100111110111011110: color_data = Z;
		19'b0100111110111011111: color_data = Z;
		19'b0101000000100011010: color_data = Z;
		19'b0101000000100011011: color_data = Z;
		19'b0101000000100011100: color_data = Z;
		19'b0101000000100011101: color_data = Z;
		19'b0101000000100011110: color_data = Z;
		19'b0101000000100011111: color_data = Z;
		19'b0101000000100100000: color_data = Z;
		19'b0101000000100100001: color_data = Z;
		19'b0101000000100101010: color_data = Z;
		19'b0101000000100101011: color_data = Z;
		19'b0101000000100101100: color_data = Z;
		19'b0101000000100101101: color_data = Z;
		19'b0101000000100101110: color_data = Z;
		19'b0101000000100101111: color_data = Z;
		19'b0101000000100110000: color_data = Z;
		19'b0101000000100110001: color_data = Z;
		19'b0101000000100110010: color_data = Z;
		19'b0101000000100110011: color_data = Z;
		19'b0101000000100110100: color_data = Z;
		19'b0101000000100110101: color_data = Z;
		19'b0101000000100110110: color_data = Z;
		19'b0101000000100110111: color_data = Z;
		19'b0101000000100111000: color_data = Z;
		19'b0101000000100111001: color_data = Z;
		19'b0101000000100111010: color_data = Z;
		19'b0101000000100111011: color_data = Z;
		19'b0101000000100111100: color_data = Z;
		19'b0101000000100111101: color_data = Z;
		19'b0101000000100111110: color_data = Z;
		19'b0101000000100111111: color_data = Z;
		19'b0101000000101000000: color_data = Z;
		19'b0101000000101000001: color_data = Z;
		19'b0101000000101000010: color_data = Z;
		19'b0101000000101000011: color_data = Z;
		19'b0101000000101000100: color_data = Z;
		19'b0101000000101000101: color_data = Z;
		19'b0101000000101000110: color_data = Z;
		19'b0101000000101000111: color_data = Z;
		19'b0101000000101001000: color_data = Z;
		19'b0101000000101001001: color_data = Z;
		19'b0101000000101001010: color_data = Z;
		19'b0101000000101001011: color_data = Z;
		19'b0101000000101001100: color_data = Z;
		19'b0101000000101001101: color_data = Z;
		19'b0101000000101001110: color_data = Z;
		19'b0101000000101001111: color_data = Z;
		19'b0101000000101010000: color_data = Z;
		19'b0101000000101010001: color_data = Z;
		19'b0101000000101010010: color_data = Z;
		19'b0101000000101010011: color_data = Z;
		19'b0101000000101010100: color_data = Z;
		19'b0101000000101010101: color_data = Z;
		19'b0101000000101010110: color_data = Z;
		19'b0101000000101010111: color_data = Z;
		19'b0101000000101011000: color_data = Z;
		19'b0101000000101011001: color_data = Z;
		19'b0101000000101011010: color_data = Z;
		19'b0101000000101011011: color_data = Z;
		19'b0101000000101011100: color_data = Z;
		19'b0101000000101011101: color_data = Z;
		19'b0101000000101011110: color_data = Z;
		19'b0101000000101011111: color_data = Z;
		19'b0101000000101100000: color_data = Z;
		19'b0101000000101100001: color_data = Z;
		19'b0101000000101100010: color_data = Z;
		19'b0101000000101100011: color_data = Z;
		19'b0101000000101100100: color_data = Z;
		19'b0101000000101100101: color_data = Z;
		19'b0101000000101100110: color_data = Z;
		19'b0101000000101100111: color_data = Z;
		19'b0101000000101101000: color_data = Z;
		19'b0101000000101101001: color_data = Z;
		19'b0101000000101101010: color_data = Z;
		19'b0101000000101101011: color_data = Z;
		19'b0101000000101101100: color_data = Z;
		19'b0101000000101101101: color_data = Z;
		19'b0101000000101101110: color_data = Z;
		19'b0101000000101101111: color_data = Z;
		19'b0101000000101110000: color_data = Z;
		19'b0101000000101110001: color_data = Z;
		19'b0101000000101110010: color_data = Z;
		19'b0101000000101110011: color_data = Z;
		19'b0101000000101110100: color_data = Z;
		19'b0101000000101110101: color_data = Z;
		19'b0101000000101110110: color_data = Z;
		19'b0101000000101110111: color_data = Z;
		19'b0101000000101111000: color_data = Z;
		19'b0101000000101111001: color_data = Z;
		19'b0101000000101111010: color_data = Z;
		19'b0101000000101111011: color_data = Z;
		19'b0101000000101111100: color_data = Z;
		19'b0101000000101111101: color_data = Z;
		19'b0101000000101111110: color_data = Z;
		19'b0101000000101111111: color_data = Z;
		19'b0101000000110000000: color_data = Z;
		19'b0101000000111001110: color_data = Z;
		19'b0101000000111001111: color_data = Z;
		19'b0101000000111010000: color_data = Z;
		19'b0101000000111010001: color_data = Z;
		19'b0101000000111010010: color_data = Z;
		19'b0101000000111010011: color_data = Z;
		19'b0101000000111010100: color_data = Z;
		19'b0101000000111010110: color_data = Z;
		19'b0101000000111010111: color_data = Z;
		19'b0101000000111011000: color_data = Z;
		19'b0101000000111011001: color_data = Z;
		19'b0101000000111011010: color_data = Z;
		19'b0101000000111011011: color_data = Z;
		19'b0101000000111011100: color_data = Z;
		19'b0101000000111011101: color_data = Z;
		19'b0101000000111011110: color_data = Z;
		19'b0101000000111100001: color_data = Z;
		19'b0101000010100011011: color_data = Z;
		19'b0101000010100011100: color_data = Z;
		19'b0101000010100011101: color_data = Z;
		19'b0101000010100011110: color_data = Z;
		19'b0101000010100011111: color_data = Z;
		19'b0101000010100100000: color_data = Z;
		19'b0101000010100100001: color_data = Z;
		19'b0101000010100101010: color_data = Z;
		19'b0101000010100101011: color_data = Z;
		19'b0101000010100101100: color_data = Z;
		19'b0101000010100101101: color_data = Z;
		19'b0101000010100101110: color_data = Z;
		19'b0101000010100101111: color_data = Z;
		19'b0101000010100110000: color_data = Z;
		19'b0101000010100110001: color_data = Z;
		19'b0101000010100110010: color_data = Z;
		19'b0101000010100110011: color_data = Z;
		19'b0101000010100110100: color_data = Z;
		19'b0101000010100110101: color_data = Z;
		19'b0101000010100110110: color_data = Z;
		19'b0101000010100110111: color_data = Z;
		19'b0101000010100111000: color_data = Z;
		19'b0101000010100111001: color_data = Z;
		19'b0101000010100111010: color_data = Z;
		19'b0101000010100111011: color_data = Z;
		19'b0101000010100111100: color_data = Z;
		19'b0101000010100111101: color_data = Z;
		19'b0101000010100111110: color_data = Z;
		19'b0101000010100111111: color_data = Z;
		19'b0101000010101000000: color_data = Z;
		19'b0101000010101000001: color_data = Z;
		19'b0101000010101000010: color_data = Z;
		19'b0101000010101000011: color_data = Z;
		19'b0101000010101000100: color_data = Z;
		19'b0101000010101000101: color_data = Z;
		19'b0101000010101000110: color_data = Z;
		19'b0101000010101000111: color_data = Z;
		19'b0101000010101001000: color_data = Z;
		19'b0101000010101001001: color_data = Z;
		19'b0101000010101001010: color_data = Z;
		19'b0101000010101001011: color_data = Z;
		19'b0101000010101001100: color_data = Z;
		19'b0101000010101001101: color_data = Z;
		19'b0101000010101001110: color_data = Z;
		19'b0101000010101001111: color_data = Z;
		19'b0101000010101010000: color_data = Z;
		19'b0101000010101010001: color_data = Z;
		19'b0101000010101010010: color_data = Z;
		19'b0101000010101010011: color_data = Z;
		19'b0101000010101010100: color_data = Z;
		19'b0101000010101010101: color_data = Z;
		19'b0101000010101010110: color_data = Z;
		19'b0101000010101010111: color_data = Z;
		19'b0101000010101011000: color_data = Z;
		19'b0101000010101011001: color_data = Z;
		19'b0101000010101011010: color_data = Z;
		19'b0101000010101011011: color_data = Z;
		19'b0101000010101011100: color_data = Z;
		19'b0101000010101011101: color_data = Z;
		19'b0101000010101011110: color_data = Z;
		19'b0101000010101011111: color_data = Z;
		19'b0101000010101100000: color_data = Z;
		19'b0101000010101100001: color_data = Z;
		19'b0101000010101100010: color_data = Z;
		19'b0101000010101100011: color_data = Z;
		19'b0101000010101100100: color_data = Z;
		19'b0101000010101100101: color_data = Z;
		19'b0101000010101100110: color_data = Z;
		19'b0101000010101100111: color_data = Z;
		19'b0101000010101101000: color_data = Z;
		19'b0101000010101101001: color_data = Z;
		19'b0101000010101101010: color_data = Z;
		19'b0101000010101101011: color_data = Z;
		19'b0101000010101101100: color_data = Z;
		19'b0101000010101101101: color_data = Z;
		19'b0101000010101101110: color_data = Z;
		19'b0101000010101101111: color_data = Z;
		19'b0101000010101110000: color_data = Z;
		19'b0101000010101110001: color_data = Z;
		19'b0101000010101110010: color_data = Z;
		19'b0101000010101110011: color_data = Z;
		19'b0101000010101110100: color_data = Z;
		19'b0101000010101110101: color_data = Z;
		19'b0101000010101110110: color_data = Z;
		19'b0101000010101110111: color_data = Z;
		19'b0101000010101111000: color_data = Z;
		19'b0101000010101111001: color_data = Z;
		19'b0101000010101111010: color_data = Z;
		19'b0101000010101111011: color_data = Z;
		19'b0101000010101111100: color_data = Z;
		19'b0101000010101111101: color_data = Z;
		19'b0101000010101111110: color_data = Z;
		19'b0101000010101111111: color_data = Z;
		19'b0101000010110000000: color_data = Z;
		19'b0101000010111001111: color_data = Z;
		19'b0101000010111010000: color_data = Z;
		19'b0101000010111010001: color_data = Z;
		19'b0101000010111010010: color_data = Z;
		19'b0101000010111010011: color_data = Z;
		19'b0101000010111010100: color_data = Z;
		19'b0101000010111010110: color_data = Z;
		19'b0101000010111010111: color_data = Z;
		19'b0101000010111011000: color_data = Z;
		19'b0101000010111011001: color_data = Z;
		19'b0101000010111011010: color_data = Z;
		19'b0101000010111011011: color_data = Z;
		19'b0101000010111011100: color_data = Z;
		19'b0101000010111011101: color_data = Z;
		19'b0101000010111011110: color_data = Z;
		19'b0101000010111100001: color_data = Z;
		19'b0101000100100011100: color_data = Z;
		19'b0101000100100011101: color_data = Z;
		19'b0101000100100011110: color_data = Z;
		19'b0101000100100011111: color_data = Z;
		19'b0101000100100100000: color_data = Z;
		19'b0101000100100100001: color_data = Z;
		19'b0101000100100101010: color_data = Z;
		19'b0101000100100101011: color_data = Z;
		19'b0101000100100101100: color_data = Z;
		19'b0101000100100101101: color_data = Z;
		19'b0101000100100101110: color_data = Z;
		19'b0101000100100101111: color_data = Z;
		19'b0101000100100110000: color_data = Z;
		19'b0101000100100110001: color_data = Z;
		19'b0101000100100110010: color_data = Z;
		19'b0101000100100110011: color_data = Z;
		19'b0101000100100110100: color_data = Z;
		19'b0101000100100110101: color_data = Z;
		19'b0101000100100110110: color_data = Z;
		19'b0101000100100110111: color_data = Z;
		19'b0101000100100111000: color_data = Z;
		19'b0101000100100111001: color_data = Z;
		19'b0101000100100111010: color_data = Z;
		19'b0101000100100111011: color_data = Z;
		19'b0101000100100111100: color_data = Z;
		19'b0101000100100111101: color_data = Z;
		19'b0101000100100111110: color_data = Z;
		19'b0101000100100111111: color_data = Z;
		19'b0101000100101000000: color_data = Z;
		19'b0101000100101000001: color_data = Z;
		19'b0101000100101000010: color_data = Z;
		19'b0101000100101000011: color_data = Z;
		19'b0101000100101000100: color_data = Z;
		19'b0101000100101000101: color_data = Z;
		19'b0101000100101000110: color_data = Z;
		19'b0101000100101000111: color_data = Z;
		19'b0101000100101001000: color_data = Z;
		19'b0101000100101001001: color_data = Z;
		19'b0101000100101001010: color_data = Z;
		19'b0101000100101001011: color_data = Z;
		19'b0101000100101001100: color_data = Z;
		19'b0101000100101001101: color_data = Z;
		19'b0101000100101001110: color_data = Z;
		19'b0101000100101001111: color_data = Z;
		19'b0101000100101010000: color_data = Z;
		19'b0101000100101010001: color_data = Z;
		19'b0101000100101010010: color_data = Z;
		19'b0101000100101010011: color_data = Z;
		19'b0101000100101010100: color_data = Z;
		19'b0101000100101010101: color_data = Z;
		19'b0101000100101010110: color_data = Z;
		19'b0101000100101010111: color_data = Z;
		19'b0101000100101011000: color_data = Z;
		19'b0101000100101011001: color_data = Z;
		19'b0101000100101011010: color_data = Z;
		19'b0101000100101011011: color_data = Z;
		19'b0101000100101011100: color_data = Z;
		19'b0101000100101011101: color_data = Z;
		19'b0101000100101011110: color_data = Z;
		19'b0101000100101011111: color_data = Z;
		19'b0101000100101100000: color_data = Z;
		19'b0101000100101100001: color_data = Z;
		19'b0101000100101100010: color_data = Z;
		19'b0101000100101100011: color_data = Z;
		19'b0101000100101100100: color_data = Z;
		19'b0101000100101100101: color_data = Z;
		19'b0101000100101100110: color_data = Z;
		19'b0101000100101100111: color_data = Z;
		19'b0101000100101101000: color_data = Z;
		19'b0101000100101101001: color_data = Z;
		19'b0101000100101101010: color_data = Z;
		19'b0101000100101101011: color_data = Z;
		19'b0101000100101101100: color_data = Z;
		19'b0101000100101101101: color_data = Z;
		19'b0101000100101101110: color_data = Z;
		19'b0101000100101101111: color_data = Z;
		19'b0101000100101110000: color_data = Z;
		19'b0101000100101110001: color_data = Z;
		19'b0101000100101110010: color_data = Z;
		19'b0101000100101110011: color_data = Z;
		19'b0101000100101110100: color_data = Z;
		19'b0101000100101110101: color_data = Z;
		19'b0101000100101110110: color_data = Z;
		19'b0101000100101110111: color_data = Z;
		19'b0101000100101111000: color_data = Z;
		19'b0101000100101111001: color_data = Z;
		19'b0101000100101111010: color_data = Z;
		19'b0101000100101111011: color_data = Z;
		19'b0101000100101111100: color_data = Z;
		19'b0101000100101111101: color_data = Z;
		19'b0101000100101111110: color_data = Z;
		19'b0101000100101111111: color_data = Z;
		19'b0101000100110000000: color_data = Z;
		19'b0101000100111001111: color_data = Z;
		19'b0101000100111010000: color_data = Z;
		19'b0101000100111010001: color_data = Z;
		19'b0101000100111010010: color_data = Z;
		19'b0101000100111010011: color_data = Z;
		19'b0101000100111010110: color_data = Z;
		19'b0101000100111010111: color_data = Z;
		19'b0101000100111011000: color_data = Z;
		19'b0101000100111011001: color_data = Z;
		19'b0101000100111011010: color_data = Z;
		19'b0101000100111011011: color_data = Z;
		19'b0101000100111011100: color_data = Z;
		19'b0101000110100011101: color_data = Z;
		19'b0101000110100011110: color_data = Z;
		19'b0101000110100011111: color_data = Z;
		19'b0101000110100100000: color_data = Z;
		19'b0101000110100100001: color_data = Z;
		19'b0101000110100100010: color_data = Z;
		19'b0101000110100101010: color_data = Z;
		19'b0101000110100101011: color_data = Z;
		19'b0101000110100101100: color_data = Z;
		19'b0101000110100101101: color_data = Z;
		19'b0101000110100101110: color_data = Z;
		19'b0101000110100101111: color_data = Z;
		19'b0101000110100110000: color_data = Z;
		19'b0101000110100110001: color_data = Z;
		19'b0101000110100110010: color_data = Z;
		19'b0101000110100110011: color_data = Z;
		19'b0101000110100110100: color_data = Z;
		19'b0101000110100110101: color_data = Z;
		19'b0101000110100110110: color_data = Z;
		19'b0101000110100110111: color_data = Z;
		19'b0101000110100111000: color_data = Z;
		19'b0101000110100111001: color_data = Z;
		19'b0101000110100111010: color_data = Z;
		19'b0101000110100111011: color_data = Z;
		19'b0101000110100111100: color_data = Z;
		19'b0101000110100111101: color_data = Z;
		19'b0101000110100111110: color_data = Z;
		19'b0101000110100111111: color_data = Z;
		19'b0101000110101000000: color_data = Z;
		19'b0101000110101000001: color_data = Z;
		19'b0101000110101000010: color_data = Z;
		19'b0101000110101000011: color_data = Z;
		19'b0101000110101000100: color_data = Z;
		19'b0101000110101000101: color_data = Z;
		19'b0101000110101000110: color_data = Z;
		19'b0101000110101000111: color_data = Z;
		19'b0101000110101001000: color_data = Z;
		19'b0101000110101001001: color_data = Z;
		19'b0101000110101001010: color_data = Z;
		19'b0101000110101001011: color_data = Z;
		19'b0101000110101001100: color_data = Z;
		19'b0101000110101001101: color_data = Z;
		19'b0101000110101001110: color_data = Z;
		19'b0101000110101001111: color_data = Z;
		19'b0101000110101010000: color_data = Z;
		19'b0101000110101010001: color_data = Z;
		19'b0101000110101010010: color_data = Z;
		19'b0101000110101010011: color_data = Z;
		19'b0101000110101010100: color_data = Z;
		19'b0101000110101010101: color_data = Z;
		19'b0101000110101010110: color_data = Z;
		19'b0101000110101010111: color_data = Z;
		19'b0101000110101011000: color_data = Z;
		19'b0101000110101011001: color_data = Z;
		19'b0101000110101011010: color_data = Z;
		19'b0101000110101011011: color_data = Z;
		19'b0101000110101011100: color_data = Z;
		19'b0101000110101011101: color_data = Z;
		19'b0101000110101011110: color_data = Z;
		19'b0101000110101011111: color_data = Z;
		19'b0101000110101100000: color_data = Z;
		19'b0101000110101100001: color_data = Z;
		19'b0101000110101100010: color_data = Z;
		19'b0101000110101100011: color_data = Z;
		19'b0101000110101100100: color_data = Z;
		19'b0101000110101100101: color_data = Z;
		19'b0101000110101100110: color_data = Z;
		19'b0101000110101100111: color_data = Z;
		19'b0101000110101101000: color_data = Z;
		19'b0101000110101101001: color_data = Z;
		19'b0101000110101101010: color_data = Z;
		19'b0101000110101101011: color_data = Z;
		19'b0101000110101101100: color_data = Z;
		19'b0101000110101101101: color_data = Z;
		19'b0101000110101101110: color_data = Z;
		19'b0101000110101101111: color_data = Z;
		19'b0101000110101110000: color_data = Z;
		19'b0101000110101110001: color_data = Z;
		19'b0101000110101110010: color_data = Z;
		19'b0101000110101110011: color_data = Z;
		19'b0101000110101110100: color_data = Z;
		19'b0101000110101110101: color_data = Z;
		19'b0101000110101110110: color_data = Z;
		19'b0101000110101110111: color_data = Z;
		19'b0101000110101111000: color_data = Z;
		19'b0101000110101111001: color_data = Z;
		19'b0101000110101111010: color_data = Z;
		19'b0101000110101111011: color_data = Z;
		19'b0101000110101111100: color_data = Z;
		19'b0101000110101111101: color_data = Z;
		19'b0101000110101111110: color_data = Z;
		19'b0101000110101111111: color_data = Z;
		19'b0101000110110000000: color_data = Z;
		19'b0101000110111001111: color_data = Z;
		19'b0101000110111010000: color_data = Z;
		19'b0101000110111010001: color_data = Z;
		19'b0101000110111010010: color_data = Z;
		19'b0101000110111010011: color_data = Z;
		19'b0101000110111010110: color_data = Z;
		19'b0101000110111010111: color_data = Z;
		19'b0101000110111011000: color_data = Z;
		19'b0101000110111011001: color_data = Z;
		19'b0101000110111011010: color_data = Z;
		19'b0101000110111011011: color_data = Z;
		19'b0101000110111011100: color_data = Z;
		19'b0101001000100011101: color_data = Z;
		19'b0101001000100011110: color_data = Z;
		19'b0101001000100011111: color_data = Z;
		19'b0101001000100100000: color_data = Z;
		19'b0101001000100100001: color_data = Z;
		19'b0101001000100100010: color_data = Z;
		19'b0101001000100100011: color_data = Z;
		19'b0101001000100100100: color_data = Z;
		19'b0101001000100101010: color_data = Z;
		19'b0101001000100101011: color_data = Z;
		19'b0101001000100101100: color_data = Z;
		19'b0101001000100101101: color_data = Z;
		19'b0101001000100101110: color_data = Z;
		19'b0101001000100101111: color_data = Z;
		19'b0101001000100110000: color_data = Z;
		19'b0101001000100110001: color_data = Z;
		19'b0101001000100110010: color_data = Z;
		19'b0101001000100110011: color_data = Z;
		19'b0101001000100110100: color_data = Z;
		19'b0101001000100110101: color_data = Z;
		19'b0101001000100110110: color_data = Z;
		19'b0101001000100110111: color_data = Z;
		19'b0101001000100111000: color_data = Z;
		19'b0101001000100111001: color_data = Z;
		19'b0101001000100111010: color_data = Z;
		19'b0101001000100111011: color_data = Z;
		19'b0101001000100111100: color_data = Z;
		19'b0101001000100111101: color_data = Z;
		19'b0101001000100111110: color_data = Z;
		19'b0101001000100111111: color_data = Z;
		19'b0101001000101000000: color_data = Z;
		19'b0101001000101000001: color_data = Z;
		19'b0101001000101000010: color_data = Z;
		19'b0101001000101000011: color_data = Z;
		19'b0101001000101000100: color_data = Z;
		19'b0101001000101000101: color_data = Z;
		19'b0101001000101000110: color_data = Z;
		19'b0101001000101000111: color_data = Z;
		19'b0101001000101001000: color_data = Z;
		19'b0101001000101001001: color_data = Z;
		19'b0101001000101001010: color_data = Z;
		19'b0101001000101001011: color_data = Z;
		19'b0101001000101001100: color_data = Z;
		19'b0101001000101001101: color_data = Z;
		19'b0101001000101001110: color_data = Z;
		19'b0101001000101001111: color_data = Z;
		19'b0101001000101010000: color_data = Z;
		19'b0101001000101010001: color_data = Z;
		19'b0101001000101010010: color_data = Z;
		19'b0101001000101010011: color_data = Z;
		19'b0101001000101010100: color_data = Z;
		19'b0101001000101010101: color_data = Z;
		19'b0101001000101010110: color_data = Z;
		19'b0101001000101010111: color_data = Z;
		19'b0101001000101011000: color_data = Z;
		19'b0101001000101011001: color_data = Z;
		19'b0101001000101011010: color_data = Z;
		19'b0101001000101011011: color_data = Z;
		19'b0101001000101011100: color_data = Z;
		19'b0101001000101011101: color_data = Z;
		19'b0101001000101011110: color_data = Z;
		19'b0101001000101011111: color_data = Z;
		19'b0101001000101100000: color_data = Z;
		19'b0101001000101100001: color_data = Z;
		19'b0101001000101100010: color_data = Z;
		19'b0101001000101100011: color_data = Z;
		19'b0101001000101100100: color_data = Z;
		19'b0101001000101100101: color_data = Z;
		19'b0101001000101100110: color_data = Z;
		19'b0101001000101100111: color_data = Z;
		19'b0101001000101101000: color_data = Z;
		19'b0101001000101101001: color_data = Z;
		19'b0101001000101101010: color_data = Z;
		19'b0101001000101101011: color_data = Z;
		19'b0101001000101101100: color_data = Z;
		19'b0101001000101101101: color_data = Z;
		19'b0101001000101101110: color_data = Z;
		19'b0101001000101101111: color_data = Z;
		19'b0101001000101110000: color_data = Z;
		19'b0101001000101110001: color_data = Z;
		19'b0101001000101110010: color_data = Z;
		19'b0101001000101110011: color_data = Z;
		19'b0101001000101110100: color_data = Z;
		19'b0101001000101110101: color_data = Z;
		19'b0101001000101110110: color_data = Z;
		19'b0101001000101110111: color_data = Z;
		19'b0101001000101111000: color_data = Z;
		19'b0101001000101111001: color_data = Z;
		19'b0101001000101111010: color_data = Z;
		19'b0101001000101111011: color_data = Z;
		19'b0101001000101111100: color_data = Z;
		19'b0101001000101111101: color_data = Z;
		19'b0101001000101111110: color_data = Z;
		19'b0101001000101111111: color_data = Z;
		19'b0101001000110000000: color_data = Z;
		19'b0101001000111001111: color_data = Z;
		19'b0101001000111010000: color_data = Z;
		19'b0101001000111010001: color_data = Z;
		19'b0101001000111010010: color_data = Z;
		19'b0101001000111010011: color_data = Z;
		19'b0101001000111010100: color_data = Z;
		19'b0101001000111010110: color_data = Z;
		19'b0101001000111010111: color_data = Z;
		19'b0101001000111011000: color_data = Z;
		19'b0101001000111011001: color_data = Z;
		19'b0101001000111011010: color_data = Z;
		19'b0101001000111011011: color_data = Z;
		19'b0101001000111011100: color_data = Z;
		19'b0101001000111011101: color_data = Z;
		19'b0101001000111100000: color_data = Z;
		19'b0101001010100011110: color_data = Z;
		19'b0101001010100011111: color_data = Z;
		19'b0101001010100100000: color_data = Z;
		19'b0101001010100100001: color_data = Z;
		19'b0101001010100100010: color_data = Z;
		19'b0101001010100100011: color_data = Z;
		19'b0101001010100100100: color_data = Z;
		19'b0101001010100101010: color_data = Z;
		19'b0101001010100101011: color_data = Z;
		19'b0101001010100101100: color_data = Z;
		19'b0101001010100101101: color_data = Z;
		19'b0101001010100101110: color_data = Z;
		19'b0101001010100101111: color_data = Z;
		19'b0101001010100110000: color_data = Z;
		19'b0101001010100110001: color_data = Z;
		19'b0101001010100110010: color_data = Z;
		19'b0101001010100110011: color_data = Z;
		19'b0101001010100110100: color_data = Z;
		19'b0101001010100110101: color_data = Z;
		19'b0101001010100110110: color_data = Z;
		19'b0101001010100110111: color_data = Z;
		19'b0101001010100111000: color_data = Z;
		19'b0101001010100111001: color_data = Z;
		19'b0101001010100111010: color_data = Z;
		19'b0101001010100111011: color_data = Z;
		19'b0101001010100111100: color_data = Z;
		19'b0101001010100111101: color_data = Z;
		19'b0101001010100111110: color_data = Z;
		19'b0101001010100111111: color_data = Z;
		19'b0101001010101000000: color_data = Z;
		19'b0101001010101000001: color_data = Z;
		19'b0101001010101000010: color_data = Z;
		19'b0101001010101000011: color_data = Z;
		19'b0101001010101000100: color_data = Z;
		19'b0101001010101000101: color_data = Z;
		19'b0101001010101000110: color_data = Z;
		19'b0101001010101000111: color_data = Z;
		19'b0101001010101001000: color_data = Z;
		19'b0101001010101001001: color_data = Z;
		19'b0101001010101001010: color_data = Z;
		19'b0101001010101001011: color_data = Z;
		19'b0101001010101001100: color_data = Z;
		19'b0101001010101001101: color_data = Z;
		19'b0101001010101001110: color_data = Z;
		19'b0101001010101001111: color_data = Z;
		19'b0101001010101010000: color_data = Z;
		19'b0101001010101010001: color_data = Z;
		19'b0101001010101010010: color_data = Z;
		19'b0101001010101010011: color_data = Z;
		19'b0101001010101010100: color_data = Z;
		19'b0101001010101010101: color_data = Z;
		19'b0101001010101010110: color_data = Z;
		19'b0101001010101010111: color_data = Z;
		19'b0101001010101011000: color_data = Z;
		19'b0101001010101011001: color_data = Z;
		19'b0101001010101011010: color_data = Z;
		19'b0101001010101011011: color_data = Z;
		19'b0101001010101011100: color_data = Z;
		19'b0101001010101011101: color_data = Z;
		19'b0101001010101011110: color_data = Z;
		19'b0101001010101011111: color_data = Z;
		19'b0101001010101100000: color_data = Z;
		19'b0101001010101100001: color_data = Z;
		19'b0101001010101100010: color_data = Z;
		19'b0101001010101100011: color_data = Z;
		19'b0101001010101100100: color_data = Z;
		19'b0101001010101100101: color_data = Z;
		19'b0101001010101100110: color_data = Z;
		19'b0101001010101100111: color_data = Z;
		19'b0101001010101101000: color_data = Z;
		19'b0101001010101101001: color_data = Z;
		19'b0101001010101101010: color_data = Z;
		19'b0101001010101101011: color_data = Z;
		19'b0101001010101101100: color_data = Z;
		19'b0101001010101101101: color_data = Z;
		19'b0101001010101101110: color_data = Z;
		19'b0101001010101101111: color_data = Z;
		19'b0101001010101110000: color_data = Z;
		19'b0101001010101110001: color_data = Z;
		19'b0101001010101110010: color_data = Z;
		19'b0101001010101110011: color_data = Z;
		19'b0101001010101110100: color_data = Z;
		19'b0101001010101110101: color_data = Z;
		19'b0101001010101110110: color_data = Z;
		19'b0101001010101110111: color_data = Z;
		19'b0101001010101111000: color_data = Z;
		19'b0101001010101111001: color_data = Z;
		19'b0101001010101111010: color_data = Z;
		19'b0101001010101111011: color_data = Z;
		19'b0101001010101111100: color_data = Z;
		19'b0101001010101111101: color_data = Z;
		19'b0101001010101111110: color_data = Z;
		19'b0101001010101111111: color_data = Z;
		19'b0101001010110000000: color_data = Z;
		19'b0101001010111001111: color_data = Z;
		19'b0101001010111010000: color_data = Z;
		19'b0101001010111010001: color_data = Z;
		19'b0101001010111010010: color_data = Z;
		19'b0101001010111010011: color_data = Z;
		19'b0101001010111010100: color_data = Z;
		19'b0101001010111010110: color_data = Z;
		19'b0101001010111010111: color_data = Z;
		19'b0101001010111011000: color_data = Z;
		19'b0101001010111011001: color_data = Z;
		19'b0101001010111011010: color_data = Z;
		19'b0101001010111011011: color_data = Z;
		19'b0101001010111011100: color_data = Z;
		19'b0101001010111011101: color_data = Z;
		19'b0101001100100011110: color_data = Z;
		19'b0101001100100011111: color_data = Z;
		19'b0101001100100100000: color_data = Z;
		19'b0101001100100100001: color_data = Z;
		19'b0101001100100100010: color_data = Z;
		19'b0101001100100100011: color_data = Z;
		19'b0101001100100100100: color_data = Z;
		19'b0101001100100100101: color_data = Z;
		19'b0101001100100101010: color_data = Z;
		19'b0101001100100101011: color_data = Z;
		19'b0101001100100101100: color_data = Z;
		19'b0101001100100101101: color_data = Z;
		19'b0101001100100101110: color_data = Z;
		19'b0101001100100101111: color_data = Z;
		19'b0101001100100110000: color_data = Z;
		19'b0101001100100110001: color_data = Z;
		19'b0101001100100110010: color_data = Z;
		19'b0101001100100110011: color_data = Z;
		19'b0101001100100110100: color_data = Z;
		19'b0101001100100110101: color_data = Z;
		19'b0101001100100110110: color_data = Z;
		19'b0101001100100110111: color_data = Z;
		19'b0101001100100111000: color_data = Z;
		19'b0101001100100111001: color_data = Z;
		19'b0101001100100111010: color_data = Z;
		19'b0101001100100111011: color_data = Z;
		19'b0101001100100111100: color_data = Z;
		19'b0101001100100111101: color_data = Z;
		19'b0101001100100111110: color_data = Z;
		19'b0101001100100111111: color_data = Z;
		19'b0101001100101000000: color_data = Z;
		19'b0101001100101000001: color_data = Z;
		19'b0101001100101000010: color_data = Z;
		19'b0101001100101000011: color_data = Z;
		19'b0101001100101000100: color_data = Z;
		19'b0101001100101000101: color_data = Z;
		19'b0101001100101000110: color_data = Z;
		19'b0101001100101000111: color_data = Z;
		19'b0101001100101001000: color_data = Z;
		19'b0101001100101001001: color_data = Z;
		19'b0101001100101001010: color_data = Z;
		19'b0101001100101001011: color_data = Z;
		19'b0101001100101001100: color_data = Z;
		19'b0101001100101001101: color_data = Z;
		19'b0101001100101001110: color_data = Z;
		19'b0101001100101001111: color_data = Z;
		19'b0101001100101010000: color_data = Z;
		19'b0101001100101010001: color_data = Z;
		19'b0101001100101010010: color_data = Z;
		19'b0101001100101010011: color_data = Z;
		19'b0101001100101010100: color_data = Z;
		19'b0101001100101010101: color_data = Z;
		19'b0101001100101010110: color_data = Z;
		19'b0101001100101010111: color_data = Z;
		19'b0101001100101011000: color_data = Z;
		19'b0101001100101011001: color_data = Z;
		19'b0101001100101011010: color_data = Z;
		19'b0101001100101011011: color_data = Z;
		19'b0101001100101011100: color_data = Z;
		19'b0101001100101011101: color_data = Z;
		19'b0101001100101011110: color_data = Z;
		19'b0101001100101011111: color_data = Z;
		19'b0101001100101100000: color_data = Z;
		19'b0101001100101100001: color_data = Z;
		19'b0101001100101100010: color_data = Z;
		19'b0101001100101100011: color_data = Z;
		19'b0101001100101100100: color_data = Z;
		19'b0101001100101100101: color_data = Z;
		19'b0101001100101100110: color_data = Z;
		19'b0101001100101100111: color_data = Z;
		19'b0101001100101101000: color_data = Z;
		19'b0101001100101101001: color_data = Z;
		19'b0101001100101101010: color_data = Z;
		19'b0101001100101101011: color_data = Z;
		19'b0101001100101101100: color_data = Z;
		19'b0101001100101101101: color_data = Z;
		19'b0101001100101101110: color_data = Z;
		19'b0101001100101101111: color_data = Z;
		19'b0101001100101110000: color_data = Z;
		19'b0101001100101110001: color_data = Z;
		19'b0101001100101110010: color_data = Z;
		19'b0101001100101110011: color_data = Z;
		19'b0101001100101110100: color_data = Z;
		19'b0101001100101110101: color_data = Z;
		19'b0101001100101110110: color_data = Z;
		19'b0101001100101110111: color_data = Z;
		19'b0101001100101111000: color_data = Z;
		19'b0101001100101111001: color_data = Z;
		19'b0101001100101111010: color_data = Z;
		19'b0101001100101111011: color_data = Z;
		19'b0101001100101111100: color_data = Z;
		19'b0101001100101111101: color_data = Z;
		19'b0101001100101111110: color_data = Z;
		19'b0101001100101111111: color_data = Z;
		19'b0101001100110000000: color_data = Z;
		19'b0101001100111001111: color_data = Z;
		19'b0101001100111010000: color_data = Z;
		19'b0101001100111010001: color_data = Z;
		19'b0101001100111010010: color_data = Z;
		19'b0101001100111010011: color_data = Z;
		19'b0101001100111010100: color_data = Z;
		19'b0101001100111010110: color_data = Z;
		19'b0101001100111010111: color_data = Z;
		19'b0101001100111011000: color_data = Z;
		19'b0101001100111011001: color_data = Z;
		19'b0101001100111011010: color_data = Z;
		19'b0101001100111011011: color_data = Z;
		19'b0101001100111011100: color_data = Z;
		19'b0101001100111011101: color_data = Z;
		19'b0101001110100011110: color_data = Z;
		19'b0101001110100011111: color_data = Z;
		19'b0101001110100100000: color_data = Z;
		19'b0101001110100100001: color_data = Z;
		19'b0101001110100100010: color_data = Z;
		19'b0101001110100100011: color_data = Z;
		19'b0101001110100100100: color_data = Z;
		19'b0101001110100100101: color_data = Z;
		19'b0101001110100101010: color_data = Z;
		19'b0101001110100101011: color_data = Z;
		19'b0101001110100101100: color_data = Z;
		19'b0101001110100101101: color_data = Z;
		19'b0101001110100101110: color_data = Z;
		19'b0101001110100101111: color_data = Z;
		19'b0101001110100110000: color_data = Z;
		19'b0101001110100110001: color_data = Z;
		19'b0101001110100110010: color_data = Z;
		19'b0101001110100110011: color_data = Z;
		19'b0101001110100110100: color_data = Z;
		19'b0101001110100110101: color_data = Z;
		19'b0101001110100110110: color_data = Z;
		19'b0101001110100110111: color_data = Z;
		19'b0101001110100111000: color_data = Z;
		19'b0101001110100111001: color_data = Z;
		19'b0101001110100111010: color_data = Z;
		19'b0101001110100111011: color_data = Z;
		19'b0101001110100111100: color_data = Z;
		19'b0101001110100111101: color_data = Z;
		19'b0101001110100111110: color_data = Z;
		19'b0101001110100111111: color_data = Z;
		19'b0101001110101000000: color_data = Z;
		19'b0101001110101000001: color_data = Z;
		19'b0101001110101000010: color_data = Z;
		19'b0101001110101000011: color_data = Z;
		19'b0101001110101000100: color_data = Z;
		19'b0101001110101000101: color_data = Z;
		19'b0101001110101000110: color_data = Z;
		19'b0101001110101000111: color_data = Z;
		19'b0101001110101001000: color_data = Z;
		19'b0101001110101001001: color_data = Z;
		19'b0101001110101001010: color_data = Z;
		19'b0101001110101001011: color_data = Z;
		19'b0101001110101001100: color_data = Z;
		19'b0101001110101001101: color_data = Z;
		19'b0101001110101001110: color_data = Z;
		19'b0101001110101001111: color_data = Z;
		19'b0101001110101010000: color_data = Z;
		19'b0101001110101010001: color_data = Z;
		19'b0101001110101010010: color_data = Z;
		19'b0101001110101010011: color_data = Z;
		19'b0101001110101010100: color_data = Z;
		19'b0101001110101010101: color_data = Z;
		19'b0101001110101010110: color_data = Z;
		19'b0101001110101010111: color_data = Z;
		19'b0101001110101011000: color_data = Z;
		19'b0101001110101011001: color_data = Z;
		19'b0101001110101011010: color_data = Z;
		19'b0101001110101011011: color_data = Z;
		19'b0101001110101011100: color_data = Z;
		19'b0101001110101011101: color_data = Z;
		19'b0101001110101011110: color_data = Z;
		19'b0101001110101011111: color_data = Z;
		19'b0101001110101100000: color_data = Z;
		19'b0101001110101100001: color_data = Z;
		19'b0101001110101100010: color_data = Z;
		19'b0101001110101100011: color_data = Z;
		19'b0101001110101100100: color_data = Z;
		19'b0101001110101100101: color_data = Z;
		19'b0101001110101100110: color_data = Z;
		19'b0101001110101100111: color_data = Z;
		19'b0101001110101101000: color_data = Z;
		19'b0101001110101101001: color_data = Z;
		19'b0101001110101101010: color_data = Z;
		19'b0101001110101101011: color_data = Z;
		19'b0101001110101101100: color_data = Z;
		19'b0101001110101101101: color_data = Z;
		19'b0101001110101101110: color_data = Z;
		19'b0101001110101101111: color_data = Z;
		19'b0101001110101110000: color_data = Z;
		19'b0101001110101110001: color_data = Z;
		19'b0101001110101110010: color_data = Z;
		19'b0101001110101110011: color_data = Z;
		19'b0101001110101110100: color_data = Z;
		19'b0101001110101110101: color_data = Z;
		19'b0101001110101110110: color_data = Z;
		19'b0101001110101110111: color_data = Z;
		19'b0101001110101111000: color_data = Z;
		19'b0101001110101111001: color_data = Z;
		19'b0101001110101111010: color_data = Z;
		19'b0101001110101111011: color_data = Z;
		19'b0101001110101111100: color_data = Z;
		19'b0101001110101111101: color_data = Z;
		19'b0101001110101111110: color_data = Z;
		19'b0101001110101111111: color_data = Z;
		19'b0101001110110000000: color_data = Z;
		19'b0101001110111001111: color_data = Z;
		19'b0101001110111010000: color_data = Z;
		19'b0101001110111010001: color_data = Z;
		19'b0101001110111010010: color_data = Z;
		19'b0101001110111010011: color_data = Z;
		19'b0101001110111010100: color_data = Z;
		19'b0101001110111010110: color_data = Z;
		19'b0101001110111010111: color_data = Z;
		19'b0101001110111011000: color_data = Z;
		19'b0101001110111011001: color_data = Z;
		19'b0101001110111011010: color_data = Z;
		19'b0101001110111011011: color_data = Z;
		19'b0101001110111011100: color_data = Z;
		19'b0101001110111011101: color_data = Z;
		19'b0101001110111100001: color_data = Z;
		19'b0101010000100011110: color_data = Z;
		19'b0101010000100011111: color_data = Z;
		19'b0101010000100100000: color_data = Z;
		19'b0101010000100100001: color_data = Z;
		19'b0101010000100100010: color_data = Z;
		19'b0101010000100100011: color_data = Z;
		19'b0101010000100101010: color_data = Z;
		19'b0101010000100101011: color_data = Z;
		19'b0101010000100101100: color_data = Z;
		19'b0101010000100101101: color_data = Z;
		19'b0101010000100101110: color_data = Z;
		19'b0101010000100101111: color_data = Z;
		19'b0101010000100110000: color_data = Z;
		19'b0101010000100110001: color_data = Z;
		19'b0101010000100110010: color_data = Z;
		19'b0101010000100110011: color_data = Z;
		19'b0101010000100110100: color_data = Z;
		19'b0101010000100110101: color_data = Z;
		19'b0101010000100110110: color_data = Z;
		19'b0101010000100110111: color_data = Z;
		19'b0101010000100111000: color_data = Z;
		19'b0101010000100111001: color_data = Z;
		19'b0101010000100111010: color_data = Z;
		19'b0101010000100111011: color_data = Z;
		19'b0101010000100111100: color_data = Z;
		19'b0101010000100111101: color_data = Z;
		19'b0101010000100111110: color_data = Z;
		19'b0101010000100111111: color_data = Z;
		19'b0101010000101000000: color_data = Z;
		19'b0101010000101000001: color_data = Z;
		19'b0101010000101000010: color_data = Z;
		19'b0101010000101000011: color_data = Z;
		19'b0101010000101000100: color_data = Z;
		19'b0101010000101000101: color_data = Z;
		19'b0101010000101000110: color_data = Z;
		19'b0101010000101000111: color_data = Z;
		19'b0101010000101001000: color_data = Z;
		19'b0101010000101001001: color_data = Z;
		19'b0101010000101001010: color_data = Z;
		19'b0101010000101001011: color_data = Z;
		19'b0101010000101001100: color_data = Z;
		19'b0101010000101001101: color_data = Z;
		19'b0101010000101001110: color_data = Z;
		19'b0101010000101001111: color_data = Z;
		19'b0101010000101010000: color_data = Z;
		19'b0101010000101010001: color_data = Z;
		19'b0101010000101010010: color_data = Z;
		19'b0101010000101010011: color_data = Z;
		19'b0101010000101010100: color_data = Z;
		19'b0101010000101010101: color_data = Z;
		19'b0101010000101010110: color_data = Z;
		19'b0101010000101010111: color_data = Z;
		19'b0101010000101011000: color_data = Z;
		19'b0101010000101011001: color_data = Z;
		19'b0101010000101011010: color_data = Z;
		19'b0101010000101011011: color_data = Z;
		19'b0101010000101011100: color_data = Z;
		19'b0101010000101011101: color_data = Z;
		19'b0101010000101011110: color_data = Z;
		19'b0101010000101011111: color_data = Z;
		19'b0101010000101100000: color_data = Z;
		19'b0101010000101100001: color_data = Z;
		19'b0101010000101100010: color_data = Z;
		19'b0101010000101100011: color_data = Z;
		19'b0101010000101100100: color_data = Z;
		19'b0101010000101100101: color_data = Z;
		19'b0101010000101100110: color_data = Z;
		19'b0101010000101100111: color_data = Z;
		19'b0101010000101101000: color_data = Z;
		19'b0101010000101101001: color_data = Z;
		19'b0101010000101101010: color_data = Z;
		19'b0101010000101101011: color_data = Z;
		19'b0101010000101101100: color_data = Z;
		19'b0101010000101101101: color_data = Z;
		19'b0101010000101101110: color_data = Z;
		19'b0101010000101101111: color_data = Z;
		19'b0101010000101110000: color_data = Z;
		19'b0101010000101110001: color_data = Z;
		19'b0101010000101110010: color_data = Z;
		19'b0101010000101110011: color_data = Z;
		19'b0101010000101110100: color_data = Z;
		19'b0101010000101110101: color_data = Z;
		19'b0101010000101110110: color_data = Z;
		19'b0101010000101110111: color_data = Z;
		19'b0101010000101111000: color_data = Z;
		19'b0101010000101111001: color_data = Z;
		19'b0101010000101111010: color_data = Z;
		19'b0101010000101111011: color_data = Z;
		19'b0101010000101111100: color_data = Z;
		19'b0101010000101111101: color_data = Z;
		19'b0101010000101111110: color_data = Z;
		19'b0101010000101111111: color_data = Z;
		19'b0101010000110000000: color_data = Z;
		19'b0101010000110000001: color_data = Z;
		19'b0101010000111001111: color_data = Z;
		19'b0101010000111010000: color_data = Z;
		19'b0101010000111010001: color_data = Z;
		19'b0101010000111010010: color_data = Z;
		19'b0101010000111010011: color_data = Z;
		19'b0101010000111010100: color_data = Z;
		19'b0101010000111010110: color_data = Z;
		19'b0101010000111010111: color_data = Z;
		19'b0101010000111011000: color_data = Z;
		19'b0101010000111011001: color_data = Z;
		19'b0101010000111011010: color_data = Z;
		19'b0101010000111011011: color_data = Z;
		19'b0101010000111011100: color_data = Z;
		19'b0101010000111011101: color_data = Z;
		19'b0101010010100011110: color_data = Z;
		19'b0101010010100011111: color_data = Z;
		19'b0101010010100100000: color_data = Z;
		19'b0101010010100100001: color_data = Z;
		19'b0101010010100100010: color_data = Z;
		19'b0101010010100100011: color_data = Z;
		19'b0101010010100100101: color_data = Z;
		19'b0101010010100101001: color_data = Z;
		19'b0101010010100101010: color_data = Z;
		19'b0101010010100101011: color_data = Z;
		19'b0101010010100101100: color_data = Z;
		19'b0101010010100101101: color_data = Z;
		19'b0101010010100101110: color_data = Z;
		19'b0101010010100101111: color_data = Z;
		19'b0101010010100110000: color_data = Z;
		19'b0101010010100110001: color_data = Z;
		19'b0101010010100110010: color_data = Z;
		19'b0101010010100110011: color_data = Z;
		19'b0101010010100110100: color_data = Z;
		19'b0101010010100110101: color_data = Z;
		19'b0101010010100110110: color_data = Z;
		19'b0101010010100110111: color_data = Z;
		19'b0101010010100111000: color_data = Z;
		19'b0101010010100111001: color_data = Z;
		19'b0101010010100111010: color_data = Z;
		19'b0101010010100111011: color_data = Z;
		19'b0101010010100111100: color_data = Z;
		19'b0101010010100111101: color_data = Z;
		19'b0101010010100111110: color_data = Z;
		19'b0101010010100111111: color_data = Z;
		19'b0101010010101000000: color_data = Z;
		19'b0101010010101000001: color_data = Z;
		19'b0101010010101000010: color_data = Z;
		19'b0101010010101000011: color_data = Z;
		19'b0101010010101000100: color_data = Z;
		19'b0101010010101000101: color_data = Z;
		19'b0101010010101000110: color_data = Z;
		19'b0101010010101000111: color_data = Z;
		19'b0101010010101001000: color_data = Z;
		19'b0101010010101001001: color_data = Z;
		19'b0101010010101001010: color_data = Z;
		19'b0101010010101001011: color_data = Z;
		19'b0101010010101001100: color_data = Z;
		19'b0101010010101001101: color_data = Z;
		19'b0101010010101001110: color_data = Z;
		19'b0101010010101001111: color_data = Z;
		19'b0101010010101010000: color_data = Z;
		19'b0101010010101010001: color_data = Z;
		19'b0101010010101010010: color_data = Z;
		19'b0101010010101010011: color_data = Z;
		19'b0101010010101010100: color_data = Z;
		19'b0101010010101010101: color_data = Z;
		19'b0101010010101010110: color_data = Z;
		19'b0101010010101010111: color_data = Z;
		19'b0101010010101011000: color_data = Z;
		19'b0101010010101011001: color_data = Z;
		19'b0101010010101011010: color_data = Z;
		19'b0101010010101011011: color_data = Z;
		19'b0101010010101011100: color_data = Z;
		19'b0101010010101011101: color_data = Z;
		19'b0101010010101011110: color_data = Z;
		19'b0101010010101011111: color_data = Z;
		19'b0101010010101100000: color_data = Z;
		19'b0101010010101100001: color_data = Z;
		19'b0101010010101100010: color_data = Z;
		19'b0101010010101100011: color_data = Z;
		19'b0101010010101100100: color_data = Z;
		19'b0101010010101100101: color_data = Z;
		19'b0101010010101100110: color_data = Z;
		19'b0101010010101100111: color_data = Z;
		19'b0101010010101101000: color_data = Z;
		19'b0101010010101101001: color_data = Z;
		19'b0101010010101101010: color_data = Z;
		19'b0101010010101101011: color_data = Z;
		19'b0101010010101101100: color_data = Z;
		19'b0101010010101101101: color_data = Z;
		19'b0101010010101101110: color_data = Z;
		19'b0101010010101101111: color_data = Z;
		19'b0101010010101110000: color_data = Z;
		19'b0101010010101110001: color_data = Z;
		19'b0101010010101110010: color_data = Z;
		19'b0101010010101110011: color_data = Z;
		19'b0101010010101110100: color_data = Z;
		19'b0101010010101110101: color_data = Z;
		19'b0101010010101110110: color_data = Z;
		19'b0101010010101110111: color_data = Z;
		19'b0101010010101111000: color_data = Z;
		19'b0101010010101111001: color_data = Z;
		19'b0101010010101111010: color_data = Z;
		19'b0101010010101111011: color_data = Z;
		19'b0101010010101111100: color_data = Z;
		19'b0101010010101111101: color_data = Z;
		19'b0101010010101111110: color_data = Z;
		19'b0101010010101111111: color_data = Z;
		19'b0101010010110000000: color_data = Z;
		19'b0101010010110000001: color_data = Z;
		19'b0101010010111001111: color_data = Z;
		19'b0101010010111010000: color_data = Z;
		19'b0101010010111010001: color_data = Z;
		19'b0101010010111010010: color_data = Z;
		19'b0101010010111010011: color_data = Z;
		19'b0101010010111010100: color_data = Z;
		19'b0101010010111010110: color_data = Z;
		19'b0101010010111010111: color_data = Z;
		19'b0101010010111011000: color_data = Z;
		19'b0101010010111011001: color_data = Z;
		19'b0101010010111011010: color_data = Z;
		19'b0101010010111011011: color_data = Z;
		19'b0101010010111011100: color_data = Z;
		19'b0101010100100011110: color_data = Z;
		19'b0101010100100011111: color_data = Z;
		19'b0101010100100100000: color_data = Z;
		19'b0101010100100100001: color_data = Z;
		19'b0101010100100100010: color_data = Z;
		19'b0101010100100100011: color_data = Z;
		19'b0101010100100100100: color_data = Z;
		19'b0101010100100101000: color_data = Z;
		19'b0101010100100101001: color_data = Z;
		19'b0101010100100101010: color_data = Z;
		19'b0101010100100101011: color_data = Z;
		19'b0101010100100101100: color_data = Z;
		19'b0101010100100101101: color_data = Z;
		19'b0101010100100101110: color_data = Z;
		19'b0101010100100101111: color_data = Z;
		19'b0101010100100110000: color_data = Z;
		19'b0101010100100110001: color_data = Z;
		19'b0101010100100110010: color_data = Z;
		19'b0101010100100110011: color_data = Z;
		19'b0101010100100110100: color_data = Z;
		19'b0101010100100110101: color_data = Z;
		19'b0101010100100110110: color_data = Z;
		19'b0101010100100110111: color_data = Z;
		19'b0101010100100111000: color_data = Z;
		19'b0101010100100111001: color_data = Z;
		19'b0101010100100111010: color_data = Z;
		19'b0101010100100111011: color_data = Z;
		19'b0101010100100111100: color_data = Z;
		19'b0101010100100111101: color_data = Z;
		19'b0101010100100111110: color_data = Z;
		19'b0101010100100111111: color_data = Z;
		19'b0101010100101000000: color_data = Z;
		19'b0101010100101000001: color_data = Z;
		19'b0101010100101000010: color_data = Z;
		19'b0101010100101000011: color_data = Z;
		19'b0101010100101000100: color_data = Z;
		19'b0101010100101000101: color_data = Z;
		19'b0101010100101000110: color_data = Z;
		19'b0101010100101000111: color_data = Z;
		19'b0101010100101001000: color_data = Z;
		19'b0101010100101001001: color_data = Z;
		19'b0101010100101001010: color_data = Z;
		19'b0101010100101001011: color_data = Z;
		19'b0101010100101001100: color_data = Z;
		19'b0101010100101001101: color_data = Z;
		19'b0101010100101001110: color_data = Z;
		19'b0101010100101001111: color_data = Z;
		19'b0101010100101010000: color_data = Z;
		19'b0101010100101010001: color_data = Z;
		19'b0101010100101010010: color_data = Z;
		19'b0101010100101010011: color_data = Z;
		19'b0101010100101010100: color_data = Z;
		19'b0101010100101010101: color_data = Z;
		19'b0101010100101010110: color_data = Z;
		19'b0101010100101010111: color_data = Z;
		19'b0101010100101011000: color_data = Z;
		19'b0101010100101011001: color_data = Z;
		19'b0101010100101011010: color_data = Z;
		19'b0101010100101011011: color_data = Z;
		19'b0101010100101011100: color_data = Z;
		19'b0101010100101011101: color_data = Z;
		19'b0101010100101011110: color_data = Z;
		19'b0101010100101011111: color_data = Z;
		19'b0101010100101100000: color_data = Z;
		19'b0101010100101100001: color_data = Z;
		19'b0101010100101100010: color_data = Z;
		19'b0101010100101100011: color_data = Z;
		19'b0101010100101100100: color_data = Z;
		19'b0101010100101100101: color_data = Z;
		19'b0101010100101100110: color_data = Z;
		19'b0101010100101100111: color_data = Z;
		19'b0101010100101101000: color_data = Z;
		19'b0101010100101101001: color_data = Z;
		19'b0101010100101101010: color_data = Z;
		19'b0101010100101101011: color_data = Z;
		19'b0101010100101101100: color_data = Z;
		19'b0101010100101101101: color_data = Z;
		19'b0101010100101101110: color_data = Z;
		19'b0101010100101101111: color_data = Z;
		19'b0101010100101110000: color_data = Z;
		19'b0101010100101110001: color_data = Z;
		19'b0101010100101110010: color_data = Z;
		19'b0101010100101110011: color_data = Z;
		19'b0101010100101110100: color_data = Z;
		19'b0101010100101110101: color_data = Z;
		19'b0101010100101110110: color_data = Z;
		19'b0101010100101110111: color_data = Z;
		19'b0101010100101111000: color_data = Z;
		19'b0101010100101111001: color_data = Z;
		19'b0101010100101111010: color_data = Z;
		19'b0101010100101111011: color_data = Z;
		19'b0101010100101111100: color_data = Z;
		19'b0101010100101111101: color_data = Z;
		19'b0101010100101111110: color_data = Z;
		19'b0101010100101111111: color_data = Z;
		19'b0101010100110000000: color_data = Z;
		19'b0101010100110000001: color_data = Z;
		19'b0101010100111001111: color_data = Z;
		19'b0101010100111010000: color_data = Z;
		19'b0101010100111010001: color_data = Z;
		19'b0101010100111010010: color_data = Z;
		19'b0101010100111010011: color_data = Z;
		19'b0101010100111010100: color_data = Z;
		19'b0101010100111010110: color_data = Z;
		19'b0101010100111010111: color_data = Z;
		19'b0101010100111011000: color_data = Z;
		19'b0101010100111011001: color_data = Z;
		19'b0101010100111011010: color_data = Z;
		19'b0101010100111011011: color_data = Z;
		19'b0101010110100011110: color_data = Z;
		19'b0101010110100011111: color_data = Z;
		19'b0101010110100100000: color_data = Z;
		19'b0101010110100100001: color_data = Z;
		19'b0101010110100100010: color_data = Z;
		19'b0101010110100100011: color_data = Z;
		19'b0101010110100100100: color_data = Z;
		19'b0101010110100100111: color_data = Z;
		19'b0101010110100101000: color_data = Z;
		19'b0101010110100101001: color_data = Z;
		19'b0101010110100101010: color_data = Z;
		19'b0101010110100101011: color_data = Z;
		19'b0101010110100101100: color_data = Z;
		19'b0101010110100101101: color_data = Z;
		19'b0101010110100101110: color_data = Z;
		19'b0101010110100101111: color_data = Z;
		19'b0101010110100110000: color_data = Z;
		19'b0101010110100110001: color_data = Z;
		19'b0101010110100110010: color_data = Z;
		19'b0101010110100110011: color_data = Z;
		19'b0101010110100110100: color_data = Z;
		19'b0101010110100110101: color_data = Z;
		19'b0101010110100110110: color_data = Z;
		19'b0101010110100110111: color_data = Z;
		19'b0101010110100111000: color_data = Z;
		19'b0101010110100111001: color_data = Z;
		19'b0101010110100111010: color_data = Z;
		19'b0101010110100111011: color_data = Z;
		19'b0101010110100111100: color_data = Z;
		19'b0101010110100111101: color_data = Z;
		19'b0101010110100111110: color_data = Z;
		19'b0101010110100111111: color_data = Z;
		19'b0101010110101000000: color_data = Z;
		19'b0101010110101000001: color_data = Z;
		19'b0101010110101000010: color_data = Z;
		19'b0101010110101000011: color_data = Z;
		19'b0101010110101000100: color_data = Z;
		19'b0101010110101000101: color_data = Z;
		19'b0101010110101000110: color_data = Z;
		19'b0101010110101000111: color_data = Z;
		19'b0101010110101001000: color_data = Z;
		19'b0101010110101001001: color_data = Z;
		19'b0101010110101001010: color_data = Z;
		19'b0101010110101001011: color_data = Z;
		19'b0101010110101001100: color_data = Z;
		19'b0101010110101001101: color_data = Z;
		19'b0101010110101001110: color_data = Z;
		19'b0101010110101001111: color_data = Z;
		19'b0101010110101010000: color_data = Z;
		19'b0101010110101010001: color_data = Z;
		19'b0101010110101010010: color_data = Z;
		19'b0101010110101010011: color_data = Z;
		19'b0101010110101010100: color_data = Z;
		19'b0101010110101010101: color_data = Z;
		19'b0101010110101010110: color_data = Z;
		19'b0101010110101010111: color_data = Z;
		19'b0101010110101011000: color_data = Z;
		19'b0101010110101011001: color_data = Z;
		19'b0101010110101011010: color_data = Z;
		19'b0101010110101011011: color_data = Z;
		19'b0101010110101011100: color_data = Z;
		19'b0101010110101011101: color_data = Z;
		19'b0101010110101011110: color_data = Z;
		19'b0101010110101011111: color_data = Z;
		19'b0101010110101100000: color_data = Z;
		19'b0101010110101100001: color_data = Z;
		19'b0101010110101100010: color_data = Z;
		19'b0101010110101100011: color_data = Z;
		19'b0101010110101100100: color_data = Z;
		19'b0101010110101100101: color_data = Z;
		19'b0101010110101100110: color_data = Z;
		19'b0101010110101100111: color_data = Z;
		19'b0101010110101101000: color_data = Z;
		19'b0101010110101101001: color_data = Z;
		19'b0101010110101101010: color_data = Z;
		19'b0101010110101101011: color_data = Z;
		19'b0101010110101101100: color_data = Z;
		19'b0101010110101101101: color_data = Z;
		19'b0101010110101101110: color_data = Z;
		19'b0101010110101101111: color_data = Z;
		19'b0101010110101110000: color_data = Z;
		19'b0101010110101110001: color_data = Z;
		19'b0101010110101110010: color_data = Z;
		19'b0101010110101110011: color_data = Z;
		19'b0101010110101110100: color_data = Z;
		19'b0101010110101110101: color_data = Z;
		19'b0101010110101110110: color_data = Z;
		19'b0101010110101110111: color_data = Z;
		19'b0101010110101111000: color_data = Z;
		19'b0101010110101111001: color_data = Z;
		19'b0101010110101111010: color_data = Z;
		19'b0101010110101111011: color_data = Z;
		19'b0101010110101111100: color_data = Z;
		19'b0101010110101111101: color_data = Z;
		19'b0101010110101111110: color_data = Z;
		19'b0101010110101111111: color_data = Z;
		19'b0101010110110000000: color_data = Z;
		19'b0101010110110000001: color_data = Z;
		19'b0101010110111001111: color_data = Z;
		19'b0101010110111010000: color_data = Z;
		19'b0101010110111010001: color_data = Z;
		19'b0101010110111010010: color_data = Z;
		19'b0101010110111010011: color_data = Z;
		19'b0101010110111010100: color_data = Z;
		19'b0101010110111010110: color_data = Z;
		19'b0101010110111010111: color_data = Z;
		19'b0101010110111011000: color_data = Z;
		19'b0101010110111011001: color_data = Z;
		19'b0101010110111011010: color_data = Z;
		19'b0101010110111011011: color_data = Z;
		19'b0101011000100011111: color_data = Z;
		19'b0101011000100100000: color_data = Z;
		19'b0101011000100100001: color_data = Z;
		19'b0101011000100100010: color_data = Z;
		19'b0101011000100100011: color_data = Z;
		19'b0101011000100100100: color_data = Z;
		19'b0101011000100100101: color_data = Z;
		19'b0101011000100100110: color_data = Z;
		19'b0101011000100100111: color_data = Z;
		19'b0101011000100101000: color_data = Z;
		19'b0101011000100101001: color_data = Z;
		19'b0101011000100101010: color_data = Z;
		19'b0101011000100101011: color_data = Z;
		19'b0101011000100101100: color_data = Z;
		19'b0101011000100101101: color_data = Z;
		19'b0101011000100101110: color_data = Z;
		19'b0101011000100101111: color_data = Z;
		19'b0101011000100110000: color_data = Z;
		19'b0101011000100110001: color_data = Z;
		19'b0101011000100110010: color_data = Z;
		19'b0101011000100110011: color_data = Z;
		19'b0101011000100110100: color_data = Z;
		19'b0101011000100110101: color_data = Z;
		19'b0101011000100110110: color_data = Z;
		19'b0101011000100110111: color_data = Z;
		19'b0101011000100111000: color_data = Z;
		19'b0101011000100111001: color_data = Z;
		19'b0101011000100111010: color_data = Z;
		19'b0101011000100111011: color_data = Z;
		19'b0101011000100111100: color_data = Z;
		19'b0101011000100111101: color_data = Z;
		19'b0101011000100111110: color_data = Z;
		19'b0101011000100111111: color_data = Z;
		19'b0101011000101000000: color_data = Z;
		19'b0101011000101000001: color_data = Z;
		19'b0101011000101000010: color_data = Z;
		19'b0101011000101000011: color_data = Z;
		19'b0101011000101000100: color_data = Z;
		19'b0101011000101000101: color_data = Z;
		19'b0101011000101000110: color_data = Z;
		19'b0101011000101000111: color_data = Z;
		19'b0101011000101001000: color_data = Z;
		19'b0101011000101001001: color_data = Z;
		19'b0101011000101001010: color_data = Z;
		19'b0101011000101001011: color_data = Z;
		19'b0101011000101001100: color_data = Z;
		19'b0101011000101001101: color_data = Z;
		19'b0101011000101001110: color_data = Z;
		19'b0101011000101001111: color_data = Z;
		19'b0101011000101010000: color_data = Z;
		19'b0101011000101010001: color_data = Z;
		19'b0101011000101010010: color_data = Z;
		19'b0101011000101010011: color_data = Z;
		19'b0101011000101010100: color_data = Z;
		19'b0101011000101010101: color_data = Z;
		19'b0101011000101010110: color_data = Z;
		19'b0101011000101010111: color_data = Z;
		19'b0101011000101011000: color_data = Z;
		19'b0101011000101011001: color_data = Z;
		19'b0101011000101011010: color_data = Z;
		19'b0101011000101011011: color_data = Z;
		19'b0101011000101011100: color_data = Z;
		19'b0101011000101011101: color_data = Z;
		19'b0101011000101011110: color_data = Z;
		19'b0101011000101011111: color_data = Z;
		19'b0101011000101100000: color_data = Z;
		19'b0101011000101100001: color_data = Z;
		19'b0101011000101100010: color_data = Z;
		19'b0101011000101100011: color_data = Z;
		19'b0101011000101100100: color_data = Z;
		19'b0101011000101100101: color_data = Z;
		19'b0101011000101100110: color_data = Z;
		19'b0101011000101100111: color_data = Z;
		19'b0101011000101101000: color_data = Z;
		19'b0101011000101101001: color_data = Z;
		19'b0101011000101101010: color_data = Z;
		19'b0101011000101101011: color_data = Z;
		19'b0101011000101101100: color_data = Z;
		19'b0101011000101101101: color_data = Z;
		19'b0101011000101101110: color_data = Z;
		19'b0101011000101101111: color_data = Z;
		19'b0101011000101110000: color_data = Z;
		19'b0101011000101110001: color_data = Z;
		19'b0101011000101110010: color_data = Z;
		19'b0101011000101110011: color_data = Z;
		19'b0101011000101110100: color_data = Z;
		19'b0101011000101110101: color_data = Z;
		19'b0101011000101110110: color_data = Z;
		19'b0101011000101110111: color_data = Z;
		19'b0101011000101111000: color_data = Z;
		19'b0101011000101111001: color_data = Z;
		19'b0101011000101111010: color_data = Z;
		19'b0101011000101111011: color_data = Z;
		19'b0101011000101111100: color_data = Z;
		19'b0101011000101111101: color_data = Z;
		19'b0101011000101111110: color_data = Z;
		19'b0101011000101111111: color_data = Z;
		19'b0101011000110000000: color_data = Z;
		19'b0101011000110000001: color_data = Z;
		19'b0101011000110000010: color_data = Z;
		19'b0101011000111001111: color_data = Z;
		19'b0101011000111010000: color_data = Z;
		19'b0101011000111010001: color_data = Z;
		19'b0101011000111010010: color_data = Z;
		19'b0101011000111010011: color_data = Z;
		19'b0101011000111010100: color_data = Z;
		19'b0101011000111010101: color_data = Z;
		19'b0101011000111010110: color_data = Z;
		19'b0101011000111010111: color_data = Z;
		19'b0101011000111011000: color_data = Z;
		19'b0101011000111011001: color_data = Z;
		19'b0101011000111011010: color_data = Z;
		19'b0101011000111011011: color_data = Z;
		19'b0101011010100011111: color_data = Z;
		19'b0101011010100100000: color_data = Z;
		19'b0101011010100100001: color_data = Z;
		19'b0101011010100100010: color_data = Z;
		19'b0101011010100100011: color_data = Z;
		19'b0101011010100100100: color_data = Z;
		19'b0101011010100100101: color_data = Z;
		19'b0101011010100100110: color_data = Z;
		19'b0101011010100100111: color_data = Z;
		19'b0101011010100101000: color_data = Z;
		19'b0101011010100101001: color_data = Z;
		19'b0101011010100101010: color_data = Z;
		19'b0101011010100101011: color_data = Z;
		19'b0101011010100101100: color_data = Z;
		19'b0101011010100101101: color_data = Z;
		19'b0101011010100101110: color_data = Z;
		19'b0101011010100101111: color_data = Z;
		19'b0101011010100110000: color_data = Z;
		19'b0101011010100110001: color_data = Z;
		19'b0101011010100110010: color_data = Z;
		19'b0101011010100110011: color_data = Z;
		19'b0101011010100110100: color_data = Z;
		19'b0101011010100110101: color_data = Z;
		19'b0101011010100110110: color_data = Z;
		19'b0101011010100110111: color_data = Z;
		19'b0101011010100111000: color_data = Z;
		19'b0101011010100111001: color_data = Z;
		19'b0101011010100111010: color_data = Z;
		19'b0101011010100111011: color_data = Z;
		19'b0101011010100111100: color_data = Z;
		19'b0101011010100111101: color_data = Z;
		19'b0101011010100111110: color_data = Z;
		19'b0101011010100111111: color_data = Z;
		19'b0101011010101000000: color_data = Z;
		19'b0101011010101000001: color_data = Z;
		19'b0101011010101000010: color_data = Z;
		19'b0101011010101000011: color_data = Z;
		19'b0101011010101000100: color_data = Z;
		19'b0101011010101000101: color_data = Z;
		19'b0101011010101000110: color_data = Z;
		19'b0101011010101000111: color_data = Z;
		19'b0101011010101001000: color_data = Z;
		19'b0101011010101001001: color_data = Z;
		19'b0101011010101001010: color_data = Z;
		19'b0101011010101001011: color_data = Z;
		19'b0101011010101001100: color_data = Z;
		19'b0101011010101001101: color_data = Z;
		19'b0101011010101001110: color_data = Z;
		19'b0101011010101001111: color_data = Z;
		19'b0101011010101010000: color_data = Z;
		19'b0101011010101010001: color_data = Z;
		19'b0101011010101010010: color_data = Z;
		19'b0101011010101010011: color_data = Z;
		19'b0101011010101010100: color_data = Z;
		19'b0101011010101010101: color_data = Z;
		19'b0101011010101010110: color_data = Z;
		19'b0101011010101010111: color_data = Z;
		19'b0101011010101011000: color_data = Z;
		19'b0101011010101011001: color_data = Z;
		19'b0101011010101011010: color_data = Z;
		19'b0101011010101011011: color_data = Z;
		19'b0101011010101011100: color_data = Z;
		19'b0101011010101011101: color_data = Z;
		19'b0101011010101011110: color_data = Z;
		19'b0101011010101011111: color_data = Z;
		19'b0101011010101100000: color_data = Z;
		19'b0101011010101100001: color_data = Z;
		19'b0101011010101100010: color_data = Z;
		19'b0101011010101100011: color_data = Z;
		19'b0101011010101100100: color_data = Z;
		19'b0101011010101100101: color_data = Z;
		19'b0101011010101100110: color_data = Z;
		19'b0101011010101100111: color_data = Z;
		19'b0101011010101101000: color_data = Z;
		19'b0101011010101101001: color_data = Z;
		19'b0101011010101101010: color_data = Z;
		19'b0101011010101101011: color_data = Z;
		19'b0101011010101101100: color_data = Z;
		19'b0101011010101101101: color_data = Z;
		19'b0101011010101101110: color_data = Z;
		19'b0101011010101101111: color_data = Z;
		19'b0101011010101110000: color_data = Z;
		19'b0101011010101110001: color_data = Z;
		19'b0101011010101110010: color_data = Z;
		19'b0101011010101110011: color_data = Z;
		19'b0101011010101110100: color_data = Z;
		19'b0101011010101110101: color_data = Z;
		19'b0101011010101110110: color_data = Z;
		19'b0101011010101110111: color_data = Z;
		19'b0101011010101111000: color_data = Z;
		19'b0101011010101111001: color_data = Z;
		19'b0101011010101111010: color_data = Z;
		19'b0101011010101111011: color_data = Z;
		19'b0101011010101111100: color_data = Z;
		19'b0101011010101111101: color_data = Z;
		19'b0101011010101111110: color_data = Z;
		19'b0101011010101111111: color_data = Z;
		19'b0101011010110000000: color_data = Z;
		19'b0101011010110000001: color_data = Z;
		19'b0101011010110000010: color_data = Z;
		19'b0101011010111001111: color_data = Z;
		19'b0101011010111010000: color_data = Z;
		19'b0101011010111010001: color_data = Z;
		19'b0101011010111010010: color_data = Z;
		19'b0101011010111010011: color_data = Z;
		19'b0101011010111010100: color_data = Z;
		19'b0101011010111010101: color_data = Z;
		19'b0101011010111010110: color_data = Z;
		19'b0101011010111010111: color_data = Z;
		19'b0101011010111011000: color_data = Z;
		19'b0101011010111011001: color_data = Z;
		19'b0101011010111011010: color_data = Z;
		19'b0101011010111011011: color_data = Z;
		19'b0101011100100011111: color_data = Z;
		19'b0101011100100100000: color_data = Z;
		19'b0101011100100100001: color_data = Z;
		19'b0101011100100100010: color_data = Z;
		19'b0101011100100100011: color_data = Z;
		19'b0101011100100100100: color_data = Z;
		19'b0101011100100100101: color_data = Z;
		19'b0101011100100100110: color_data = Z;
		19'b0101011100100100111: color_data = Z;
		19'b0101011100100101000: color_data = Z;
		19'b0101011100100101001: color_data = Z;
		19'b0101011100100101010: color_data = Z;
		19'b0101011100100101011: color_data = Z;
		19'b0101011100100101100: color_data = Z;
		19'b0101011100100101101: color_data = Z;
		19'b0101011100100101110: color_data = Z;
		19'b0101011100100101111: color_data = Z;
		19'b0101011100100110000: color_data = Z;
		19'b0101011100100110001: color_data = Z;
		19'b0101011100100110010: color_data = Z;
		19'b0101011100100110011: color_data = Z;
		19'b0101011100100110100: color_data = Z;
		19'b0101011100100110101: color_data = Z;
		19'b0101011100100110110: color_data = Z;
		19'b0101011100100110111: color_data = Z;
		19'b0101011100100111000: color_data = Z;
		19'b0101011100100111001: color_data = Z;
		19'b0101011100100111010: color_data = Z;
		19'b0101011100100111011: color_data = Z;
		19'b0101011100100111100: color_data = Z;
		19'b0101011100100111101: color_data = Z;
		19'b0101011100100111110: color_data = Z;
		19'b0101011100100111111: color_data = Z;
		19'b0101011100101000000: color_data = Z;
		19'b0101011100101000001: color_data = Z;
		19'b0101011100101000010: color_data = Z;
		19'b0101011100101000011: color_data = Z;
		19'b0101011100101000100: color_data = Z;
		19'b0101011100101000101: color_data = Z;
		19'b0101011100101000110: color_data = Z;
		19'b0101011100101000111: color_data = Z;
		19'b0101011100101001000: color_data = Z;
		19'b0101011100101001001: color_data = Z;
		19'b0101011100101001010: color_data = Z;
		19'b0101011100101001011: color_data = Z;
		19'b0101011100101001100: color_data = Z;
		19'b0101011100101001101: color_data = Z;
		19'b0101011100101001110: color_data = Z;
		19'b0101011100101001111: color_data = Z;
		19'b0101011100101010000: color_data = Z;
		19'b0101011100101010001: color_data = Z;
		19'b0101011100101010010: color_data = Z;
		19'b0101011100101010011: color_data = Z;
		19'b0101011100101010100: color_data = Z;
		19'b0101011100101010101: color_data = Z;
		19'b0101011100101010110: color_data = Z;
		19'b0101011100101010111: color_data = Z;
		19'b0101011100101011000: color_data = Z;
		19'b0101011100101011001: color_data = Z;
		19'b0101011100101011010: color_data = Z;
		19'b0101011100101011011: color_data = Z;
		19'b0101011100101011100: color_data = Z;
		19'b0101011100101011101: color_data = Z;
		19'b0101011100101011110: color_data = Z;
		19'b0101011100101011111: color_data = Z;
		19'b0101011100101100000: color_data = Z;
		19'b0101011100101100001: color_data = Z;
		19'b0101011100101100010: color_data = Z;
		19'b0101011100101100011: color_data = Z;
		19'b0101011100101100100: color_data = Z;
		19'b0101011100101100101: color_data = Z;
		19'b0101011100101100110: color_data = Z;
		19'b0101011100101100111: color_data = Z;
		19'b0101011100101101000: color_data = Z;
		19'b0101011100101101001: color_data = Z;
		19'b0101011100101101010: color_data = Z;
		19'b0101011100101101011: color_data = Z;
		19'b0101011100101101100: color_data = Z;
		19'b0101011100101101101: color_data = Z;
		19'b0101011100101101110: color_data = Z;
		19'b0101011100101101111: color_data = Z;
		19'b0101011100101110000: color_data = Z;
		19'b0101011100101110001: color_data = Z;
		19'b0101011100101110010: color_data = Z;
		19'b0101011100101110011: color_data = Z;
		19'b0101011100101110100: color_data = Z;
		19'b0101011100101110101: color_data = Z;
		19'b0101011100101110110: color_data = Z;
		19'b0101011100101110111: color_data = Z;
		19'b0101011100101111000: color_data = Z;
		19'b0101011100101111001: color_data = Z;
		19'b0101011100101111010: color_data = Z;
		19'b0101011100101111011: color_data = Z;
		19'b0101011100101111100: color_data = Z;
		19'b0101011100101111101: color_data = Z;
		19'b0101011100101111110: color_data = Z;
		19'b0101011100101111111: color_data = Z;
		19'b0101011100110000000: color_data = Z;
		19'b0101011100110000001: color_data = Z;
		19'b0101011100110000010: color_data = Z;
		19'b0101011100111001111: color_data = Z;
		19'b0101011100111010000: color_data = Z;
		19'b0101011100111010001: color_data = Z;
		19'b0101011100111010010: color_data = Z;
		19'b0101011100111010011: color_data = Z;
		19'b0101011100111010100: color_data = Z;
		19'b0101011100111010101: color_data = Z;
		19'b0101011100111010110: color_data = Z;
		19'b0101011100111010111: color_data = Z;
		19'b0101011100111011000: color_data = Z;
		19'b0101011100111011001: color_data = Z;
		19'b0101011100111011010: color_data = Z;
		19'b0101011100111011011: color_data = Z;
		19'b0101011110100011111: color_data = Z;
		19'b0101011110100100000: color_data = Z;
		19'b0101011110100100001: color_data = Z;
		19'b0101011110100100010: color_data = Z;
		19'b0101011110100100011: color_data = Z;
		19'b0101011110100100100: color_data = Z;
		19'b0101011110100100101: color_data = Z;
		19'b0101011110100100110: color_data = Z;
		19'b0101011110100100111: color_data = Z;
		19'b0101011110100101000: color_data = Z;
		19'b0101011110100101001: color_data = Z;
		19'b0101011110100101010: color_data = Z;
		19'b0101011110100101011: color_data = Z;
		19'b0101011110100101100: color_data = Z;
		19'b0101011110100101101: color_data = Z;
		19'b0101011110100101110: color_data = Z;
		19'b0101011110100101111: color_data = Z;
		19'b0101011110100110000: color_data = Z;
		19'b0101011110100110001: color_data = Z;
		19'b0101011110100110010: color_data = Z;
		19'b0101011110100110011: color_data = Z;
		19'b0101011110100110100: color_data = Z;
		19'b0101011110100110101: color_data = Z;
		19'b0101011110100110110: color_data = Z;
		19'b0101011110100110111: color_data = Z;
		19'b0101011110100111000: color_data = Z;
		19'b0101011110100111001: color_data = Z;
		19'b0101011110100111010: color_data = Z;
		19'b0101011110100111011: color_data = Z;
		19'b0101011110100111100: color_data = Z;
		19'b0101011110100111101: color_data = Z;
		19'b0101011110100111110: color_data = Z;
		19'b0101011110100111111: color_data = Z;
		19'b0101011110101000000: color_data = Z;
		19'b0101011110101000001: color_data = Z;
		19'b0101011110101000010: color_data = Z;
		19'b0101011110101000011: color_data = Z;
		19'b0101011110101000100: color_data = Z;
		19'b0101011110101000101: color_data = Z;
		19'b0101011110101000110: color_data = Z;
		19'b0101011110101000111: color_data = Z;
		19'b0101011110101001000: color_data = Z;
		19'b0101011110101001001: color_data = Z;
		19'b0101011110101001010: color_data = Z;
		19'b0101011110101001011: color_data = Z;
		19'b0101011110101001100: color_data = Z;
		19'b0101011110101001101: color_data = Z;
		19'b0101011110101001110: color_data = Z;
		19'b0101011110101001111: color_data = Z;
		19'b0101011110101010000: color_data = Z;
		19'b0101011110101010001: color_data = Z;
		19'b0101011110101010010: color_data = Z;
		19'b0101011110101010011: color_data = Z;
		19'b0101011110101010100: color_data = Z;
		19'b0101011110101010101: color_data = Z;
		19'b0101011110101010110: color_data = Z;
		19'b0101011110101010111: color_data = Z;
		19'b0101011110101011000: color_data = Z;
		19'b0101011110101011001: color_data = Z;
		19'b0101011110101011010: color_data = Z;
		19'b0101011110101011011: color_data = Z;
		19'b0101011110101011100: color_data = Z;
		19'b0101011110101011101: color_data = Z;
		19'b0101011110101011110: color_data = Z;
		19'b0101011110101011111: color_data = Z;
		19'b0101011110101100000: color_data = Z;
		19'b0101011110101100001: color_data = Z;
		19'b0101011110101100010: color_data = Z;
		19'b0101011110101100011: color_data = Z;
		19'b0101011110101100100: color_data = Z;
		19'b0101011110101100101: color_data = Z;
		19'b0101011110101100110: color_data = Z;
		19'b0101011110101100111: color_data = Z;
		19'b0101011110101101000: color_data = Z;
		19'b0101011110101101001: color_data = Z;
		19'b0101011110101101010: color_data = Z;
		19'b0101011110101101011: color_data = Z;
		19'b0101011110101101100: color_data = Z;
		19'b0101011110101101101: color_data = Z;
		19'b0101011110101101110: color_data = Z;
		19'b0101011110101101111: color_data = Z;
		19'b0101011110101110000: color_data = Z;
		19'b0101011110101110001: color_data = Z;
		19'b0101011110101110010: color_data = Z;
		19'b0101011110101110011: color_data = Z;
		19'b0101011110101110100: color_data = Z;
		19'b0101011110101110101: color_data = Z;
		19'b0101011110101110110: color_data = Z;
		19'b0101011110101110111: color_data = Z;
		19'b0101011110101111000: color_data = Z;
		19'b0101011110101111001: color_data = Z;
		19'b0101011110101111010: color_data = Z;
		19'b0101011110101111011: color_data = Z;
		19'b0101011110101111100: color_data = Z;
		19'b0101011110101111101: color_data = Z;
		19'b0101011110101111110: color_data = Z;
		19'b0101011110101111111: color_data = Z;
		19'b0101011110110000000: color_data = Z;
		19'b0101011110110000001: color_data = Z;
		19'b0101011110110000010: color_data = Z;
		19'b0101011110111001111: color_data = Z;
		19'b0101011110111010000: color_data = Z;
		19'b0101011110111010001: color_data = Z;
		19'b0101011110111010010: color_data = Z;
		19'b0101011110111010011: color_data = Z;
		19'b0101011110111010100: color_data = Z;
		19'b0101011110111010101: color_data = Z;
		19'b0101011110111010110: color_data = Z;
		19'b0101011110111010111: color_data = Z;
		19'b0101011110111011000: color_data = Z;
		19'b0101011110111011001: color_data = Z;
		19'b0101011110111011010: color_data = Z;
		19'b0101011110111011011: color_data = Z;
		19'b0101100000100011111: color_data = Z;
		19'b0101100000100100000: color_data = Z;
		19'b0101100000100100001: color_data = Z;
		19'b0101100000100100010: color_data = Z;
		19'b0101100000100100011: color_data = Z;
		19'b0101100000100100100: color_data = Z;
		19'b0101100000100100110: color_data = Z;
		19'b0101100000100100111: color_data = Z;
		19'b0101100000100101000: color_data = Z;
		19'b0101100000100101001: color_data = Z;
		19'b0101100000100101010: color_data = Z;
		19'b0101100000100101011: color_data = Z;
		19'b0101100000100101100: color_data = Z;
		19'b0101100000100101101: color_data = Z;
		19'b0101100000100101110: color_data = Z;
		19'b0101100000100101111: color_data = Z;
		19'b0101100000100110000: color_data = Z;
		19'b0101100000100110001: color_data = Z;
		19'b0101100000100110010: color_data = Z;
		19'b0101100000100110011: color_data = Z;
		19'b0101100000100110100: color_data = Z;
		19'b0101100000100110101: color_data = Z;
		19'b0101100000100110110: color_data = Z;
		19'b0101100000100110111: color_data = Z;
		19'b0101100000100111000: color_data = Z;
		19'b0101100000100111001: color_data = Z;
		19'b0101100000100111010: color_data = Z;
		19'b0101100000100111011: color_data = Z;
		19'b0101100000100111100: color_data = Z;
		19'b0101100000100111101: color_data = Z;
		19'b0101100000100111110: color_data = Z;
		19'b0101100000100111111: color_data = Z;
		19'b0101100000101000000: color_data = Z;
		19'b0101100000101000001: color_data = Z;
		19'b0101100000101000010: color_data = Z;
		19'b0101100000101000011: color_data = Z;
		19'b0101100000101000100: color_data = Z;
		19'b0101100000101000101: color_data = Z;
		19'b0101100000101000110: color_data = Z;
		19'b0101100000101000111: color_data = Z;
		19'b0101100000101001000: color_data = Z;
		19'b0101100000101001001: color_data = Z;
		19'b0101100000101001010: color_data = Z;
		19'b0101100000101001011: color_data = Z;
		19'b0101100000101001100: color_data = Z;
		19'b0101100000101001101: color_data = Z;
		19'b0101100000101001110: color_data = Z;
		19'b0101100000101001111: color_data = Z;
		19'b0101100000101010000: color_data = Z;
		19'b0101100000101010001: color_data = Z;
		19'b0101100000101010010: color_data = Z;
		19'b0101100000101010011: color_data = Z;
		19'b0101100000101010100: color_data = Z;
		19'b0101100000101010101: color_data = Z;
		19'b0101100000101010110: color_data = Z;
		19'b0101100000101010111: color_data = Z;
		19'b0101100000101011000: color_data = Z;
		19'b0101100000101011001: color_data = Z;
		19'b0101100000101011010: color_data = Z;
		19'b0101100000101011011: color_data = Z;
		19'b0101100000101011100: color_data = Z;
		19'b0101100000101011101: color_data = Z;
		19'b0101100000101011110: color_data = Z;
		19'b0101100000101011111: color_data = Z;
		19'b0101100000101100000: color_data = Z;
		19'b0101100000101100001: color_data = Z;
		19'b0101100000101100010: color_data = Z;
		19'b0101100000101100011: color_data = Z;
		19'b0101100000101100100: color_data = Z;
		19'b0101100000101100101: color_data = Z;
		19'b0101100000101100110: color_data = Z;
		19'b0101100000101100111: color_data = Z;
		19'b0101100000101101000: color_data = Z;
		19'b0101100000101101001: color_data = Z;
		19'b0101100000101101010: color_data = Z;
		19'b0101100000101101011: color_data = Z;
		19'b0101100000101101100: color_data = Z;
		19'b0101100000101101101: color_data = Z;
		19'b0101100000101101110: color_data = Z;
		19'b0101100000101101111: color_data = Z;
		19'b0101100000101110000: color_data = Z;
		19'b0101100000101110001: color_data = Z;
		19'b0101100000101110010: color_data = Z;
		19'b0101100000101110011: color_data = Z;
		19'b0101100000101110100: color_data = Z;
		19'b0101100000101110101: color_data = Z;
		19'b0101100000101110110: color_data = Z;
		19'b0101100000101110111: color_data = Z;
		19'b0101100000101111000: color_data = Z;
		19'b0101100000101111001: color_data = Z;
		19'b0101100000101111010: color_data = Z;
		19'b0101100000101111011: color_data = Z;
		19'b0101100000101111100: color_data = Z;
		19'b0101100000101111101: color_data = Z;
		19'b0101100000101111110: color_data = Z;
		19'b0101100000101111111: color_data = Z;
		19'b0101100000110000000: color_data = Z;
		19'b0101100000110000001: color_data = Z;
		19'b0101100000110000010: color_data = Z;
		19'b0101100000111001111: color_data = Z;
		19'b0101100000111010000: color_data = Z;
		19'b0101100000111010001: color_data = Z;
		19'b0101100000111010010: color_data = Z;
		19'b0101100000111010011: color_data = Z;
		19'b0101100000111010100: color_data = Z;
		19'b0101100000111010101: color_data = Z;
		19'b0101100000111010110: color_data = Z;
		19'b0101100000111010111: color_data = Z;
		19'b0101100000111011000: color_data = Z;
		19'b0101100000111011001: color_data = Z;
		19'b0101100000111011010: color_data = Z;
		19'b0101100000111011011: color_data = Z;
		19'b0101100010100011111: color_data = Z;
		19'b0101100010100100000: color_data = Z;
		19'b0101100010100100001: color_data = Z;
		19'b0101100010100100010: color_data = Z;
		19'b0101100010100100011: color_data = Z;
		19'b0101100010100100100: color_data = Z;
		19'b0101100010100100110: color_data = Z;
		19'b0101100010100100111: color_data = Z;
		19'b0101100010100101000: color_data = Z;
		19'b0101100010100101001: color_data = Z;
		19'b0101100010100101010: color_data = Z;
		19'b0101100010100101011: color_data = Z;
		19'b0101100010100101100: color_data = Z;
		19'b0101100010100101101: color_data = Z;
		19'b0101100010100101110: color_data = Z;
		19'b0101100010100101111: color_data = Z;
		19'b0101100010100110000: color_data = Z;
		19'b0101100010100110001: color_data = Z;
		19'b0101100010100110010: color_data = Z;
		19'b0101100010100110011: color_data = Z;
		19'b0101100010100110100: color_data = Z;
		19'b0101100010100110101: color_data = Z;
		19'b0101100010100110110: color_data = Z;
		19'b0101100010100110111: color_data = Z;
		19'b0101100010100111000: color_data = Z;
		19'b0101100010100111001: color_data = Z;
		19'b0101100010100111010: color_data = Z;
		19'b0101100010100111011: color_data = Z;
		19'b0101100010100111100: color_data = Z;
		19'b0101100010100111101: color_data = Z;
		19'b0101100010100111110: color_data = Z;
		19'b0101100010100111111: color_data = Z;
		19'b0101100010101000000: color_data = Z;
		19'b0101100010101000001: color_data = Z;
		19'b0101100010101000010: color_data = Z;
		19'b0101100010101000011: color_data = Z;
		19'b0101100010101000100: color_data = Z;
		19'b0101100010101000101: color_data = Z;
		19'b0101100010101000110: color_data = Z;
		19'b0101100010101000111: color_data = Z;
		19'b0101100010101001000: color_data = Z;
		19'b0101100010101001001: color_data = Z;
		19'b0101100010101001010: color_data = Z;
		19'b0101100010101001011: color_data = Z;
		19'b0101100010101001100: color_data = Z;
		19'b0101100010101001101: color_data = Z;
		19'b0101100010101001110: color_data = Z;
		19'b0101100010101001111: color_data = Z;
		19'b0101100010101010000: color_data = Z;
		19'b0101100010101010001: color_data = Z;
		19'b0101100010101010010: color_data = Z;
		19'b0101100010101010011: color_data = Z;
		19'b0101100010101010100: color_data = Z;
		19'b0101100010101010101: color_data = Z;
		19'b0101100010101010110: color_data = Z;
		19'b0101100010101010111: color_data = Z;
		19'b0101100010101011000: color_data = Z;
		19'b0101100010101011001: color_data = Z;
		19'b0101100010101011010: color_data = Z;
		19'b0101100010101011011: color_data = Z;
		19'b0101100010101011100: color_data = Z;
		19'b0101100010101011101: color_data = Z;
		19'b0101100010101011110: color_data = Z;
		19'b0101100010101011111: color_data = Z;
		19'b0101100010101100000: color_data = Z;
		19'b0101100010101100001: color_data = Z;
		19'b0101100010101100010: color_data = Z;
		19'b0101100010101100011: color_data = Z;
		19'b0101100010101100100: color_data = Z;
		19'b0101100010101100101: color_data = Z;
		19'b0101100010101100110: color_data = Z;
		19'b0101100010101100111: color_data = Z;
		19'b0101100010101101000: color_data = Z;
		19'b0101100010101101001: color_data = Z;
		19'b0101100010101101010: color_data = Z;
		19'b0101100010101101011: color_data = Z;
		19'b0101100010101101100: color_data = Z;
		19'b0101100010101101101: color_data = Z;
		19'b0101100010101101110: color_data = Z;
		19'b0101100010101101111: color_data = Z;
		19'b0101100010101110000: color_data = Z;
		19'b0101100010101110001: color_data = Z;
		19'b0101100010101110010: color_data = Z;
		19'b0101100010101110011: color_data = Z;
		19'b0101100010101110101: color_data = Z;
		19'b0101100010101110110: color_data = Z;
		19'b0101100010101110111: color_data = Z;
		19'b0101100010101111000: color_data = Z;
		19'b0101100010101111001: color_data = Z;
		19'b0101100010101111010: color_data = Z;
		19'b0101100010101111011: color_data = Z;
		19'b0101100010101111100: color_data = Z;
		19'b0101100010101111101: color_data = Z;
		19'b0101100010101111110: color_data = Z;
		19'b0101100010101111111: color_data = Z;
		19'b0101100010110000000: color_data = Z;
		19'b0101100010110000001: color_data = Z;
		19'b0101100010110000010: color_data = Z;
		19'b0101100010110000011: color_data = Z;
		19'b0101100010111001111: color_data = Z;
		19'b0101100010111010000: color_data = Z;
		19'b0101100010111010001: color_data = Z;
		19'b0101100010111010010: color_data = Z;
		19'b0101100010111010011: color_data = Z;
		19'b0101100010111010100: color_data = Z;
		19'b0101100010111010101: color_data = Z;
		19'b0101100010111010110: color_data = Z;
		19'b0101100010111010111: color_data = Z;
		19'b0101100010111011000: color_data = Z;
		19'b0101100010111011001: color_data = Z;
		19'b0101100010111011010: color_data = Z;
		19'b0101100010111011011: color_data = Z;
		19'b0101100100100011111: color_data = Z;
		19'b0101100100100100000: color_data = Z;
		19'b0101100100100100001: color_data = Z;
		19'b0101100100100100010: color_data = Z;
		19'b0101100100100100011: color_data = Z;
		19'b0101100100100100110: color_data = Z;
		19'b0101100100100100111: color_data = Z;
		19'b0101100100100101000: color_data = Z;
		19'b0101100100100101001: color_data = Z;
		19'b0101100100100101010: color_data = Z;
		19'b0101100100100101011: color_data = Z;
		19'b0101100100100101100: color_data = Z;
		19'b0101100100100101101: color_data = Z;
		19'b0101100100100101110: color_data = Z;
		19'b0101100100100101111: color_data = Z;
		19'b0101100100100110000: color_data = Z;
		19'b0101100100100110001: color_data = Z;
		19'b0101100100100110010: color_data = Z;
		19'b0101100100100110011: color_data = Z;
		19'b0101100100100110100: color_data = Z;
		19'b0101100100100110101: color_data = Z;
		19'b0101100100100110110: color_data = Z;
		19'b0101100100100110111: color_data = Z;
		19'b0101100100100111000: color_data = Z;
		19'b0101100100100111001: color_data = Z;
		19'b0101100100100111010: color_data = Z;
		19'b0101100100100111011: color_data = Z;
		19'b0101100100100111100: color_data = Z;
		19'b0101100100100111101: color_data = Z;
		19'b0101100100100111110: color_data = Z;
		19'b0101100100100111111: color_data = Z;
		19'b0101100100101000000: color_data = Z;
		19'b0101100100101000001: color_data = Z;
		19'b0101100100101000010: color_data = Z;
		19'b0101100100101000011: color_data = Z;
		19'b0101100100101000100: color_data = Z;
		19'b0101100100101000101: color_data = Z;
		19'b0101100100101000110: color_data = Z;
		19'b0101100100101000111: color_data = Z;
		19'b0101100100101001000: color_data = Z;
		19'b0101100100101001001: color_data = Z;
		19'b0101100100101001010: color_data = Z;
		19'b0101100100101001011: color_data = Z;
		19'b0101100100101001100: color_data = Z;
		19'b0101100100101001101: color_data = Z;
		19'b0101100100101001110: color_data = Z;
		19'b0101100100101001111: color_data = Z;
		19'b0101100100101010000: color_data = Z;
		19'b0101100100101010001: color_data = Z;
		19'b0101100100101010010: color_data = Z;
		19'b0101100100101010011: color_data = Z;
		19'b0101100100101010100: color_data = Z;
		19'b0101100100101010101: color_data = Z;
		19'b0101100100101010110: color_data = Z;
		19'b0101100100101010111: color_data = Z;
		19'b0101100100101011000: color_data = Z;
		19'b0101100100101011001: color_data = Z;
		19'b0101100100101011010: color_data = Z;
		19'b0101100100101011011: color_data = Z;
		19'b0101100100101011100: color_data = Z;
		19'b0101100100101011101: color_data = Z;
		19'b0101100100101011110: color_data = Z;
		19'b0101100100101011111: color_data = Z;
		19'b0101100100101100000: color_data = Z;
		19'b0101100100101100001: color_data = Z;
		19'b0101100100101100010: color_data = Z;
		19'b0101100100101100011: color_data = Z;
		19'b0101100100101100100: color_data = Z;
		19'b0101100100101100101: color_data = Z;
		19'b0101100100101100110: color_data = Z;
		19'b0101100100101100111: color_data = Z;
		19'b0101100100101101000: color_data = Z;
		19'b0101100100101101001: color_data = Z;
		19'b0101100100101101010: color_data = Z;
		19'b0101100100101101011: color_data = Z;
		19'b0101100100101101100: color_data = Z;
		19'b0101100100101101101: color_data = Z;
		19'b0101100100101101110: color_data = Z;
		19'b0101100100101101111: color_data = Z;
		19'b0101100100101110000: color_data = Z;
		19'b0101100100101110001: color_data = Z;
		19'b0101100100101110010: color_data = Z;
		19'b0101100100101110011: color_data = Z;
		19'b0101100100101110111: color_data = Z;
		19'b0101100100101111000: color_data = Z;
		19'b0101100100101111010: color_data = Z;
		19'b0101100100101111011: color_data = Z;
		19'b0101100100101111100: color_data = Z;
		19'b0101100100101111101: color_data = Z;
		19'b0101100100101111110: color_data = Z;
		19'b0101100100101111111: color_data = Z;
		19'b0101100100110000000: color_data = Z;
		19'b0101100100110000001: color_data = Z;
		19'b0101100100110000010: color_data = Z;
		19'b0101100100110000011: color_data = Z;
		19'b0101100100111001111: color_data = Z;
		19'b0101100100111010000: color_data = Z;
		19'b0101100100111010001: color_data = Z;
		19'b0101100100111010010: color_data = Z;
		19'b0101100100111010011: color_data = Z;
		19'b0101100100111010100: color_data = Z;
		19'b0101100100111010101: color_data = Z;
		19'b0101100100111010110: color_data = Z;
		19'b0101100100111010111: color_data = Z;
		19'b0101100100111011000: color_data = Z;
		19'b0101100100111011001: color_data = Z;
		19'b0101100100111011010: color_data = Z;
		19'b0101100100111011011: color_data = Z;
		19'b0101100110100011111: color_data = Z;
		19'b0101100110100100000: color_data = Z;
		19'b0101100110100100001: color_data = Z;
		19'b0101100110100100010: color_data = Z;
		19'b0101100110100100011: color_data = Z;
		19'b0101100110100100100: color_data = Z;
		19'b0101100110100100110: color_data = Z;
		19'b0101100110100100111: color_data = Z;
		19'b0101100110100101000: color_data = Z;
		19'b0101100110100101001: color_data = Z;
		19'b0101100110100101010: color_data = Z;
		19'b0101100110100101011: color_data = Z;
		19'b0101100110100101100: color_data = Z;
		19'b0101100110100101101: color_data = Z;
		19'b0101100110100101110: color_data = Z;
		19'b0101100110100101111: color_data = Z;
		19'b0101100110100110000: color_data = Z;
		19'b0101100110100110001: color_data = Z;
		19'b0101100110100110010: color_data = Z;
		19'b0101100110100110011: color_data = Z;
		19'b0101100110100110100: color_data = Z;
		19'b0101100110100110101: color_data = Z;
		19'b0101100110100110110: color_data = Z;
		19'b0101100110100110111: color_data = Z;
		19'b0101100110100111000: color_data = Z;
		19'b0101100110100111001: color_data = Z;
		19'b0101100110100111010: color_data = Z;
		19'b0101100110100111011: color_data = Z;
		19'b0101100110100111100: color_data = Z;
		19'b0101100110100111101: color_data = Z;
		19'b0101100110100111110: color_data = Z;
		19'b0101100110100111111: color_data = Z;
		19'b0101100110101000000: color_data = Z;
		19'b0101100110101000001: color_data = Z;
		19'b0101100110101000010: color_data = Z;
		19'b0101100110101000011: color_data = Z;
		19'b0101100110101000100: color_data = Z;
		19'b0101100110101000101: color_data = Z;
		19'b0101100110101000110: color_data = Z;
		19'b0101100110101000111: color_data = Z;
		19'b0101100110101001000: color_data = Z;
		19'b0101100110101001001: color_data = Z;
		19'b0101100110101001010: color_data = Z;
		19'b0101100110101001011: color_data = Z;
		19'b0101100110101001100: color_data = Z;
		19'b0101100110101001101: color_data = Z;
		19'b0101100110101001110: color_data = Z;
		19'b0101100110101001111: color_data = Z;
		19'b0101100110101010000: color_data = Z;
		19'b0101100110101010001: color_data = Z;
		19'b0101100110101010010: color_data = Z;
		19'b0101100110101010011: color_data = Z;
		19'b0101100110101010100: color_data = Z;
		19'b0101100110101010101: color_data = Z;
		19'b0101100110101010110: color_data = Z;
		19'b0101100110101010111: color_data = Z;
		19'b0101100110101011000: color_data = Z;
		19'b0101100110101011001: color_data = Z;
		19'b0101100110101011010: color_data = Z;
		19'b0101100110101011011: color_data = Z;
		19'b0101100110101011100: color_data = Z;
		19'b0101100110101011101: color_data = Z;
		19'b0101100110101011110: color_data = Z;
		19'b0101100110101011111: color_data = Z;
		19'b0101100110101100000: color_data = Z;
		19'b0101100110101100001: color_data = Z;
		19'b0101100110101100010: color_data = Z;
		19'b0101100110101100011: color_data = Z;
		19'b0101100110101100100: color_data = Z;
		19'b0101100110101100101: color_data = Z;
		19'b0101100110101100110: color_data = Z;
		19'b0101100110101100111: color_data = Z;
		19'b0101100110101101000: color_data = Z;
		19'b0101100110101101001: color_data = Z;
		19'b0101100110101101010: color_data = Z;
		19'b0101100110101101011: color_data = Z;
		19'b0101100110101101100: color_data = Z;
		19'b0101100110101101101: color_data = Z;
		19'b0101100110101101110: color_data = Z;
		19'b0101100110101101111: color_data = Z;
		19'b0101100110101110000: color_data = Z;
		19'b0101100110101110001: color_data = Z;
		19'b0101100110101110010: color_data = Z;
		19'b0101100110101110011: color_data = Z;
		19'b0101100110101110111: color_data = Z;
		19'b0101100110101111000: color_data = Z;
		19'b0101100110101111010: color_data = Z;
		19'b0101100110101111011: color_data = Z;
		19'b0101100110101111100: color_data = Z;
		19'b0101100110101111101: color_data = Z;
		19'b0101100110101111110: color_data = Z;
		19'b0101100110101111111: color_data = Z;
		19'b0101100110110000000: color_data = Z;
		19'b0101100110110000001: color_data = Z;
		19'b0101100110110000010: color_data = Z;
		19'b0101100110110000011: color_data = Z;
		19'b0101100110111001111: color_data = Z;
		19'b0101100110111010000: color_data = Z;
		19'b0101100110111010001: color_data = Z;
		19'b0101100110111010010: color_data = Z;
		19'b0101100110111010011: color_data = Z;
		19'b0101100110111010100: color_data = Z;
		19'b0101100110111010101: color_data = Z;
		19'b0101100110111010110: color_data = Z;
		19'b0101100110111010111: color_data = Z;
		19'b0101100110111011000: color_data = Z;
		19'b0101100110111011001: color_data = Z;
		19'b0101100110111011010: color_data = Z;
		19'b0101100110111011011: color_data = Z;
		19'b0101101000100011111: color_data = Z;
		19'b0101101000100100000: color_data = Z;
		19'b0101101000100100001: color_data = Z;
		19'b0101101000100100010: color_data = Z;
		19'b0101101000100100011: color_data = Z;
		19'b0101101000100100100: color_data = Z;
		19'b0101101000100100110: color_data = Z;
		19'b0101101000100100111: color_data = Z;
		19'b0101101000100101000: color_data = Z;
		19'b0101101000100101001: color_data = Z;
		19'b0101101000100101010: color_data = Z;
		19'b0101101000100101011: color_data = Z;
		19'b0101101000100101100: color_data = Z;
		19'b0101101000100101101: color_data = Z;
		19'b0101101000100101110: color_data = Z;
		19'b0101101000100101111: color_data = Z;
		19'b0101101000100110000: color_data = Z;
		19'b0101101000100110001: color_data = Z;
		19'b0101101000100110010: color_data = Z;
		19'b0101101000100110011: color_data = Z;
		19'b0101101000100110100: color_data = Z;
		19'b0101101000100110101: color_data = Z;
		19'b0101101000100110110: color_data = Z;
		19'b0101101000100110111: color_data = Z;
		19'b0101101000100111000: color_data = Z;
		19'b0101101000100111001: color_data = Z;
		19'b0101101000100111010: color_data = Z;
		19'b0101101000100111011: color_data = Z;
		19'b0101101000100111100: color_data = Z;
		19'b0101101000100111101: color_data = Z;
		19'b0101101000100111110: color_data = Z;
		19'b0101101000100111111: color_data = Z;
		19'b0101101000101000000: color_data = Z;
		19'b0101101000101000001: color_data = Z;
		19'b0101101000101000010: color_data = Z;
		19'b0101101000101000011: color_data = Z;
		19'b0101101000101000100: color_data = Z;
		19'b0101101000101000101: color_data = Z;
		19'b0101101000101000110: color_data = Z;
		19'b0101101000101000111: color_data = Z;
		19'b0101101000101001000: color_data = Z;
		19'b0101101000101001001: color_data = Z;
		19'b0101101000101001010: color_data = Z;
		19'b0101101000101001011: color_data = Z;
		19'b0101101000101001100: color_data = Z;
		19'b0101101000101001101: color_data = Z;
		19'b0101101000101001110: color_data = Z;
		19'b0101101000101001111: color_data = Z;
		19'b0101101000101010000: color_data = Z;
		19'b0101101000101010001: color_data = Z;
		19'b0101101000101010010: color_data = Z;
		19'b0101101000101010011: color_data = Z;
		19'b0101101000101010100: color_data = Z;
		19'b0101101000101010101: color_data = Z;
		19'b0101101000101010110: color_data = Z;
		19'b0101101000101010111: color_data = Z;
		19'b0101101000101011000: color_data = Z;
		19'b0101101000101011001: color_data = Z;
		19'b0101101000101011010: color_data = Z;
		19'b0101101000101011011: color_data = Z;
		19'b0101101000101011100: color_data = Z;
		19'b0101101000101011101: color_data = Z;
		19'b0101101000101011110: color_data = Z;
		19'b0101101000101011111: color_data = Z;
		19'b0101101000101100000: color_data = Z;
		19'b0101101000101100001: color_data = Z;
		19'b0101101000101100010: color_data = Z;
		19'b0101101000101100011: color_data = Z;
		19'b0101101000101100100: color_data = Z;
		19'b0101101000101100101: color_data = Z;
		19'b0101101000101100110: color_data = Z;
		19'b0101101000101100111: color_data = Z;
		19'b0101101000101101000: color_data = Z;
		19'b0101101000101101001: color_data = Z;
		19'b0101101000101101010: color_data = Z;
		19'b0101101000101101011: color_data = Z;
		19'b0101101000101101100: color_data = Z;
		19'b0101101000101101101: color_data = Z;
		19'b0101101000101101110: color_data = Z;
		19'b0101101000101101111: color_data = Z;
		19'b0101101000101110000: color_data = Z;
		19'b0101101000101110001: color_data = Z;
		19'b0101101000101110010: color_data = Z;
		19'b0101101000101110011: color_data = Z;
		19'b0101101000101110111: color_data = Z;
		19'b0101101000101111000: color_data = Z;
		19'b0101101000101111011: color_data = Z;
		19'b0101101000101111100: color_data = Z;
		19'b0101101000101111101: color_data = Z;
		19'b0101101000101111110: color_data = Z;
		19'b0101101000101111111: color_data = Z;
		19'b0101101000110000000: color_data = Z;
		19'b0101101000110000001: color_data = Z;
		19'b0101101000110000010: color_data = Z;
		19'b0101101000110000011: color_data = Z;
		19'b0101101000111001111: color_data = Z;
		19'b0101101000111010000: color_data = Z;
		19'b0101101000111010001: color_data = Z;
		19'b0101101000111010010: color_data = Z;
		19'b0101101000111010011: color_data = Z;
		19'b0101101000111010100: color_data = Z;
		19'b0101101000111010101: color_data = Z;
		19'b0101101000111010110: color_data = Z;
		19'b0101101000111010111: color_data = Z;
		19'b0101101000111011000: color_data = Z;
		19'b0101101000111011001: color_data = Z;
		19'b0101101000111011010: color_data = Z;
		19'b0101101000111011011: color_data = Z;
		19'b0101101010100011111: color_data = Z;
		19'b0101101010100100000: color_data = Z;
		19'b0101101010100100001: color_data = Z;
		19'b0101101010100100010: color_data = Z;
		19'b0101101010100100011: color_data = Z;
		19'b0101101010100100110: color_data = Z;
		19'b0101101010100100111: color_data = Z;
		19'b0101101010100101000: color_data = Z;
		19'b0101101010100101001: color_data = Z;
		19'b0101101010100101010: color_data = Z;
		19'b0101101010100101011: color_data = Z;
		19'b0101101010100101100: color_data = Z;
		19'b0101101010100101101: color_data = Z;
		19'b0101101010100101110: color_data = Z;
		19'b0101101010100101111: color_data = Z;
		19'b0101101010100110000: color_data = Z;
		19'b0101101010100110001: color_data = Z;
		19'b0101101010100110010: color_data = Z;
		19'b0101101010100110011: color_data = Z;
		19'b0101101010100110100: color_data = Z;
		19'b0101101010100110101: color_data = Z;
		19'b0101101010100110110: color_data = Z;
		19'b0101101010100110111: color_data = Z;
		19'b0101101010100111000: color_data = Z;
		19'b0101101010100111001: color_data = Z;
		19'b0101101010100111010: color_data = Z;
		19'b0101101010100111011: color_data = Z;
		19'b0101101010100111100: color_data = Z;
		19'b0101101010100111101: color_data = Z;
		19'b0101101010100111110: color_data = Z;
		19'b0101101010100111111: color_data = Z;
		19'b0101101010101000000: color_data = Z;
		19'b0101101010101000001: color_data = Z;
		19'b0101101010101000010: color_data = Z;
		19'b0101101010101000011: color_data = Z;
		19'b0101101010101000100: color_data = Z;
		19'b0101101010101000101: color_data = Z;
		19'b0101101010101000110: color_data = Z;
		19'b0101101010101000111: color_data = Z;
		19'b0101101010101001000: color_data = Z;
		19'b0101101010101001001: color_data = Z;
		19'b0101101010101001010: color_data = Z;
		19'b0101101010101001011: color_data = Z;
		19'b0101101010101001100: color_data = Z;
		19'b0101101010101001101: color_data = Z;
		19'b0101101010101001110: color_data = Z;
		19'b0101101010101001111: color_data = Z;
		19'b0101101010101010000: color_data = Z;
		19'b0101101010101010001: color_data = Z;
		19'b0101101010101010010: color_data = Z;
		19'b0101101010101010011: color_data = Z;
		19'b0101101010101010100: color_data = Z;
		19'b0101101010101010101: color_data = Z;
		19'b0101101010101010110: color_data = Z;
		19'b0101101010101010111: color_data = Z;
		19'b0101101010101011000: color_data = Z;
		19'b0101101010101011001: color_data = Z;
		19'b0101101010101011010: color_data = Z;
		19'b0101101010101011011: color_data = Z;
		19'b0101101010101011100: color_data = Z;
		19'b0101101010101011101: color_data = Z;
		19'b0101101010101011110: color_data = Z;
		19'b0101101010101011111: color_data = Z;
		19'b0101101010101100000: color_data = Z;
		19'b0101101010101100001: color_data = Z;
		19'b0101101010101100010: color_data = Z;
		19'b0101101010101100011: color_data = Z;
		19'b0101101010101100100: color_data = Z;
		19'b0101101010101100101: color_data = Z;
		19'b0101101010101100110: color_data = Z;
		19'b0101101010101100111: color_data = Z;
		19'b0101101010101101000: color_data = Z;
		19'b0101101010101101001: color_data = Z;
		19'b0101101010101101010: color_data = Z;
		19'b0101101010101101011: color_data = Z;
		19'b0101101010101101100: color_data = Z;
		19'b0101101010101101101: color_data = Z;
		19'b0101101010101101110: color_data = Z;
		19'b0101101010101101111: color_data = Z;
		19'b0101101010101110000: color_data = Z;
		19'b0101101010101110001: color_data = Z;
		19'b0101101010101110010: color_data = Z;
		19'b0101101010101110011: color_data = Z;
		19'b0101101010101110111: color_data = Z;
		19'b0101101010101111000: color_data = Z;
		19'b0101101010101111011: color_data = Z;
		19'b0101101010101111100: color_data = Z;
		19'b0101101010101111101: color_data = Z;
		19'b0101101010101111110: color_data = Z;
		19'b0101101010101111111: color_data = Z;
		19'b0101101010110000000: color_data = Z;
		19'b0101101010110000001: color_data = Z;
		19'b0101101010110000010: color_data = Z;
		19'b0101101010110000011: color_data = Z;
		19'b0101101010111001111: color_data = Z;
		19'b0101101010111010000: color_data = Z;
		19'b0101101010111010001: color_data = Z;
		19'b0101101010111010010: color_data = Z;
		19'b0101101010111010011: color_data = Z;
		19'b0101101010111010100: color_data = Z;
		19'b0101101010111010101: color_data = Z;
		19'b0101101010111010110: color_data = Z;
		19'b0101101010111010111: color_data = Z;
		19'b0101101010111011000: color_data = Z;
		19'b0101101010111011001: color_data = Z;
		19'b0101101010111011010: color_data = Z;
		19'b0101101010111011011: color_data = Z;
		19'b0101101100100011111: color_data = Z;
		19'b0101101100100100000: color_data = Z;
		19'b0101101100100100001: color_data = Z;
		19'b0101101100100100010: color_data = Z;
		19'b0101101100100100011: color_data = Z;
		19'b0101101100100100110: color_data = Z;
		19'b0101101100100100111: color_data = Z;
		19'b0101101100100101000: color_data = Z;
		19'b0101101100100101001: color_data = Z;
		19'b0101101100100101010: color_data = Z;
		19'b0101101100100101011: color_data = Z;
		19'b0101101100100101100: color_data = Z;
		19'b0101101100100101101: color_data = Z;
		19'b0101101100100101110: color_data = Z;
		19'b0101101100100101111: color_data = Z;
		19'b0101101100100110000: color_data = Z;
		19'b0101101100100110001: color_data = Z;
		19'b0101101100100110010: color_data = Z;
		19'b0101101100100110011: color_data = Z;
		19'b0101101100100110100: color_data = Z;
		19'b0101101100100110101: color_data = Z;
		19'b0101101100100110110: color_data = Z;
		19'b0101101100100110111: color_data = Z;
		19'b0101101100100111000: color_data = Z;
		19'b0101101100100111001: color_data = Z;
		19'b0101101100100111010: color_data = Z;
		19'b0101101100100111011: color_data = Z;
		19'b0101101100100111100: color_data = Z;
		19'b0101101100100111101: color_data = Z;
		19'b0101101100100111110: color_data = Z;
		19'b0101101100100111111: color_data = Z;
		19'b0101101100101000000: color_data = Z;
		19'b0101101100101000001: color_data = Z;
		19'b0101101100101000010: color_data = Z;
		19'b0101101100101000011: color_data = Z;
		19'b0101101100101000100: color_data = Z;
		19'b0101101100101000101: color_data = Z;
		19'b0101101100101000110: color_data = Z;
		19'b0101101100101000111: color_data = Z;
		19'b0101101100101001000: color_data = Z;
		19'b0101101100101001001: color_data = Z;
		19'b0101101100101001010: color_data = Z;
		19'b0101101100101001011: color_data = Z;
		19'b0101101100101001100: color_data = Z;
		19'b0101101100101001101: color_data = Z;
		19'b0101101100101001110: color_data = Z;
		19'b0101101100101001111: color_data = Z;
		19'b0101101100101010000: color_data = Z;
		19'b0101101100101010001: color_data = Z;
		19'b0101101100101010010: color_data = Z;
		19'b0101101100101010011: color_data = Z;
		19'b0101101100101010100: color_data = Z;
		19'b0101101100101010101: color_data = Z;
		19'b0101101100101010110: color_data = Z;
		19'b0101101100101010111: color_data = Z;
		19'b0101101100101011000: color_data = Z;
		19'b0101101100101011001: color_data = Z;
		19'b0101101100101011010: color_data = Z;
		19'b0101101100101011011: color_data = Z;
		19'b0101101100101011100: color_data = Z;
		19'b0101101100101011101: color_data = Z;
		19'b0101101100101011110: color_data = Z;
		19'b0101101100101011111: color_data = Z;
		19'b0101101100101100000: color_data = Z;
		19'b0101101100101100001: color_data = Z;
		19'b0101101100101100010: color_data = Z;
		19'b0101101100101100011: color_data = Z;
		19'b0101101100101100100: color_data = Z;
		19'b0101101100101100101: color_data = Z;
		19'b0101101100101100110: color_data = Z;
		19'b0101101100101100111: color_data = Z;
		19'b0101101100101101000: color_data = Z;
		19'b0101101100101101001: color_data = Z;
		19'b0101101100101101010: color_data = Z;
		19'b0101101100101101011: color_data = Z;
		19'b0101101100101101100: color_data = Z;
		19'b0101101100101101101: color_data = Z;
		19'b0101101100101101110: color_data = Z;
		19'b0101101100101101111: color_data = Z;
		19'b0101101100101110000: color_data = Z;
		19'b0101101100101110001: color_data = Z;
		19'b0101101100101110010: color_data = Z;
		19'b0101101100101110011: color_data = Z;
		19'b0101101100101110111: color_data = Z;
		19'b0101101100101111000: color_data = Z;
		19'b0101101100101111001: color_data = Z;
		19'b0101101100101111100: color_data = Z;
		19'b0101101100101111101: color_data = Z;
		19'b0101101100101111110: color_data = Z;
		19'b0101101100101111111: color_data = Z;
		19'b0101101100110000000: color_data = Z;
		19'b0101101100110000001: color_data = Z;
		19'b0101101100110000010: color_data = Z;
		19'b0101101100110000011: color_data = Z;
		19'b0101101100110000100: color_data = Z;
		19'b0101101100111001111: color_data = Z;
		19'b0101101100111010000: color_data = Z;
		19'b0101101100111010001: color_data = Z;
		19'b0101101100111010010: color_data = Z;
		19'b0101101100111010011: color_data = Z;
		19'b0101101100111010100: color_data = Z;
		19'b0101101100111010101: color_data = Z;
		19'b0101101100111010110: color_data = Z;
		19'b0101101100111010111: color_data = Z;
		19'b0101101100111011000: color_data = Z;
		19'b0101101100111011001: color_data = Z;
		19'b0101101100111011010: color_data = Z;
		19'b0101101100111011011: color_data = Z;
		19'b0101101110100011111: color_data = Z;
		19'b0101101110100100000: color_data = Z;
		19'b0101101110100100001: color_data = Z;
		19'b0101101110100100010: color_data = Z;
		19'b0101101110100100011: color_data = Z;
		19'b0101101110100100110: color_data = Z;
		19'b0101101110100100111: color_data = Z;
		19'b0101101110100101000: color_data = Z;
		19'b0101101110100101001: color_data = Z;
		19'b0101101110100101010: color_data = Z;
		19'b0101101110100101011: color_data = Z;
		19'b0101101110100101100: color_data = Z;
		19'b0101101110100101101: color_data = Z;
		19'b0101101110100101110: color_data = Z;
		19'b0101101110100101111: color_data = Z;
		19'b0101101110100110000: color_data = Z;
		19'b0101101110100110001: color_data = Z;
		19'b0101101110100110010: color_data = Z;
		19'b0101101110100110011: color_data = Z;
		19'b0101101110100110100: color_data = Z;
		19'b0101101110100110101: color_data = Z;
		19'b0101101110100110110: color_data = Z;
		19'b0101101110100110111: color_data = Z;
		19'b0101101110100111000: color_data = Z;
		19'b0101101110100111001: color_data = Z;
		19'b0101101110100111010: color_data = Z;
		19'b0101101110100111011: color_data = Z;
		19'b0101101110100111100: color_data = Z;
		19'b0101101110100111101: color_data = Z;
		19'b0101101110100111110: color_data = Z;
		19'b0101101110100111111: color_data = Z;
		19'b0101101110101000000: color_data = Z;
		19'b0101101110101000001: color_data = Z;
		19'b0101101110101000010: color_data = Z;
		19'b0101101110101000011: color_data = Z;
		19'b0101101110101000100: color_data = Z;
		19'b0101101110101000101: color_data = Z;
		19'b0101101110101000110: color_data = Z;
		19'b0101101110101000111: color_data = Z;
		19'b0101101110101001000: color_data = Z;
		19'b0101101110101001001: color_data = Z;
		19'b0101101110101001010: color_data = Z;
		19'b0101101110101001011: color_data = Z;
		19'b0101101110101001100: color_data = Z;
		19'b0101101110101001101: color_data = Z;
		19'b0101101110101001110: color_data = Z;
		19'b0101101110101001111: color_data = Z;
		19'b0101101110101010000: color_data = Z;
		19'b0101101110101010001: color_data = Z;
		19'b0101101110101010010: color_data = Z;
		19'b0101101110101010011: color_data = Z;
		19'b0101101110101010100: color_data = Z;
		19'b0101101110101010101: color_data = Z;
		19'b0101101110101010110: color_data = Z;
		19'b0101101110101010111: color_data = Z;
		19'b0101101110101011000: color_data = Z;
		19'b0101101110101011001: color_data = Z;
		19'b0101101110101011010: color_data = Z;
		19'b0101101110101011011: color_data = Z;
		19'b0101101110101011100: color_data = Z;
		19'b0101101110101011101: color_data = Z;
		19'b0101101110101011110: color_data = Z;
		19'b0101101110101011111: color_data = Z;
		19'b0101101110101100000: color_data = Z;
		19'b0101101110101100001: color_data = Z;
		19'b0101101110101100010: color_data = Z;
		19'b0101101110101100011: color_data = Z;
		19'b0101101110101100100: color_data = Z;
		19'b0101101110101100101: color_data = Z;
		19'b0101101110101100110: color_data = Z;
		19'b0101101110101100111: color_data = Z;
		19'b0101101110101101000: color_data = Z;
		19'b0101101110101101001: color_data = Z;
		19'b0101101110101101010: color_data = Z;
		19'b0101101110101101011: color_data = Z;
		19'b0101101110101101100: color_data = Z;
		19'b0101101110101101101: color_data = Z;
		19'b0101101110101101110: color_data = Z;
		19'b0101101110101101111: color_data = Z;
		19'b0101101110101110000: color_data = Z;
		19'b0101101110101110001: color_data = Z;
		19'b0101101110101110010: color_data = Z;
		19'b0101101110101110011: color_data = Z;
		19'b0101101110101110111: color_data = Z;
		19'b0101101110101111000: color_data = Z;
		19'b0101101110101111101: color_data = Z;
		19'b0101101110101111110: color_data = Z;
		19'b0101101110101111111: color_data = Z;
		19'b0101101110110000000: color_data = Z;
		19'b0101101110110000001: color_data = Z;
		19'b0101101110110000010: color_data = Z;
		19'b0101101110110000011: color_data = Z;
		19'b0101101110110000100: color_data = Z;
		19'b0101101110111001111: color_data = Z;
		19'b0101101110111010000: color_data = Z;
		19'b0101101110111010001: color_data = Z;
		19'b0101101110111010010: color_data = Z;
		19'b0101101110111010011: color_data = Z;
		19'b0101101110111010100: color_data = Z;
		19'b0101101110111010101: color_data = Z;
		19'b0101101110111010110: color_data = Z;
		19'b0101101110111010111: color_data = Z;
		19'b0101101110111011000: color_data = Z;
		19'b0101101110111011001: color_data = Z;
		19'b0101101110111011010: color_data = Z;
		19'b0101101110111011011: color_data = Z;
		19'b0101110000100011111: color_data = Z;
		19'b0101110000100100000: color_data = Z;
		19'b0101110000100100001: color_data = Z;
		19'b0101110000100100010: color_data = Z;
		19'b0101110000100100011: color_data = Z;
		19'b0101110000100100110: color_data = Z;
		19'b0101110000100100111: color_data = Z;
		19'b0101110000100101000: color_data = Z;
		19'b0101110000100101001: color_data = Z;
		19'b0101110000100101010: color_data = Z;
		19'b0101110000100101011: color_data = Z;
		19'b0101110000100101100: color_data = Z;
		19'b0101110000100101101: color_data = Z;
		19'b0101110000100101110: color_data = Z;
		19'b0101110000100101111: color_data = Z;
		19'b0101110000100110000: color_data = Z;
		19'b0101110000100110001: color_data = Z;
		19'b0101110000100110010: color_data = Z;
		19'b0101110000100110011: color_data = Z;
		19'b0101110000100110100: color_data = Z;
		19'b0101110000100110101: color_data = Z;
		19'b0101110000100110110: color_data = Z;
		19'b0101110000100110111: color_data = Z;
		19'b0101110000100111000: color_data = Z;
		19'b0101110000100111001: color_data = Z;
		19'b0101110000100111010: color_data = Z;
		19'b0101110000100111011: color_data = Z;
		19'b0101110000100111100: color_data = Z;
		19'b0101110000100111101: color_data = Z;
		19'b0101110000100111110: color_data = Z;
		19'b0101110000100111111: color_data = Z;
		19'b0101110000101000000: color_data = Z;
		19'b0101110000101000001: color_data = Z;
		19'b0101110000101000010: color_data = Z;
		19'b0101110000101000011: color_data = Z;
		19'b0101110000101000100: color_data = Z;
		19'b0101110000101000101: color_data = Z;
		19'b0101110000101000110: color_data = Z;
		19'b0101110000101000111: color_data = Z;
		19'b0101110000101001000: color_data = Z;
		19'b0101110000101001001: color_data = Z;
		19'b0101110000101001010: color_data = Z;
		19'b0101110000101001011: color_data = Z;
		19'b0101110000101001100: color_data = Z;
		19'b0101110000101001101: color_data = Z;
		19'b0101110000101001110: color_data = Z;
		19'b0101110000101001111: color_data = Z;
		19'b0101110000101010000: color_data = Z;
		19'b0101110000101010001: color_data = Z;
		19'b0101110000101010010: color_data = Z;
		19'b0101110000101010011: color_data = Z;
		19'b0101110000101010100: color_data = Z;
		19'b0101110000101010101: color_data = Z;
		19'b0101110000101010110: color_data = Z;
		19'b0101110000101010111: color_data = Z;
		19'b0101110000101011000: color_data = Z;
		19'b0101110000101011001: color_data = Z;
		19'b0101110000101011010: color_data = Z;
		19'b0101110000101011011: color_data = Z;
		19'b0101110000101011100: color_data = Z;
		19'b0101110000101011101: color_data = Z;
		19'b0101110000101011110: color_data = Z;
		19'b0101110000101011111: color_data = Z;
		19'b0101110000101100000: color_data = Z;
		19'b0101110000101100001: color_data = Z;
		19'b0101110000101100010: color_data = Z;
		19'b0101110000101100011: color_data = Z;
		19'b0101110000101100100: color_data = Z;
		19'b0101110000101100101: color_data = Z;
		19'b0101110000101100110: color_data = Z;
		19'b0101110000101100111: color_data = Z;
		19'b0101110000101101000: color_data = Z;
		19'b0101110000101101001: color_data = Z;
		19'b0101110000101101010: color_data = Z;
		19'b0101110000101101011: color_data = Z;
		19'b0101110000101101100: color_data = Z;
		19'b0101110000101101101: color_data = Z;
		19'b0101110000101101110: color_data = Z;
		19'b0101110000101101111: color_data = Z;
		19'b0101110000101110000: color_data = Z;
		19'b0101110000101110001: color_data = Z;
		19'b0101110000101110010: color_data = Z;
		19'b0101110000101110011: color_data = Z;
		19'b0101110000101111000: color_data = Z;
		19'b0101110000101111110: color_data = Z;
		19'b0101110000101111111: color_data = Z;
		19'b0101110000110000000: color_data = Z;
		19'b0101110000110000001: color_data = Z;
		19'b0101110000110000010: color_data = Z;
		19'b0101110000110000011: color_data = Z;
		19'b0101110000110000100: color_data = Z;
		19'b0101110000111010000: color_data = Z;
		19'b0101110000111010001: color_data = Z;
		19'b0101110000111010010: color_data = Z;
		19'b0101110000111010011: color_data = Z;
		19'b0101110000111010100: color_data = Z;
		19'b0101110000111010101: color_data = Z;
		19'b0101110000111010110: color_data = Z;
		19'b0101110000111010111: color_data = Z;
		19'b0101110000111011000: color_data = Z;
		19'b0101110000111011001: color_data = Z;
		19'b0101110000111011010: color_data = Z;
		19'b0101110000111011011: color_data = Z;
		19'b0101110010100011111: color_data = Z;
		19'b0101110010100100000: color_data = Z;
		19'b0101110010100100001: color_data = Z;
		19'b0101110010100100010: color_data = Z;
		19'b0101110010100100011: color_data = Z;
		19'b0101110010100100110: color_data = Z;
		19'b0101110010100100111: color_data = Z;
		19'b0101110010100101000: color_data = Z;
		19'b0101110010100101001: color_data = Z;
		19'b0101110010100101010: color_data = Z;
		19'b0101110010100101011: color_data = Z;
		19'b0101110010100101100: color_data = Z;
		19'b0101110010100101101: color_data = Z;
		19'b0101110010100101110: color_data = Z;
		19'b0101110010100101111: color_data = Z;
		19'b0101110010100110000: color_data = Z;
		19'b0101110010100110001: color_data = Z;
		19'b0101110010100110010: color_data = Z;
		19'b0101110010100110011: color_data = Z;
		19'b0101110010100110100: color_data = Z;
		19'b0101110010100110101: color_data = Z;
		19'b0101110010100110110: color_data = Z;
		19'b0101110010100110111: color_data = Z;
		19'b0101110010100111000: color_data = Z;
		19'b0101110010100111001: color_data = Z;
		19'b0101110010100111010: color_data = Z;
		19'b0101110010100111011: color_data = Z;
		19'b0101110010100111100: color_data = Z;
		19'b0101110010100111101: color_data = Z;
		19'b0101110010100111110: color_data = Z;
		19'b0101110010100111111: color_data = Z;
		19'b0101110010101000000: color_data = Z;
		19'b0101110010101000001: color_data = Z;
		19'b0101110010101000010: color_data = Z;
		19'b0101110010101000011: color_data = Z;
		19'b0101110010101000100: color_data = Z;
		19'b0101110010101000101: color_data = Z;
		19'b0101110010101000110: color_data = Z;
		19'b0101110010101000111: color_data = Z;
		19'b0101110010101001000: color_data = Z;
		19'b0101110010101001001: color_data = Z;
		19'b0101110010101001010: color_data = Z;
		19'b0101110010101001011: color_data = Z;
		19'b0101110010101001100: color_data = Z;
		19'b0101110010101001101: color_data = Z;
		19'b0101110010101001110: color_data = Z;
		19'b0101110010101001111: color_data = Z;
		19'b0101110010101010000: color_data = Z;
		19'b0101110010101010001: color_data = Z;
		19'b0101110010101010010: color_data = Z;
		19'b0101110010101010011: color_data = Z;
		19'b0101110010101010100: color_data = Z;
		19'b0101110010101010101: color_data = Z;
		19'b0101110010101010110: color_data = Z;
		19'b0101110010101010111: color_data = Z;
		19'b0101110010101011000: color_data = Z;
		19'b0101110010101011001: color_data = Z;
		19'b0101110010101011010: color_data = Z;
		19'b0101110010101011011: color_data = Z;
		19'b0101110010101011100: color_data = Z;
		19'b0101110010101011101: color_data = Z;
		19'b0101110010101011110: color_data = Z;
		19'b0101110010101011111: color_data = Z;
		19'b0101110010101100000: color_data = Z;
		19'b0101110010101100001: color_data = Z;
		19'b0101110010101100010: color_data = Z;
		19'b0101110010101100011: color_data = Z;
		19'b0101110010101100100: color_data = Z;
		19'b0101110010101100101: color_data = Z;
		19'b0101110010101100110: color_data = Z;
		19'b0101110010101100111: color_data = Z;
		19'b0101110010101101000: color_data = Z;
		19'b0101110010101101001: color_data = Z;
		19'b0101110010101101010: color_data = Z;
		19'b0101110010101101011: color_data = Z;
		19'b0101110010101101100: color_data = Z;
		19'b0101110010101101101: color_data = Z;
		19'b0101110010101101110: color_data = Z;
		19'b0101110010101101111: color_data = Z;
		19'b0101110010101110000: color_data = Z;
		19'b0101110010101110001: color_data = Z;
		19'b0101110010101110010: color_data = Z;
		19'b0101110010101110011: color_data = Z;
		19'b0101110010101111000: color_data = Z;
		19'b0101110010101111110: color_data = Z;
		19'b0101110010101111111: color_data = Z;
		19'b0101110010110000000: color_data = Z;
		19'b0101110010110000001: color_data = Z;
		19'b0101110010110000010: color_data = Z;
		19'b0101110010110000011: color_data = Z;
		19'b0101110010110000100: color_data = Z;
		19'b0101110010110000101: color_data = Z;
		19'b0101110010111010000: color_data = Z;
		19'b0101110010111010001: color_data = Z;
		19'b0101110010111010010: color_data = Z;
		19'b0101110010111010011: color_data = Z;
		19'b0101110010111010100: color_data = Z;
		19'b0101110010111010101: color_data = Z;
		19'b0101110010111010110: color_data = Z;
		19'b0101110010111010111: color_data = Z;
		19'b0101110010111011000: color_data = Z;
		19'b0101110010111011001: color_data = Z;
		19'b0101110010111011010: color_data = Z;
		19'b0101110010111011011: color_data = Z;
		19'b0101110100100011110: color_data = Z;
		19'b0101110100100011111: color_data = Z;
		19'b0101110100100100000: color_data = Z;
		19'b0101110100100100001: color_data = Z;
		19'b0101110100100100010: color_data = Z;
		19'b0101110100100100011: color_data = Z;
		19'b0101110100100100110: color_data = Z;
		19'b0101110100100100111: color_data = Z;
		19'b0101110100100101000: color_data = Z;
		19'b0101110100100101001: color_data = Z;
		19'b0101110100100101010: color_data = Z;
		19'b0101110100100101011: color_data = Z;
		19'b0101110100100101100: color_data = Z;
		19'b0101110100100101101: color_data = Z;
		19'b0101110100100101110: color_data = Z;
		19'b0101110100100101111: color_data = Z;
		19'b0101110100100110000: color_data = Z;
		19'b0101110100100110001: color_data = Z;
		19'b0101110100100110010: color_data = Z;
		19'b0101110100100110011: color_data = Z;
		19'b0101110100100110100: color_data = Z;
		19'b0101110100100110101: color_data = Z;
		19'b0101110100100110110: color_data = Z;
		19'b0101110100100110111: color_data = Z;
		19'b0101110100100111000: color_data = Z;
		19'b0101110100100111001: color_data = Z;
		19'b0101110100100111010: color_data = Z;
		19'b0101110100100111011: color_data = Z;
		19'b0101110100100111100: color_data = Z;
		19'b0101110100100111101: color_data = Z;
		19'b0101110100100111110: color_data = Z;
		19'b0101110100100111111: color_data = Z;
		19'b0101110100101000000: color_data = Z;
		19'b0101110100101000001: color_data = Z;
		19'b0101110100101000010: color_data = Z;
		19'b0101110100101000011: color_data = Z;
		19'b0101110100101000100: color_data = Z;
		19'b0101110100101000101: color_data = Z;
		19'b0101110100101000110: color_data = Z;
		19'b0101110100101000111: color_data = Z;
		19'b0101110100101001000: color_data = Z;
		19'b0101110100101001001: color_data = Z;
		19'b0101110100101001010: color_data = Z;
		19'b0101110100101001011: color_data = Z;
		19'b0101110100101001100: color_data = Z;
		19'b0101110100101001101: color_data = Z;
		19'b0101110100101001110: color_data = Z;
		19'b0101110100101001111: color_data = Z;
		19'b0101110100101010000: color_data = Z;
		19'b0101110100101010001: color_data = Z;
		19'b0101110100101010010: color_data = Z;
		19'b0101110100101010011: color_data = Z;
		19'b0101110100101010100: color_data = Z;
		19'b0101110100101010101: color_data = Z;
		19'b0101110100101010110: color_data = Z;
		19'b0101110100101010111: color_data = Z;
		19'b0101110100101011000: color_data = Z;
		19'b0101110100101011001: color_data = Z;
		19'b0101110100101011010: color_data = Z;
		19'b0101110100101011011: color_data = Z;
		19'b0101110100101011100: color_data = Z;
		19'b0101110100101011101: color_data = Z;
		19'b0101110100101011110: color_data = Z;
		19'b0101110100101011111: color_data = Z;
		19'b0101110100101100000: color_data = Z;
		19'b0101110100101100001: color_data = Z;
		19'b0101110100101100010: color_data = Z;
		19'b0101110100101100011: color_data = Z;
		19'b0101110100101100100: color_data = Z;
		19'b0101110100101100101: color_data = Z;
		19'b0101110100101100110: color_data = Z;
		19'b0101110100101100111: color_data = Z;
		19'b0101110100101101000: color_data = Z;
		19'b0101110100101101001: color_data = Z;
		19'b0101110100101101010: color_data = Z;
		19'b0101110100101101011: color_data = Z;
		19'b0101110100101101100: color_data = Z;
		19'b0101110100101101101: color_data = Z;
		19'b0101110100101101110: color_data = Z;
		19'b0101110100101101111: color_data = Z;
		19'b0101110100101110000: color_data = Z;
		19'b0101110100101110001: color_data = Z;
		19'b0101110100101110010: color_data = Z;
		19'b0101110100101110011: color_data = Z;
		19'b0101110100101111000: color_data = Z;
		19'b0101110100101111001: color_data = Z;
		19'b0101110100101111111: color_data = Z;
		19'b0101110100110000000: color_data = Z;
		19'b0101110100110000001: color_data = Z;
		19'b0101110100110000010: color_data = Z;
		19'b0101110100110000011: color_data = Z;
		19'b0101110100110000100: color_data = Z;
		19'b0101110100110000101: color_data = Z;
		19'b0101110100111010000: color_data = Z;
		19'b0101110100111010001: color_data = Z;
		19'b0101110100111010010: color_data = Z;
		19'b0101110100111010011: color_data = Z;
		19'b0101110100111010100: color_data = Z;
		19'b0101110100111010101: color_data = Z;
		19'b0101110100111010110: color_data = Z;
		19'b0101110100111010111: color_data = Z;
		19'b0101110100111011000: color_data = Z;
		19'b0101110100111011001: color_data = Z;
		19'b0101110100111011010: color_data = Z;
		19'b0101110100111011011: color_data = Z;
		19'b0101110110100011110: color_data = Z;
		19'b0101110110100011111: color_data = Z;
		19'b0101110110100100000: color_data = Z;
		19'b0101110110100100001: color_data = Z;
		19'b0101110110100100010: color_data = Z;
		19'b0101110110100100011: color_data = Z;
		19'b0101110110100100110: color_data = Z;
		19'b0101110110100100111: color_data = Z;
		19'b0101110110100101000: color_data = Z;
		19'b0101110110100101001: color_data = Z;
		19'b0101110110100101010: color_data = Z;
		19'b0101110110100101011: color_data = Z;
		19'b0101110110100101100: color_data = Z;
		19'b0101110110100101101: color_data = Z;
		19'b0101110110100101110: color_data = Z;
		19'b0101110110100101111: color_data = Z;
		19'b0101110110100110000: color_data = Z;
		19'b0101110110100110001: color_data = Z;
		19'b0101110110100110010: color_data = Z;
		19'b0101110110100110011: color_data = Z;
		19'b0101110110100110100: color_data = Z;
		19'b0101110110100110101: color_data = Z;
		19'b0101110110100110110: color_data = Z;
		19'b0101110110100110111: color_data = Z;
		19'b0101110110100111000: color_data = Z;
		19'b0101110110100111001: color_data = Z;
		19'b0101110110100111010: color_data = Z;
		19'b0101110110100111011: color_data = Z;
		19'b0101110110100111100: color_data = Z;
		19'b0101110110100111101: color_data = Z;
		19'b0101110110100111110: color_data = Z;
		19'b0101110110100111111: color_data = Z;
		19'b0101110110101000000: color_data = Z;
		19'b0101110110101000001: color_data = Z;
		19'b0101110110101000010: color_data = Z;
		19'b0101110110101000011: color_data = Z;
		19'b0101110110101000100: color_data = Z;
		19'b0101110110101000101: color_data = Z;
		19'b0101110110101000110: color_data = Z;
		19'b0101110110101000111: color_data = Z;
		19'b0101110110101001000: color_data = Z;
		19'b0101110110101001001: color_data = Z;
		19'b0101110110101001010: color_data = Z;
		19'b0101110110101001011: color_data = Z;
		19'b0101110110101001100: color_data = Z;
		19'b0101110110101001101: color_data = Z;
		19'b0101110110101001110: color_data = Z;
		19'b0101110110101001111: color_data = Z;
		19'b0101110110101010000: color_data = Z;
		19'b0101110110101010001: color_data = Z;
		19'b0101110110101010010: color_data = Z;
		19'b0101110110101010011: color_data = Z;
		19'b0101110110101010100: color_data = Z;
		19'b0101110110101010101: color_data = Z;
		19'b0101110110101010110: color_data = Z;
		19'b0101110110101010111: color_data = Z;
		19'b0101110110101011000: color_data = Z;
		19'b0101110110101011001: color_data = Z;
		19'b0101110110101011010: color_data = Z;
		19'b0101110110101011011: color_data = Z;
		19'b0101110110101011100: color_data = Z;
		19'b0101110110101011101: color_data = Z;
		19'b0101110110101011110: color_data = Z;
		19'b0101110110101011111: color_data = Z;
		19'b0101110110101100000: color_data = Z;
		19'b0101110110101100001: color_data = Z;
		19'b0101110110101100010: color_data = Z;
		19'b0101110110101100011: color_data = Z;
		19'b0101110110101100100: color_data = Z;
		19'b0101110110101100101: color_data = Z;
		19'b0101110110101100110: color_data = Z;
		19'b0101110110101100111: color_data = Z;
		19'b0101110110101101000: color_data = Z;
		19'b0101110110101101001: color_data = Z;
		19'b0101110110101101010: color_data = Z;
		19'b0101110110101101011: color_data = Z;
		19'b0101110110101101100: color_data = Z;
		19'b0101110110101101101: color_data = Z;
		19'b0101110110101101110: color_data = Z;
		19'b0101110110101101111: color_data = Z;
		19'b0101110110101110000: color_data = Z;
		19'b0101110110101110001: color_data = Z;
		19'b0101110110101110010: color_data = Z;
		19'b0101110110101110011: color_data = Z;
		19'b0101110110101110100: color_data = Z;
		19'b0101110110101111000: color_data = Z;
		19'b0101110110101111001: color_data = Z;
		19'b0101110110110000001: color_data = Z;
		19'b0101110110110000010: color_data = Z;
		19'b0101110110110000011: color_data = Z;
		19'b0101110110110000100: color_data = Z;
		19'b0101110110110000101: color_data = Z;
		19'b0101110110110000110: color_data = Z;
		19'b0101110110111010000: color_data = Z;
		19'b0101110110111010001: color_data = Z;
		19'b0101110110111010010: color_data = Z;
		19'b0101110110111010011: color_data = Z;
		19'b0101110110111010100: color_data = Z;
		19'b0101110110111010101: color_data = Z;
		19'b0101110110111010110: color_data = Z;
		19'b0101110110111010111: color_data = Z;
		19'b0101110110111011000: color_data = Z;
		19'b0101110110111011001: color_data = Z;
		19'b0101110110111011010: color_data = Z;
		19'b0101110110111011011: color_data = Z;
		19'b0101111000100011110: color_data = Z;
		19'b0101111000100011111: color_data = Z;
		19'b0101111000100100000: color_data = Z;
		19'b0101111000100100001: color_data = Z;
		19'b0101111000100100010: color_data = Z;
		19'b0101111000100100011: color_data = Z;
		19'b0101111000100100101: color_data = Z;
		19'b0101111000100100110: color_data = Z;
		19'b0101111000100100111: color_data = Z;
		19'b0101111000100101000: color_data = Z;
		19'b0101111000100101001: color_data = Z;
		19'b0101111000100101010: color_data = Z;
		19'b0101111000100101011: color_data = Z;
		19'b0101111000100101100: color_data = Z;
		19'b0101111000100101101: color_data = Z;
		19'b0101111000100101110: color_data = Z;
		19'b0101111000100101111: color_data = Z;
		19'b0101111000100110000: color_data = Z;
		19'b0101111000100110001: color_data = Z;
		19'b0101111000100110010: color_data = Z;
		19'b0101111000100110011: color_data = Z;
		19'b0101111000100110100: color_data = Z;
		19'b0101111000100110101: color_data = Z;
		19'b0101111000100110110: color_data = Z;
		19'b0101111000100110111: color_data = Z;
		19'b0101111000100111000: color_data = Z;
		19'b0101111000100111001: color_data = Z;
		19'b0101111000100111010: color_data = Z;
		19'b0101111000100111011: color_data = Z;
		19'b0101111000100111100: color_data = Z;
		19'b0101111000100111101: color_data = Z;
		19'b0101111000100111110: color_data = Z;
		19'b0101111000100111111: color_data = Z;
		19'b0101111000101000000: color_data = Z;
		19'b0101111000101000001: color_data = Z;
		19'b0101111000101000010: color_data = Z;
		19'b0101111000101000011: color_data = Z;
		19'b0101111000101000100: color_data = Z;
		19'b0101111000101000101: color_data = Z;
		19'b0101111000101000110: color_data = Z;
		19'b0101111000101000111: color_data = Z;
		19'b0101111000101001000: color_data = Z;
		19'b0101111000101001001: color_data = Z;
		19'b0101111000101001010: color_data = Z;
		19'b0101111000101001011: color_data = Z;
		19'b0101111000101001100: color_data = Z;
		19'b0101111000101001101: color_data = Z;
		19'b0101111000101001110: color_data = Z;
		19'b0101111000101001111: color_data = Z;
		19'b0101111000101010000: color_data = Z;
		19'b0101111000101010001: color_data = Z;
		19'b0101111000101010010: color_data = Z;
		19'b0101111000101010011: color_data = Z;
		19'b0101111000101010100: color_data = Z;
		19'b0101111000101010101: color_data = Z;
		19'b0101111000101010110: color_data = Z;
		19'b0101111000101010111: color_data = Z;
		19'b0101111000101011000: color_data = Z;
		19'b0101111000101011001: color_data = Z;
		19'b0101111000101011010: color_data = Z;
		19'b0101111000101011011: color_data = Z;
		19'b0101111000101011100: color_data = Z;
		19'b0101111000101011101: color_data = Z;
		19'b0101111000101011110: color_data = Z;
		19'b0101111000101011111: color_data = Z;
		19'b0101111000101100000: color_data = Z;
		19'b0101111000101100001: color_data = Z;
		19'b0101111000101100010: color_data = Z;
		19'b0101111000101100011: color_data = Z;
		19'b0101111000101100100: color_data = Z;
		19'b0101111000101100101: color_data = Z;
		19'b0101111000101100110: color_data = Z;
		19'b0101111000101100111: color_data = Z;
		19'b0101111000101101000: color_data = Z;
		19'b0101111000101101001: color_data = Z;
		19'b0101111000101101010: color_data = Z;
		19'b0101111000101101011: color_data = Z;
		19'b0101111000101101100: color_data = Z;
		19'b0101111000101101101: color_data = Z;
		19'b0101111000101101110: color_data = Z;
		19'b0101111000101101111: color_data = Z;
		19'b0101111000101110000: color_data = Z;
		19'b0101111000101110001: color_data = Z;
		19'b0101111000101110010: color_data = Z;
		19'b0101111000101110011: color_data = Z;
		19'b0101111000101110100: color_data = Z;
		19'b0101111000101111001: color_data = Z;
		19'b0101111000110000010: color_data = Z;
		19'b0101111000110000011: color_data = Z;
		19'b0101111000110000100: color_data = Z;
		19'b0101111000110000101: color_data = Z;
		19'b0101111000110000110: color_data = Z;
		19'b0101111000110000111: color_data = Z;
		19'b0101111000111010000: color_data = Z;
		19'b0101111000111010001: color_data = Z;
		19'b0101111000111010010: color_data = Z;
		19'b0101111000111010011: color_data = Z;
		19'b0101111000111010100: color_data = Z;
		19'b0101111000111010101: color_data = Z;
		19'b0101111000111010110: color_data = Z;
		19'b0101111000111010111: color_data = Z;
		19'b0101111000111011000: color_data = Z;
		19'b0101111000111011001: color_data = Z;
		19'b0101111000111011010: color_data = Z;
		19'b0101111000111011011: color_data = Z;
		19'b0101111010100011110: color_data = Z;
		19'b0101111010100011111: color_data = Z;
		19'b0101111010100100000: color_data = Z;
		19'b0101111010100100001: color_data = Z;
		19'b0101111010100100010: color_data = Z;
		19'b0101111010100100011: color_data = Z;
		19'b0101111010100100101: color_data = Z;
		19'b0101111010100100110: color_data = Z;
		19'b0101111010100100111: color_data = Z;
		19'b0101111010100101000: color_data = Z;
		19'b0101111010100101001: color_data = Z;
		19'b0101111010100101010: color_data = Z;
		19'b0101111010100101011: color_data = Z;
		19'b0101111010100101100: color_data = Z;
		19'b0101111010100101101: color_data = Z;
		19'b0101111010100101110: color_data = Z;
		19'b0101111010100101111: color_data = Z;
		19'b0101111010100110000: color_data = Z;
		19'b0101111010100110001: color_data = Z;
		19'b0101111010100110010: color_data = Z;
		19'b0101111010100110011: color_data = Z;
		19'b0101111010100110100: color_data = Z;
		19'b0101111010100110101: color_data = Z;
		19'b0101111010100110110: color_data = Z;
		19'b0101111010100110111: color_data = Z;
		19'b0101111010100111000: color_data = Z;
		19'b0101111010100111001: color_data = Z;
		19'b0101111010100111010: color_data = Z;
		19'b0101111010100111011: color_data = Z;
		19'b0101111010100111100: color_data = Z;
		19'b0101111010100111101: color_data = Z;
		19'b0101111010100111110: color_data = Z;
		19'b0101111010100111111: color_data = Z;
		19'b0101111010101000000: color_data = Z;
		19'b0101111010101000001: color_data = Z;
		19'b0101111010101000010: color_data = Z;
		19'b0101111010101000011: color_data = Z;
		19'b0101111010101000100: color_data = Z;
		19'b0101111010101000101: color_data = Z;
		19'b0101111010101000110: color_data = Z;
		19'b0101111010101000111: color_data = Z;
		19'b0101111010101001000: color_data = Z;
		19'b0101111010101001001: color_data = Z;
		19'b0101111010101001010: color_data = Z;
		19'b0101111010101001011: color_data = Z;
		19'b0101111010101001100: color_data = Z;
		19'b0101111010101001101: color_data = Z;
		19'b0101111010101001110: color_data = Z;
		19'b0101111010101001111: color_data = Z;
		19'b0101111010101010000: color_data = Z;
		19'b0101111010101010001: color_data = Z;
		19'b0101111010101010010: color_data = Z;
		19'b0101111010101010011: color_data = Z;
		19'b0101111010101010100: color_data = Z;
		19'b0101111010101010101: color_data = Z;
		19'b0101111010101010110: color_data = Z;
		19'b0101111010101010111: color_data = Z;
		19'b0101111010101011000: color_data = Z;
		19'b0101111010101011001: color_data = Z;
		19'b0101111010101011010: color_data = Z;
		19'b0101111010101011011: color_data = Z;
		19'b0101111010101011100: color_data = Z;
		19'b0101111010101011101: color_data = Z;
		19'b0101111010101011110: color_data = Z;
		19'b0101111010101011111: color_data = Z;
		19'b0101111010101100000: color_data = Z;
		19'b0101111010101100001: color_data = Z;
		19'b0101111010101100010: color_data = Z;
		19'b0101111010101100011: color_data = Z;
		19'b0101111010101100100: color_data = Z;
		19'b0101111010101100101: color_data = Z;
		19'b0101111010101100110: color_data = Z;
		19'b0101111010101100111: color_data = Z;
		19'b0101111010101101000: color_data = Z;
		19'b0101111010101101001: color_data = Z;
		19'b0101111010101101010: color_data = Z;
		19'b0101111010101101011: color_data = Z;
		19'b0101111010101101100: color_data = Z;
		19'b0101111010101101101: color_data = Z;
		19'b0101111010101101110: color_data = Z;
		19'b0101111010101101111: color_data = Z;
		19'b0101111010101110000: color_data = Z;
		19'b0101111010101110001: color_data = Z;
		19'b0101111010101110010: color_data = Z;
		19'b0101111010101110011: color_data = Z;
		19'b0101111010101110100: color_data = Z;
		19'b0101111010110000011: color_data = Z;
		19'b0101111010110000100: color_data = Z;
		19'b0101111010110000101: color_data = Z;
		19'b0101111010110000110: color_data = Z;
		19'b0101111010110000111: color_data = Z;
		19'b0101111010111010000: color_data = Z;
		19'b0101111010111010001: color_data = Z;
		19'b0101111010111010010: color_data = Z;
		19'b0101111010111010011: color_data = Z;
		19'b0101111010111010100: color_data = Z;
		19'b0101111010111010101: color_data = Z;
		19'b0101111010111010110: color_data = Z;
		19'b0101111010111010111: color_data = Z;
		19'b0101111010111011000: color_data = Z;
		19'b0101111010111011001: color_data = Z;
		19'b0101111010111011010: color_data = Z;
		19'b0101111010111011011: color_data = Z;
		19'b0101111100100011110: color_data = Z;
		19'b0101111100100011111: color_data = Z;
		19'b0101111100100100000: color_data = Z;
		19'b0101111100100100001: color_data = Z;
		19'b0101111100100100010: color_data = Z;
		19'b0101111100100100011: color_data = Z;
		19'b0101111100100100101: color_data = Z;
		19'b0101111100100100110: color_data = Z;
		19'b0101111100100100111: color_data = Z;
		19'b0101111100100101000: color_data = Z;
		19'b0101111100100101001: color_data = Z;
		19'b0101111100100101010: color_data = Z;
		19'b0101111100100101011: color_data = Z;
		19'b0101111100100101100: color_data = Z;
		19'b0101111100100101101: color_data = Z;
		19'b0101111100100101110: color_data = Z;
		19'b0101111100100101111: color_data = Z;
		19'b0101111100100110000: color_data = Z;
		19'b0101111100100110001: color_data = Z;
		19'b0101111100100110010: color_data = Z;
		19'b0101111100100110011: color_data = Z;
		19'b0101111100100110100: color_data = Z;
		19'b0101111100100110101: color_data = Z;
		19'b0101111100100110110: color_data = Z;
		19'b0101111100100110111: color_data = Z;
		19'b0101111100100111000: color_data = Z;
		19'b0101111100100111001: color_data = Z;
		19'b0101111100100111010: color_data = Z;
		19'b0101111100100111011: color_data = Z;
		19'b0101111100100111100: color_data = Z;
		19'b0101111100100111101: color_data = Z;
		19'b0101111100100111110: color_data = Z;
		19'b0101111100100111111: color_data = Z;
		19'b0101111100101000000: color_data = Z;
		19'b0101111100101000001: color_data = Z;
		19'b0101111100101000010: color_data = Z;
		19'b0101111100101000011: color_data = Z;
		19'b0101111100101000100: color_data = Z;
		19'b0101111100101000101: color_data = Z;
		19'b0101111100101000110: color_data = Z;
		19'b0101111100101000111: color_data = Z;
		19'b0101111100101001000: color_data = Z;
		19'b0101111100101001001: color_data = Z;
		19'b0101111100101001010: color_data = Z;
		19'b0101111100101001011: color_data = Z;
		19'b0101111100101001100: color_data = Z;
		19'b0101111100101001101: color_data = Z;
		19'b0101111100101001110: color_data = Z;
		19'b0101111100101001111: color_data = Z;
		19'b0101111100101010000: color_data = Z;
		19'b0101111100101010001: color_data = Z;
		19'b0101111100101010010: color_data = Z;
		19'b0101111100101010011: color_data = Z;
		19'b0101111100101010100: color_data = Z;
		19'b0101111100101010101: color_data = Z;
		19'b0101111100101010110: color_data = Z;
		19'b0101111100101010111: color_data = Z;
		19'b0101111100101011000: color_data = Z;
		19'b0101111100101011001: color_data = Z;
		19'b0101111100101011010: color_data = Z;
		19'b0101111100101011011: color_data = Z;
		19'b0101111100101011100: color_data = Z;
		19'b0101111100101011101: color_data = Z;
		19'b0101111100101011110: color_data = Z;
		19'b0101111100101011111: color_data = Z;
		19'b0101111100101100000: color_data = Z;
		19'b0101111100101100001: color_data = Z;
		19'b0101111100101100010: color_data = Z;
		19'b0101111100101100011: color_data = Z;
		19'b0101111100101100100: color_data = Z;
		19'b0101111100101100101: color_data = Z;
		19'b0101111100101100110: color_data = Z;
		19'b0101111100101100111: color_data = Z;
		19'b0101111100101101000: color_data = Z;
		19'b0101111100101101001: color_data = Z;
		19'b0101111100101101010: color_data = Z;
		19'b0101111100101101011: color_data = Z;
		19'b0101111100101101100: color_data = Z;
		19'b0101111100101101101: color_data = Z;
		19'b0101111100101101110: color_data = Z;
		19'b0101111100101101111: color_data = Z;
		19'b0101111100101110000: color_data = Z;
		19'b0101111100101110001: color_data = Z;
		19'b0101111100101110010: color_data = Z;
		19'b0101111100101110011: color_data = Z;
		19'b0101111100101110100: color_data = Z;
		19'b0101111100101111010: color_data = Z;
		19'b0101111100110000011: color_data = Z;
		19'b0101111100110000100: color_data = Z;
		19'b0101111100110000101: color_data = Z;
		19'b0101111100110000110: color_data = Z;
		19'b0101111100110000111: color_data = Z;
		19'b0101111100110001000: color_data = Z;
		19'b0101111100111010000: color_data = Z;
		19'b0101111100111010001: color_data = Z;
		19'b0101111100111010010: color_data = Z;
		19'b0101111100111010011: color_data = Z;
		19'b0101111100111010100: color_data = Z;
		19'b0101111100111010101: color_data = Z;
		19'b0101111100111010110: color_data = Z;
		19'b0101111100111010111: color_data = Z;
		19'b0101111100111011000: color_data = Z;
		19'b0101111100111011001: color_data = Z;
		19'b0101111100111011010: color_data = Z;
		19'b0101111100111011011: color_data = Z;
		19'b0101111110100011110: color_data = Z;
		19'b0101111110100011111: color_data = Z;
		19'b0101111110100100000: color_data = Z;
		19'b0101111110100100001: color_data = Z;
		19'b0101111110100100010: color_data = Z;
		19'b0101111110100100011: color_data = Z;
		19'b0101111110100100101: color_data = Z;
		19'b0101111110100100110: color_data = Z;
		19'b0101111110100100111: color_data = Z;
		19'b0101111110100101000: color_data = Z;
		19'b0101111110100101001: color_data = Z;
		19'b0101111110100101010: color_data = Z;
		19'b0101111110100101011: color_data = Z;
		19'b0101111110100101100: color_data = Z;
		19'b0101111110100101101: color_data = Z;
		19'b0101111110100101110: color_data = Z;
		19'b0101111110100101111: color_data = Z;
		19'b0101111110100110000: color_data = Z;
		19'b0101111110100110001: color_data = Z;
		19'b0101111110100110010: color_data = Z;
		19'b0101111110100110011: color_data = Z;
		19'b0101111110100110100: color_data = Z;
		19'b0101111110100110101: color_data = Z;
		19'b0101111110100110110: color_data = Z;
		19'b0101111110100110111: color_data = Z;
		19'b0101111110100111000: color_data = Z;
		19'b0101111110100111001: color_data = Z;
		19'b0101111110100111010: color_data = Z;
		19'b0101111110100111011: color_data = Z;
		19'b0101111110100111100: color_data = Z;
		19'b0101111110100111101: color_data = Z;
		19'b0101111110100111110: color_data = Z;
		19'b0101111110100111111: color_data = Z;
		19'b0101111110101000000: color_data = Z;
		19'b0101111110101000001: color_data = Z;
		19'b0101111110101000010: color_data = Z;
		19'b0101111110101000011: color_data = Z;
		19'b0101111110101000100: color_data = Z;
		19'b0101111110101000101: color_data = Z;
		19'b0101111110101000110: color_data = Z;
		19'b0101111110101000111: color_data = Z;
		19'b0101111110101001000: color_data = Z;
		19'b0101111110101001001: color_data = Z;
		19'b0101111110101001010: color_data = Z;
		19'b0101111110101001011: color_data = Z;
		19'b0101111110101001100: color_data = Z;
		19'b0101111110101001101: color_data = Z;
		19'b0101111110101001110: color_data = Z;
		19'b0101111110101001111: color_data = Z;
		19'b0101111110101010000: color_data = Z;
		19'b0101111110101010001: color_data = Z;
		19'b0101111110101010010: color_data = Z;
		19'b0101111110101010011: color_data = Z;
		19'b0101111110101010100: color_data = Z;
		19'b0101111110101010101: color_data = Z;
		19'b0101111110101010110: color_data = Z;
		19'b0101111110101010111: color_data = Z;
		19'b0101111110101011000: color_data = Z;
		19'b0101111110101011001: color_data = Z;
		19'b0101111110101011010: color_data = Z;
		19'b0101111110101011011: color_data = Z;
		19'b0101111110101011100: color_data = Z;
		19'b0101111110101011101: color_data = Z;
		19'b0101111110101011110: color_data = Z;
		19'b0101111110101011111: color_data = Z;
		19'b0101111110101100000: color_data = Z;
		19'b0101111110101100001: color_data = Z;
		19'b0101111110101100010: color_data = Z;
		19'b0101111110101100011: color_data = Z;
		19'b0101111110101100100: color_data = Z;
		19'b0101111110101100101: color_data = Z;
		19'b0101111110101100110: color_data = Z;
		19'b0101111110101100111: color_data = Z;
		19'b0101111110101101000: color_data = Z;
		19'b0101111110101101001: color_data = Z;
		19'b0101111110101101010: color_data = Z;
		19'b0101111110101101011: color_data = Z;
		19'b0101111110101101100: color_data = Z;
		19'b0101111110101101101: color_data = Z;
		19'b0101111110101101110: color_data = Z;
		19'b0101111110101101111: color_data = Z;
		19'b0101111110101110000: color_data = Z;
		19'b0101111110101110001: color_data = Z;
		19'b0101111110101110010: color_data = Z;
		19'b0101111110101110011: color_data = Z;
		19'b0101111110101110100: color_data = Z;
		19'b0101111110101111011: color_data = Z;
		19'b0101111110110000100: color_data = Z;
		19'b0101111110110000101: color_data = Z;
		19'b0101111110110000110: color_data = Z;
		19'b0101111110110000111: color_data = Z;
		19'b0101111110110001000: color_data = Z;
		19'b0101111110111010000: color_data = Z;
		19'b0101111110111010001: color_data = Z;
		19'b0101111110111010010: color_data = Z;
		19'b0101111110111010011: color_data = Z;
		19'b0101111110111010100: color_data = Z;
		19'b0101111110111010101: color_data = Z;
		19'b0101111110111010110: color_data = Z;
		19'b0101111110111010111: color_data = Z;
		19'b0101111110111011000: color_data = Z;
		19'b0101111110111011001: color_data = Z;
		19'b0101111110111011010: color_data = Z;
		19'b0101111110111011011: color_data = Z;
		19'b0110000000100011110: color_data = Z;
		19'b0110000000100011111: color_data = Z;
		19'b0110000000100100000: color_data = Z;
		19'b0110000000100100001: color_data = Z;
		19'b0110000000100100010: color_data = Z;
		19'b0110000000100100101: color_data = Z;
		19'b0110000000100100110: color_data = Z;
		19'b0110000000100100111: color_data = Z;
		19'b0110000000100101000: color_data = Z;
		19'b0110000000100101001: color_data = Z;
		19'b0110000000100101010: color_data = Z;
		19'b0110000000100101011: color_data = Z;
		19'b0110000000100101100: color_data = Z;
		19'b0110000000100101101: color_data = Z;
		19'b0110000000100101110: color_data = Z;
		19'b0110000000100101111: color_data = Z;
		19'b0110000000100110000: color_data = Z;
		19'b0110000000100110001: color_data = Z;
		19'b0110000000100110010: color_data = Z;
		19'b0110000000100110011: color_data = Z;
		19'b0110000000100110100: color_data = Z;
		19'b0110000000100110101: color_data = Z;
		19'b0110000000100110110: color_data = Z;
		19'b0110000000100110111: color_data = Z;
		19'b0110000000100111000: color_data = Z;
		19'b0110000000100111001: color_data = Z;
		19'b0110000000100111010: color_data = Z;
		19'b0110000000100111011: color_data = Z;
		19'b0110000000100111100: color_data = Z;
		19'b0110000000100111101: color_data = Z;
		19'b0110000000100111110: color_data = Z;
		19'b0110000000100111111: color_data = Z;
		19'b0110000000101000000: color_data = Z;
		19'b0110000000101000001: color_data = Z;
		19'b0110000000101000010: color_data = Z;
		19'b0110000000101000011: color_data = Z;
		19'b0110000000101000100: color_data = Z;
		19'b0110000000101000101: color_data = Z;
		19'b0110000000101000110: color_data = Z;
		19'b0110000000101000111: color_data = Z;
		19'b0110000000101001000: color_data = Z;
		19'b0110000000101001001: color_data = Z;
		19'b0110000000101001010: color_data = Z;
		19'b0110000000101001011: color_data = Z;
		19'b0110000000101001100: color_data = Z;
		19'b0110000000101001101: color_data = Z;
		19'b0110000000101001110: color_data = Z;
		19'b0110000000101001111: color_data = Z;
		19'b0110000000101010000: color_data = Z;
		19'b0110000000101010001: color_data = Z;
		19'b0110000000101010010: color_data = Z;
		19'b0110000000101010011: color_data = Z;
		19'b0110000000101010100: color_data = Z;
		19'b0110000000101010101: color_data = Z;
		19'b0110000000101010110: color_data = Z;
		19'b0110000000101010111: color_data = Z;
		19'b0110000000101011000: color_data = Z;
		19'b0110000000101011001: color_data = Z;
		19'b0110000000101011010: color_data = Z;
		19'b0110000000101011011: color_data = Z;
		19'b0110000000101011100: color_data = Z;
		19'b0110000000101011101: color_data = Z;
		19'b0110000000101011110: color_data = Z;
		19'b0110000000101011111: color_data = Z;
		19'b0110000000101100000: color_data = Z;
		19'b0110000000101100001: color_data = Z;
		19'b0110000000101100010: color_data = Z;
		19'b0110000000101100011: color_data = Z;
		19'b0110000000101100100: color_data = Z;
		19'b0110000000101100101: color_data = Z;
		19'b0110000000101100110: color_data = Z;
		19'b0110000000101100111: color_data = Z;
		19'b0110000000101101000: color_data = Z;
		19'b0110000000101101001: color_data = Z;
		19'b0110000000101101010: color_data = Z;
		19'b0110000000101101011: color_data = Z;
		19'b0110000000101101100: color_data = Z;
		19'b0110000000101101101: color_data = Z;
		19'b0110000000101101110: color_data = Z;
		19'b0110000000101101111: color_data = Z;
		19'b0110000000101110000: color_data = Z;
		19'b0110000000101110001: color_data = Z;
		19'b0110000000101110010: color_data = Z;
		19'b0110000000101110011: color_data = Z;
		19'b0110000000101110100: color_data = Z;
		19'b0110000000101110101: color_data = Z;
		19'b0110000000101111011: color_data = Z;
		19'b0110000000101111100: color_data = Z;
		19'b0110000000110000101: color_data = Z;
		19'b0110000000110000110: color_data = Z;
		19'b0110000000110000111: color_data = Z;
		19'b0110000000110001000: color_data = Z;
		19'b0110000000111010000: color_data = Z;
		19'b0110000000111010001: color_data = Z;
		19'b0110000000111010010: color_data = Z;
		19'b0110000000111010011: color_data = Z;
		19'b0110000000111010100: color_data = Z;
		19'b0110000000111010101: color_data = Z;
		19'b0110000000111010110: color_data = Z;
		19'b0110000000111010111: color_data = Z;
		19'b0110000000111011000: color_data = Z;
		19'b0110000000111011001: color_data = Z;
		19'b0110000000111011010: color_data = Z;
		19'b0110000000111011011: color_data = Z;
		19'b0110000010100011110: color_data = Z;
		19'b0110000010100011111: color_data = Z;
		19'b0110000010100100000: color_data = Z;
		19'b0110000010100100001: color_data = Z;
		19'b0110000010100100010: color_data = Z;
		19'b0110000010100100011: color_data = Z;
		19'b0110000010100100101: color_data = Z;
		19'b0110000010100100110: color_data = Z;
		19'b0110000010100100111: color_data = Z;
		19'b0110000010100101000: color_data = Z;
		19'b0110000010100101001: color_data = Z;
		19'b0110000010100101010: color_data = Z;
		19'b0110000010100101011: color_data = Z;
		19'b0110000010100101100: color_data = Z;
		19'b0110000010100101101: color_data = Z;
		19'b0110000010100101110: color_data = Z;
		19'b0110000010100101111: color_data = Z;
		19'b0110000010100110000: color_data = Z;
		19'b0110000010100110001: color_data = Z;
		19'b0110000010100110010: color_data = Z;
		19'b0110000010100110011: color_data = Z;
		19'b0110000010100110100: color_data = Z;
		19'b0110000010100110101: color_data = Z;
		19'b0110000010100110110: color_data = Z;
		19'b0110000010100110111: color_data = Z;
		19'b0110000010100111000: color_data = Z;
		19'b0110000010100111001: color_data = Z;
		19'b0110000010100111010: color_data = Z;
		19'b0110000010100111011: color_data = Z;
		19'b0110000010100111100: color_data = Z;
		19'b0110000010100111101: color_data = Z;
		19'b0110000010100111110: color_data = Z;
		19'b0110000010100111111: color_data = Z;
		19'b0110000010101000000: color_data = Z;
		19'b0110000010101000001: color_data = Z;
		19'b0110000010101000010: color_data = Z;
		19'b0110000010101000011: color_data = Z;
		19'b0110000010101000100: color_data = Z;
		19'b0110000010101000101: color_data = Z;
		19'b0110000010101000110: color_data = Z;
		19'b0110000010101000111: color_data = Z;
		19'b0110000010101001000: color_data = Z;
		19'b0110000010101001001: color_data = Z;
		19'b0110000010101001010: color_data = Z;
		19'b0110000010101001011: color_data = Z;
		19'b0110000010101001100: color_data = Z;
		19'b0110000010101001101: color_data = Z;
		19'b0110000010101001110: color_data = Z;
		19'b0110000010101001111: color_data = Z;
		19'b0110000010101010000: color_data = Z;
		19'b0110000010101010001: color_data = Z;
		19'b0110000010101010010: color_data = Z;
		19'b0110000010101010011: color_data = Z;
		19'b0110000010101010100: color_data = Z;
		19'b0110000010101010101: color_data = Z;
		19'b0110000010101010110: color_data = Z;
		19'b0110000010101010111: color_data = Z;
		19'b0110000010101011000: color_data = Z;
		19'b0110000010101011001: color_data = Z;
		19'b0110000010101011010: color_data = Z;
		19'b0110000010101011011: color_data = Z;
		19'b0110000010101011100: color_data = Z;
		19'b0110000010101011101: color_data = Z;
		19'b0110000010101011110: color_data = Z;
		19'b0110000010101011111: color_data = Z;
		19'b0110000010101100000: color_data = Z;
		19'b0110000010101100001: color_data = Z;
		19'b0110000010101100010: color_data = Z;
		19'b0110000010101100011: color_data = Z;
		19'b0110000010101100100: color_data = Z;
		19'b0110000010101100101: color_data = Z;
		19'b0110000010101100110: color_data = Z;
		19'b0110000010101100111: color_data = Z;
		19'b0110000010101101000: color_data = Z;
		19'b0110000010101101001: color_data = Z;
		19'b0110000010101101010: color_data = Z;
		19'b0110000010101101011: color_data = Z;
		19'b0110000010101101100: color_data = Z;
		19'b0110000010101101101: color_data = Z;
		19'b0110000010101101110: color_data = Z;
		19'b0110000010101101111: color_data = Z;
		19'b0110000010101110000: color_data = Z;
		19'b0110000010101110001: color_data = Z;
		19'b0110000010101110010: color_data = Z;
		19'b0110000010101110011: color_data = Z;
		19'b0110000010101110100: color_data = Z;
		19'b0110000010101110101: color_data = Z;
		19'b0110000010101111011: color_data = Z;
		19'b0110000010110000110: color_data = Z;
		19'b0110000010110000111: color_data = Z;
		19'b0110000010110001000: color_data = Z;
		19'b0110000010111010000: color_data = Z;
		19'b0110000010111010001: color_data = Z;
		19'b0110000010111010010: color_data = Z;
		19'b0110000010111010011: color_data = Z;
		19'b0110000010111010100: color_data = Z;
		19'b0110000010111010101: color_data = Z;
		19'b0110000010111010110: color_data = Z;
		19'b0110000010111010111: color_data = Z;
		19'b0110000010111011000: color_data = Z;
		19'b0110000010111011001: color_data = Z;
		19'b0110000010111011010: color_data = Z;
		19'b0110000010111011011: color_data = Z;
		19'b0110000100100011101: color_data = Z;
		19'b0110000100100011110: color_data = Z;
		19'b0110000100100011111: color_data = Z;
		19'b0110000100100100000: color_data = Z;
		19'b0110000100100100001: color_data = Z;
		19'b0110000100100100010: color_data = Z;
		19'b0110000100100100011: color_data = Z;
		19'b0110000100100100100: color_data = Z;
		19'b0110000100100100101: color_data = Z;
		19'b0110000100100100110: color_data = Z;
		19'b0110000100100100111: color_data = Z;
		19'b0110000100100101000: color_data = Z;
		19'b0110000100100101001: color_data = Z;
		19'b0110000100100101010: color_data = Z;
		19'b0110000100100101011: color_data = Z;
		19'b0110000100100101100: color_data = Z;
		19'b0110000100100101101: color_data = Z;
		19'b0110000100100101110: color_data = Z;
		19'b0110000100100101111: color_data = Z;
		19'b0110000100100110000: color_data = Z;
		19'b0110000100100110001: color_data = Z;
		19'b0110000100100110010: color_data = Z;
		19'b0110000100100110011: color_data = Z;
		19'b0110000100100110100: color_data = Z;
		19'b0110000100100110101: color_data = Z;
		19'b0110000100100110110: color_data = Z;
		19'b0110000100100110111: color_data = Z;
		19'b0110000100100111000: color_data = Z;
		19'b0110000100100111001: color_data = Z;
		19'b0110000100100111010: color_data = Z;
		19'b0110000100100111011: color_data = Z;
		19'b0110000100100111100: color_data = Z;
		19'b0110000100100111101: color_data = Z;
		19'b0110000100100111110: color_data = Z;
		19'b0110000100100111111: color_data = Z;
		19'b0110000100101000000: color_data = Z;
		19'b0110000100101000001: color_data = Z;
		19'b0110000100101000010: color_data = Z;
		19'b0110000100101000011: color_data = Z;
		19'b0110000100101000100: color_data = Z;
		19'b0110000100101000101: color_data = Z;
		19'b0110000100101000110: color_data = Z;
		19'b0110000100101000111: color_data = Z;
		19'b0110000100101001000: color_data = Z;
		19'b0110000100101001001: color_data = Z;
		19'b0110000100101001010: color_data = Z;
		19'b0110000100101001011: color_data = Z;
		19'b0110000100101001100: color_data = Z;
		19'b0110000100101001101: color_data = Z;
		19'b0110000100101001110: color_data = Z;
		19'b0110000100101001111: color_data = Z;
		19'b0110000100101010000: color_data = Z;
		19'b0110000100101010001: color_data = Z;
		19'b0110000100101010010: color_data = Z;
		19'b0110000100101010011: color_data = Z;
		19'b0110000100101010100: color_data = Z;
		19'b0110000100101010101: color_data = Z;
		19'b0110000100101010110: color_data = Z;
		19'b0110000100101010111: color_data = Z;
		19'b0110000100101011000: color_data = Z;
		19'b0110000100101011001: color_data = Z;
		19'b0110000100101011010: color_data = Z;
		19'b0110000100101011011: color_data = Z;
		19'b0110000100101011100: color_data = Z;
		19'b0110000100101011101: color_data = Z;
		19'b0110000100101011110: color_data = Z;
		19'b0110000100101011111: color_data = Z;
		19'b0110000100101100000: color_data = Z;
		19'b0110000100101100001: color_data = Z;
		19'b0110000100101100010: color_data = Z;
		19'b0110000100101100011: color_data = Z;
		19'b0110000100101100100: color_data = Z;
		19'b0110000100101100101: color_data = Z;
		19'b0110000100101100110: color_data = Z;
		19'b0110000100101100111: color_data = Z;
		19'b0110000100101101000: color_data = Z;
		19'b0110000100101101001: color_data = Z;
		19'b0110000100101101010: color_data = Z;
		19'b0110000100101101011: color_data = Z;
		19'b0110000100101101100: color_data = Z;
		19'b0110000100101101101: color_data = Z;
		19'b0110000100101101110: color_data = Z;
		19'b0110000100101101111: color_data = Z;
		19'b0110000100101110000: color_data = Z;
		19'b0110000100101110001: color_data = Z;
		19'b0110000100101110010: color_data = Z;
		19'b0110000100101110011: color_data = Z;
		19'b0110000100101110100: color_data = Z;
		19'b0110000100101110101: color_data = Z;
		19'b0110000100101111011: color_data = Z;
		19'b0110000100101111111: color_data = Z;
		19'b0110000100110000000: color_data = Z;
		19'b0110000100110000001: color_data = Z;
		19'b0110000100110001000: color_data = Z;
		19'b0110000100110001001: color_data = Z;
		19'b0110000100111010000: color_data = Z;
		19'b0110000100111010001: color_data = Z;
		19'b0110000100111010010: color_data = Z;
		19'b0110000100111010011: color_data = Z;
		19'b0110000100111010100: color_data = Z;
		19'b0110000100111010101: color_data = Z;
		19'b0110000100111010110: color_data = Z;
		19'b0110000100111010111: color_data = Z;
		19'b0110000100111011000: color_data = Z;
		19'b0110000100111011001: color_data = Z;
		19'b0110000100111011010: color_data = Z;
		19'b0110000100111011011: color_data = Z;
		19'b0110000100111011100: color_data = Z;
		19'b0110000110100011101: color_data = Z;
		19'b0110000110100011110: color_data = Z;
		19'b0110000110100011111: color_data = Z;
		19'b0110000110100100000: color_data = Z;
		19'b0110000110100100001: color_data = Z;
		19'b0110000110100100010: color_data = Z;
		19'b0110000110100100011: color_data = Z;
		19'b0110000110100100100: color_data = Z;
		19'b0110000110100100101: color_data = Z;
		19'b0110000110100100110: color_data = Z;
		19'b0110000110100100111: color_data = Z;
		19'b0110000110100101000: color_data = Z;
		19'b0110000110100101001: color_data = Z;
		19'b0110000110100101010: color_data = Z;
		19'b0110000110100101011: color_data = Z;
		19'b0110000110100101100: color_data = Z;
		19'b0110000110100101101: color_data = Z;
		19'b0110000110100101110: color_data = Z;
		19'b0110000110100101111: color_data = Z;
		19'b0110000110100110000: color_data = Z;
		19'b0110000110100110001: color_data = Z;
		19'b0110000110100110010: color_data = Z;
		19'b0110000110100110011: color_data = Z;
		19'b0110000110100110100: color_data = Z;
		19'b0110000110100110101: color_data = Z;
		19'b0110000110100110110: color_data = Z;
		19'b0110000110100110111: color_data = Z;
		19'b0110000110100111000: color_data = Z;
		19'b0110000110100111001: color_data = Z;
		19'b0110000110100111010: color_data = Z;
		19'b0110000110100111011: color_data = Z;
		19'b0110000110100111100: color_data = Z;
		19'b0110000110100111101: color_data = Z;
		19'b0110000110100111110: color_data = Z;
		19'b0110000110100111111: color_data = Z;
		19'b0110000110101000000: color_data = Z;
		19'b0110000110101000001: color_data = Z;
		19'b0110000110101000010: color_data = Z;
		19'b0110000110101000011: color_data = Z;
		19'b0110000110101000100: color_data = Z;
		19'b0110000110101000101: color_data = Z;
		19'b0110000110101000110: color_data = Z;
		19'b0110000110101000111: color_data = Z;
		19'b0110000110101001000: color_data = Z;
		19'b0110000110101001001: color_data = Z;
		19'b0110000110101001010: color_data = Z;
		19'b0110000110101001011: color_data = Z;
		19'b0110000110101001100: color_data = Z;
		19'b0110000110101001101: color_data = Z;
		19'b0110000110101001110: color_data = Z;
		19'b0110000110101001111: color_data = Z;
		19'b0110000110101010000: color_data = Z;
		19'b0110000110101010001: color_data = Z;
		19'b0110000110101010010: color_data = Z;
		19'b0110000110101010011: color_data = Z;
		19'b0110000110101010100: color_data = Z;
		19'b0110000110101010101: color_data = Z;
		19'b0110000110101010110: color_data = Z;
		19'b0110000110101010111: color_data = Z;
		19'b0110000110101011000: color_data = Z;
		19'b0110000110101011001: color_data = Z;
		19'b0110000110101011010: color_data = Z;
		19'b0110000110101011011: color_data = Z;
		19'b0110000110101011100: color_data = Z;
		19'b0110000110101011101: color_data = Z;
		19'b0110000110101011110: color_data = Z;
		19'b0110000110101011111: color_data = Z;
		19'b0110000110101100000: color_data = Z;
		19'b0110000110101100001: color_data = Z;
		19'b0110000110101100010: color_data = Z;
		19'b0110000110101100011: color_data = Z;
		19'b0110000110101100100: color_data = Z;
		19'b0110000110101100101: color_data = Z;
		19'b0110000110101100110: color_data = Z;
		19'b0110000110101100111: color_data = Z;
		19'b0110000110101101000: color_data = Z;
		19'b0110000110101101001: color_data = Z;
		19'b0110000110101101010: color_data = Z;
		19'b0110000110101101011: color_data = Z;
		19'b0110000110101101100: color_data = Z;
		19'b0110000110101101101: color_data = Z;
		19'b0110000110101101110: color_data = Z;
		19'b0110000110101101111: color_data = Z;
		19'b0110000110101110000: color_data = Z;
		19'b0110000110101110001: color_data = Z;
		19'b0110000110101110010: color_data = Z;
		19'b0110000110101110011: color_data = Z;
		19'b0110000110101110100: color_data = Z;
		19'b0110000110101110101: color_data = Z;
		19'b0110000110101111100: color_data = Z;
		19'b0110000110101111101: color_data = Z;
		19'b0110000110101111110: color_data = Z;
		19'b0110000110101111111: color_data = Z;
		19'b0110000110110000000: color_data = Z;
		19'b0110000110110000001: color_data = Z;
		19'b0110000110110000010: color_data = Z;
		19'b0110000110110001000: color_data = Z;
		19'b0110000110110001001: color_data = Z;
		19'b0110000110111010000: color_data = Z;
		19'b0110000110111010001: color_data = Z;
		19'b0110000110111010010: color_data = Z;
		19'b0110000110111010011: color_data = Z;
		19'b0110000110111010100: color_data = Z;
		19'b0110000110111010101: color_data = Z;
		19'b0110000110111010110: color_data = Z;
		19'b0110000110111010111: color_data = Z;
		19'b0110000110111011000: color_data = Z;
		19'b0110000110111011001: color_data = Z;
		19'b0110000110111011010: color_data = Z;
		19'b0110000110111011011: color_data = Z;
		19'b0110000110111011100: color_data = Z;
		19'b0110001000100011101: color_data = Z;
		19'b0110001000100011110: color_data = Z;
		19'b0110001000100011111: color_data = Z;
		19'b0110001000100100000: color_data = Z;
		19'b0110001000100100001: color_data = Z;
		19'b0110001000100100010: color_data = Z;
		19'b0110001000100100011: color_data = Z;
		19'b0110001000100100100: color_data = Z;
		19'b0110001000100100101: color_data = Z;
		19'b0110001000100100110: color_data = Z;
		19'b0110001000100100111: color_data = Z;
		19'b0110001000100101000: color_data = Z;
		19'b0110001000100101001: color_data = Z;
		19'b0110001000100101010: color_data = Z;
		19'b0110001000100101011: color_data = Z;
		19'b0110001000100101100: color_data = Z;
		19'b0110001000100101101: color_data = Z;
		19'b0110001000100101110: color_data = Z;
		19'b0110001000100101111: color_data = Z;
		19'b0110001000100110000: color_data = Z;
		19'b0110001000100110001: color_data = Z;
		19'b0110001000100110010: color_data = Z;
		19'b0110001000100110011: color_data = Z;
		19'b0110001000100110100: color_data = Z;
		19'b0110001000100110101: color_data = Z;
		19'b0110001000100110110: color_data = Z;
		19'b0110001000100110111: color_data = Z;
		19'b0110001000100111000: color_data = Z;
		19'b0110001000100111001: color_data = Z;
		19'b0110001000100111010: color_data = Z;
		19'b0110001000100111011: color_data = Z;
		19'b0110001000100111100: color_data = Z;
		19'b0110001000100111101: color_data = Z;
		19'b0110001000100111110: color_data = Z;
		19'b0110001000100111111: color_data = Z;
		19'b0110001000101000000: color_data = Z;
		19'b0110001000101000001: color_data = Z;
		19'b0110001000101000010: color_data = Z;
		19'b0110001000101000011: color_data = Z;
		19'b0110001000101000100: color_data = Z;
		19'b0110001000101000101: color_data = Z;
		19'b0110001000101000110: color_data = Z;
		19'b0110001000101000111: color_data = Z;
		19'b0110001000101001000: color_data = Z;
		19'b0110001000101001001: color_data = Z;
		19'b0110001000101001010: color_data = Z;
		19'b0110001000101001011: color_data = Z;
		19'b0110001000101001100: color_data = Z;
		19'b0110001000101001101: color_data = Z;
		19'b0110001000101001110: color_data = Z;
		19'b0110001000101001111: color_data = Z;
		19'b0110001000101010000: color_data = Z;
		19'b0110001000101010001: color_data = Z;
		19'b0110001000101010010: color_data = Z;
		19'b0110001000101010011: color_data = Z;
		19'b0110001000101010100: color_data = Z;
		19'b0110001000101010101: color_data = Z;
		19'b0110001000101010110: color_data = Z;
		19'b0110001000101010111: color_data = Z;
		19'b0110001000101011000: color_data = Z;
		19'b0110001000101011001: color_data = Z;
		19'b0110001000101011010: color_data = Z;
		19'b0110001000101011011: color_data = Z;
		19'b0110001000101011100: color_data = Z;
		19'b0110001000101011101: color_data = Z;
		19'b0110001000101011110: color_data = Z;
		19'b0110001000101011111: color_data = Z;
		19'b0110001000101100000: color_data = Z;
		19'b0110001000101100001: color_data = Z;
		19'b0110001000101100010: color_data = Z;
		19'b0110001000101100011: color_data = Z;
		19'b0110001000101100100: color_data = Z;
		19'b0110001000101100101: color_data = Z;
		19'b0110001000101100110: color_data = Z;
		19'b0110001000101100111: color_data = Z;
		19'b0110001000101101000: color_data = Z;
		19'b0110001000101101001: color_data = Z;
		19'b0110001000101101010: color_data = Z;
		19'b0110001000101101011: color_data = Z;
		19'b0110001000101101100: color_data = Z;
		19'b0110001000101101101: color_data = Z;
		19'b0110001000101101110: color_data = Z;
		19'b0110001000101101111: color_data = Z;
		19'b0110001000101110000: color_data = Z;
		19'b0110001000101110001: color_data = Z;
		19'b0110001000101110010: color_data = Z;
		19'b0110001000101110011: color_data = Z;
		19'b0110001000101110100: color_data = Z;
		19'b0110001000101110101: color_data = Z;
		19'b0110001000101111100: color_data = Z;
		19'b0110001000101111101: color_data = Z;
		19'b0110001000101111110: color_data = Z;
		19'b0110001000101111111: color_data = Z;
		19'b0110001000110000000: color_data = Z;
		19'b0110001000110000001: color_data = Z;
		19'b0110001000110000010: color_data = Z;
		19'b0110001000110000011: color_data = Z;
		19'b0110001000110001001: color_data = Z;
		19'b0110001000110001010: color_data = Z;
		19'b0110001000111010000: color_data = Z;
		19'b0110001000111010001: color_data = Z;
		19'b0110001000111010010: color_data = Z;
		19'b0110001000111010011: color_data = Z;
		19'b0110001000111010100: color_data = Z;
		19'b0110001000111010101: color_data = Z;
		19'b0110001000111010110: color_data = Z;
		19'b0110001000111010111: color_data = Z;
		19'b0110001000111011000: color_data = Z;
		19'b0110001000111011001: color_data = Z;
		19'b0110001000111011010: color_data = Z;
		19'b0110001000111011011: color_data = Z;
		19'b0110001010010100000: color_data = Z;
		19'b0110001010100011100: color_data = Z;
		19'b0110001010100011101: color_data = Z;
		19'b0110001010100011110: color_data = Z;
		19'b0110001010100011111: color_data = Z;
		19'b0110001010100100000: color_data = Z;
		19'b0110001010100100010: color_data = Z;
		19'b0110001010100100011: color_data = Z;
		19'b0110001010100100100: color_data = Z;
		19'b0110001010100100101: color_data = Z;
		19'b0110001010100100110: color_data = Z;
		19'b0110001010100100111: color_data = Z;
		19'b0110001010100101000: color_data = Z;
		19'b0110001010100101001: color_data = Z;
		19'b0110001010100101010: color_data = Z;
		19'b0110001010100101011: color_data = Z;
		19'b0110001010100101100: color_data = Z;
		19'b0110001010100101101: color_data = Z;
		19'b0110001010100101110: color_data = Z;
		19'b0110001010100101111: color_data = Z;
		19'b0110001010100110000: color_data = Z;
		19'b0110001010100110001: color_data = Z;
		19'b0110001010100110010: color_data = Z;
		19'b0110001010100110011: color_data = Z;
		19'b0110001010100110100: color_data = Z;
		19'b0110001010100110101: color_data = Z;
		19'b0110001010100110110: color_data = Z;
		19'b0110001010100110111: color_data = Z;
		19'b0110001010100111000: color_data = Z;
		19'b0110001010100111001: color_data = Z;
		19'b0110001010100111010: color_data = Z;
		19'b0110001010100111011: color_data = Z;
		19'b0110001010100111100: color_data = Z;
		19'b0110001010100111101: color_data = Z;
		19'b0110001010100111110: color_data = Z;
		19'b0110001010100111111: color_data = Z;
		19'b0110001010101000000: color_data = Z;
		19'b0110001010101000001: color_data = Z;
		19'b0110001010101000010: color_data = Z;
		19'b0110001010101000011: color_data = Z;
		19'b0110001010101000100: color_data = Z;
		19'b0110001010101000101: color_data = Z;
		19'b0110001010101000110: color_data = Z;
		19'b0110001010101000111: color_data = Z;
		19'b0110001010101001000: color_data = Z;
		19'b0110001010101001001: color_data = Z;
		19'b0110001010101001010: color_data = Z;
		19'b0110001010101001011: color_data = Z;
		19'b0110001010101001100: color_data = Z;
		19'b0110001010101001101: color_data = Z;
		19'b0110001010101001110: color_data = Z;
		19'b0110001010101001111: color_data = Z;
		19'b0110001010101010000: color_data = Z;
		19'b0110001010101010001: color_data = Z;
		19'b0110001010101010010: color_data = Z;
		19'b0110001010101010011: color_data = Z;
		19'b0110001010101010100: color_data = Z;
		19'b0110001010101010101: color_data = Z;
		19'b0110001010101010110: color_data = Z;
		19'b0110001010101010111: color_data = Z;
		19'b0110001010101011000: color_data = Z;
		19'b0110001010101011001: color_data = Z;
		19'b0110001010101011010: color_data = Z;
		19'b0110001010101011011: color_data = Z;
		19'b0110001010101011100: color_data = Z;
		19'b0110001010101011101: color_data = Z;
		19'b0110001010101011110: color_data = Z;
		19'b0110001010101011111: color_data = Z;
		19'b0110001010101100000: color_data = Z;
		19'b0110001010101100001: color_data = Z;
		19'b0110001010101100010: color_data = Z;
		19'b0110001010101100011: color_data = Z;
		19'b0110001010101100100: color_data = Z;
		19'b0110001010101100101: color_data = Z;
		19'b0110001010101100110: color_data = Z;
		19'b0110001010101100111: color_data = Z;
		19'b0110001010101101000: color_data = Z;
		19'b0110001010101101001: color_data = Z;
		19'b0110001010101101010: color_data = Z;
		19'b0110001010101101011: color_data = Z;
		19'b0110001010101101100: color_data = Z;
		19'b0110001010101101101: color_data = Z;
		19'b0110001010101101110: color_data = Z;
		19'b0110001010101101111: color_data = Z;
		19'b0110001010101110000: color_data = Z;
		19'b0110001010101110001: color_data = Z;
		19'b0110001010101110010: color_data = Z;
		19'b0110001010101110011: color_data = Z;
		19'b0110001010101110100: color_data = Z;
		19'b0110001010101110101: color_data = Z;
		19'b0110001010101110110: color_data = Z;
		19'b0110001010101111100: color_data = Z;
		19'b0110001010101111101: color_data = Z;
		19'b0110001010101111110: color_data = Z;
		19'b0110001010101111111: color_data = Z;
		19'b0110001010110000000: color_data = Z;
		19'b0110001010110000001: color_data = Z;
		19'b0110001010110000010: color_data = Z;
		19'b0110001010110000011: color_data = Z;
		19'b0110001010110001010: color_data = Z;
		19'b0110001010110001011: color_data = Z;
		19'b0110001010111010000: color_data = Z;
		19'b0110001010111010001: color_data = Z;
		19'b0110001010111010010: color_data = Z;
		19'b0110001010111010011: color_data = Z;
		19'b0110001010111010100: color_data = Z;
		19'b0110001010111010101: color_data = Z;
		19'b0110001010111010110: color_data = Z;
		19'b0110001010111010111: color_data = Z;
		19'b0110001010111011000: color_data = Z;
		19'b0110001010111011001: color_data = Z;
		19'b0110001010111011010: color_data = Z;
		19'b0110001010111011011: color_data = Z;
		19'b0110001100010100000: color_data = Z;
		19'b0110001100100011100: color_data = Z;
		19'b0110001100100011101: color_data = Z;
		19'b0110001100100011110: color_data = Z;
		19'b0110001100100011111: color_data = Z;
		19'b0110001100100100010: color_data = Z;
		19'b0110001100100100011: color_data = Z;
		19'b0110001100100100100: color_data = Z;
		19'b0110001100100100101: color_data = Z;
		19'b0110001100100100110: color_data = Z;
		19'b0110001100100100111: color_data = Z;
		19'b0110001100100101000: color_data = Z;
		19'b0110001100100101001: color_data = Z;
		19'b0110001100100101010: color_data = Z;
		19'b0110001100100101100: color_data = Z;
		19'b0110001100100101101: color_data = Z;
		19'b0110001100100101110: color_data = Z;
		19'b0110001100100101111: color_data = Z;
		19'b0110001100100110000: color_data = Z;
		19'b0110001100100110001: color_data = Z;
		19'b0110001100100110010: color_data = Z;
		19'b0110001100100110011: color_data = Z;
		19'b0110001100100110100: color_data = Z;
		19'b0110001100100110101: color_data = Z;
		19'b0110001100100110110: color_data = Z;
		19'b0110001100100110111: color_data = Z;
		19'b0110001100100111000: color_data = Z;
		19'b0110001100100111001: color_data = Z;
		19'b0110001100100111010: color_data = Z;
		19'b0110001100100111011: color_data = Z;
		19'b0110001100100111100: color_data = Z;
		19'b0110001100100111101: color_data = Z;
		19'b0110001100100111110: color_data = Z;
		19'b0110001100100111111: color_data = Z;
		19'b0110001100101000000: color_data = Z;
		19'b0110001100101000001: color_data = Z;
		19'b0110001100101000010: color_data = Z;
		19'b0110001100101000011: color_data = Z;
		19'b0110001100101000100: color_data = Z;
		19'b0110001100101000101: color_data = Z;
		19'b0110001100101000110: color_data = Z;
		19'b0110001100101000111: color_data = Z;
		19'b0110001100101001000: color_data = Z;
		19'b0110001100101001001: color_data = Z;
		19'b0110001100101001010: color_data = Z;
		19'b0110001100101001011: color_data = Z;
		19'b0110001100101001100: color_data = Z;
		19'b0110001100101001101: color_data = Z;
		19'b0110001100101001110: color_data = Z;
		19'b0110001100101001111: color_data = Z;
		19'b0110001100101010000: color_data = Z;
		19'b0110001100101010001: color_data = Z;
		19'b0110001100101010010: color_data = Z;
		19'b0110001100101010011: color_data = Z;
		19'b0110001100101010100: color_data = Z;
		19'b0110001100101010101: color_data = Z;
		19'b0110001100101010110: color_data = Z;
		19'b0110001100101010111: color_data = Z;
		19'b0110001100101011000: color_data = Z;
		19'b0110001100101011001: color_data = Z;
		19'b0110001100101011010: color_data = Z;
		19'b0110001100101011011: color_data = Z;
		19'b0110001100101011100: color_data = Z;
		19'b0110001100101011101: color_data = Z;
		19'b0110001100101011110: color_data = Z;
		19'b0110001100101011111: color_data = Z;
		19'b0110001100101100000: color_data = Z;
		19'b0110001100101100001: color_data = Z;
		19'b0110001100101100010: color_data = Z;
		19'b0110001100101100011: color_data = Z;
		19'b0110001100101100100: color_data = Z;
		19'b0110001100101100101: color_data = Z;
		19'b0110001100101100110: color_data = Z;
		19'b0110001100101100111: color_data = Z;
		19'b0110001100101101000: color_data = Z;
		19'b0110001100101101001: color_data = Z;
		19'b0110001100101101010: color_data = Z;
		19'b0110001100101101011: color_data = Z;
		19'b0110001100101101100: color_data = Z;
		19'b0110001100101101101: color_data = Z;
		19'b0110001100101101110: color_data = Z;
		19'b0110001100101101111: color_data = Z;
		19'b0110001100101110000: color_data = Z;
		19'b0110001100101110001: color_data = Z;
		19'b0110001100101110010: color_data = Z;
		19'b0110001100101110011: color_data = Z;
		19'b0110001100101110100: color_data = Z;
		19'b0110001100101110101: color_data = Z;
		19'b0110001100101110110: color_data = Z;
		19'b0110001100101111101: color_data = Z;
		19'b0110001100101111110: color_data = Z;
		19'b0110001100101111111: color_data = Z;
		19'b0110001100110000000: color_data = Z;
		19'b0110001100110000001: color_data = Z;
		19'b0110001100110000010: color_data = Z;
		19'b0110001100110000011: color_data = Z;
		19'b0110001100110000100: color_data = Z;
		19'b0110001100110001010: color_data = Z;
		19'b0110001100110001011: color_data = Z;
		19'b0110001100110001100: color_data = Z;
		19'b0110001100111010000: color_data = Z;
		19'b0110001100111010001: color_data = Z;
		19'b0110001100111010010: color_data = Z;
		19'b0110001100111010011: color_data = Z;
		19'b0110001100111010100: color_data = Z;
		19'b0110001100111010101: color_data = Z;
		19'b0110001100111010110: color_data = Z;
		19'b0110001100111010111: color_data = Z;
		19'b0110001100111011000: color_data = Z;
		19'b0110001100111011001: color_data = Z;
		19'b0110001100111011010: color_data = Z;
		19'b0110001100111011011: color_data = Z;
		19'b0110001110010100000: color_data = Z;
		19'b0110001110100011100: color_data = Z;
		19'b0110001110100011101: color_data = Z;
		19'b0110001110100011110: color_data = Z;
		19'b0110001110100011111: color_data = Z;
		19'b0110001110100100001: color_data = Z;
		19'b0110001110100100010: color_data = Z;
		19'b0110001110100100011: color_data = Z;
		19'b0110001110100100100: color_data = Z;
		19'b0110001110100100101: color_data = Z;
		19'b0110001110100100110: color_data = Z;
		19'b0110001110100100111: color_data = Z;
		19'b0110001110100101000: color_data = Z;
		19'b0110001110100101001: color_data = Z;
		19'b0110001110100101010: color_data = Z;
		19'b0110001110100101101: color_data = Z;
		19'b0110001110100101110: color_data = Z;
		19'b0110001110100101111: color_data = Z;
		19'b0110001110100110000: color_data = Z;
		19'b0110001110100110001: color_data = Z;
		19'b0110001110100110010: color_data = Z;
		19'b0110001110100110011: color_data = Z;
		19'b0110001110100110100: color_data = Z;
		19'b0110001110100110101: color_data = Z;
		19'b0110001110100110110: color_data = Z;
		19'b0110001110100110111: color_data = Z;
		19'b0110001110100111000: color_data = Z;
		19'b0110001110100111001: color_data = Z;
		19'b0110001110100111010: color_data = Z;
		19'b0110001110100111011: color_data = Z;
		19'b0110001110100111100: color_data = Z;
		19'b0110001110100111101: color_data = Z;
		19'b0110001110100111110: color_data = Z;
		19'b0110001110100111111: color_data = Z;
		19'b0110001110101000000: color_data = Z;
		19'b0110001110101000001: color_data = Z;
		19'b0110001110101000010: color_data = Z;
		19'b0110001110101000011: color_data = Z;
		19'b0110001110101000100: color_data = Z;
		19'b0110001110101000101: color_data = Z;
		19'b0110001110101000110: color_data = Z;
		19'b0110001110101000111: color_data = Z;
		19'b0110001110101001000: color_data = Z;
		19'b0110001110101001001: color_data = Z;
		19'b0110001110101001010: color_data = Z;
		19'b0110001110101001011: color_data = Z;
		19'b0110001110101001100: color_data = Z;
		19'b0110001110101001101: color_data = Z;
		19'b0110001110101001110: color_data = Z;
		19'b0110001110101001111: color_data = Z;
		19'b0110001110101010000: color_data = Z;
		19'b0110001110101010001: color_data = Z;
		19'b0110001110101010010: color_data = Z;
		19'b0110001110101010011: color_data = Z;
		19'b0110001110101010100: color_data = Z;
		19'b0110001110101010101: color_data = Z;
		19'b0110001110101010110: color_data = Z;
		19'b0110001110101010111: color_data = Z;
		19'b0110001110101011000: color_data = Z;
		19'b0110001110101011001: color_data = Z;
		19'b0110001110101011010: color_data = Z;
		19'b0110001110101011011: color_data = Z;
		19'b0110001110101011100: color_data = Z;
		19'b0110001110101011101: color_data = Z;
		19'b0110001110101011110: color_data = Z;
		19'b0110001110101011111: color_data = Z;
		19'b0110001110101100000: color_data = Z;
		19'b0110001110101100001: color_data = Z;
		19'b0110001110101100010: color_data = Z;
		19'b0110001110101100011: color_data = Z;
		19'b0110001110101100100: color_data = Z;
		19'b0110001110101100101: color_data = Z;
		19'b0110001110101100110: color_data = Z;
		19'b0110001110101100111: color_data = Z;
		19'b0110001110101101000: color_data = Z;
		19'b0110001110101101001: color_data = Z;
		19'b0110001110101101010: color_data = Z;
		19'b0110001110101101011: color_data = Z;
		19'b0110001110101101100: color_data = Z;
		19'b0110001110101101101: color_data = Z;
		19'b0110001110101101110: color_data = Z;
		19'b0110001110101101111: color_data = Z;
		19'b0110001110101110000: color_data = Z;
		19'b0110001110101110001: color_data = Z;
		19'b0110001110101110010: color_data = Z;
		19'b0110001110101110011: color_data = Z;
		19'b0110001110101110100: color_data = Z;
		19'b0110001110101110101: color_data = Z;
		19'b0110001110101110110: color_data = Z;
		19'b0110001110101111101: color_data = Z;
		19'b0110001110101111110: color_data = Z;
		19'b0110001110101111111: color_data = Z;
		19'b0110001110110000000: color_data = Z;
		19'b0110001110110000001: color_data = Z;
		19'b0110001110110000010: color_data = Z;
		19'b0110001110110000011: color_data = Z;
		19'b0110001110110000100: color_data = Z;
		19'b0110001110110001011: color_data = Z;
		19'b0110001110110001100: color_data = Z;
		19'b0110001110110001101: color_data = Z;
		19'b0110001110110001110: color_data = Z;
		19'b0110001110110001111: color_data = Z;
		19'b0110001110110010000: color_data = Z;
		19'b0110001110111010001: color_data = Z;
		19'b0110001110111010010: color_data = Z;
		19'b0110001110111010011: color_data = Z;
		19'b0110001110111010100: color_data = Z;
		19'b0110001110111010101: color_data = Z;
		19'b0110001110111010110: color_data = Z;
		19'b0110001110111010111: color_data = Z;
		19'b0110001110111011000: color_data = Z;
		19'b0110001110111011001: color_data = Z;
		19'b0110001110111011010: color_data = Z;
		19'b0110001110111011011: color_data = Z;
		19'b0110010000010100000: color_data = Z;
		19'b0110010000100011011: color_data = Z;
		19'b0110010000100011100: color_data = Z;
		19'b0110010000100011101: color_data = Z;
		19'b0110010000100011110: color_data = Z;
		19'b0110010000100011111: color_data = Z;
		19'b0110010000100100000: color_data = Z;
		19'b0110010000100100001: color_data = Z;
		19'b0110010000100100010: color_data = Z;
		19'b0110010000100100011: color_data = Z;
		19'b0110010000100100100: color_data = Z;
		19'b0110010000100100101: color_data = Z;
		19'b0110010000100100110: color_data = Z;
		19'b0110010000100100111: color_data = Z;
		19'b0110010000100101000: color_data = Z;
		19'b0110010000100101001: color_data = Z;
		19'b0110010000100101010: color_data = Z;
		19'b0110010000100101100: color_data = Z;
		19'b0110010000100101101: color_data = Z;
		19'b0110010000100101110: color_data = Z;
		19'b0110010000100101111: color_data = Z;
		19'b0110010000100110000: color_data = Z;
		19'b0110010000100110001: color_data = Z;
		19'b0110010000100110010: color_data = Z;
		19'b0110010000100110011: color_data = Z;
		19'b0110010000100110100: color_data = Z;
		19'b0110010000100110101: color_data = Z;
		19'b0110010000100110110: color_data = Z;
		19'b0110010000100110111: color_data = Z;
		19'b0110010000100111000: color_data = Z;
		19'b0110010000100111001: color_data = Z;
		19'b0110010000100111010: color_data = Z;
		19'b0110010000100111011: color_data = Z;
		19'b0110010000100111100: color_data = Z;
		19'b0110010000100111101: color_data = Z;
		19'b0110010000100111110: color_data = Z;
		19'b0110010000100111111: color_data = Z;
		19'b0110010000101000000: color_data = Z;
		19'b0110010000101000001: color_data = Z;
		19'b0110010000101000010: color_data = Z;
		19'b0110010000101000011: color_data = Z;
		19'b0110010000101000100: color_data = Z;
		19'b0110010000101000101: color_data = Z;
		19'b0110010000101000110: color_data = Z;
		19'b0110010000101000111: color_data = Z;
		19'b0110010000101001000: color_data = Z;
		19'b0110010000101001001: color_data = Z;
		19'b0110010000101001010: color_data = Z;
		19'b0110010000101001011: color_data = Z;
		19'b0110010000101001100: color_data = Z;
		19'b0110010000101001101: color_data = Z;
		19'b0110010000101001110: color_data = Z;
		19'b0110010000101001111: color_data = Z;
		19'b0110010000101010000: color_data = Z;
		19'b0110010000101010001: color_data = Z;
		19'b0110010000101010010: color_data = Z;
		19'b0110010000101010011: color_data = Z;
		19'b0110010000101010100: color_data = Z;
		19'b0110010000101010101: color_data = Z;
		19'b0110010000101010110: color_data = Z;
		19'b0110010000101010111: color_data = Z;
		19'b0110010000101011000: color_data = Z;
		19'b0110010000101011001: color_data = Z;
		19'b0110010000101011010: color_data = Z;
		19'b0110010000101011011: color_data = Z;
		19'b0110010000101011100: color_data = Z;
		19'b0110010000101011101: color_data = Z;
		19'b0110010000101011110: color_data = Z;
		19'b0110010000101011111: color_data = Z;
		19'b0110010000101100000: color_data = Z;
		19'b0110010000101100001: color_data = Z;
		19'b0110010000101100010: color_data = Z;
		19'b0110010000101100011: color_data = Z;
		19'b0110010000101100100: color_data = Z;
		19'b0110010000101100101: color_data = Z;
		19'b0110010000101100110: color_data = Z;
		19'b0110010000101100111: color_data = Z;
		19'b0110010000101101000: color_data = Z;
		19'b0110010000101101001: color_data = Z;
		19'b0110010000101101010: color_data = Z;
		19'b0110010000101101011: color_data = Z;
		19'b0110010000101101100: color_data = Z;
		19'b0110010000101101101: color_data = Z;
		19'b0110010000101101110: color_data = Z;
		19'b0110010000101101111: color_data = Z;
		19'b0110010000101110000: color_data = Z;
		19'b0110010000101110001: color_data = Z;
		19'b0110010000101110010: color_data = Z;
		19'b0110010000101110011: color_data = Z;
		19'b0110010000101110100: color_data = Z;
		19'b0110010000101110101: color_data = Z;
		19'b0110010000101110110: color_data = Z;
		19'b0110010000101111101: color_data = Z;
		19'b0110010000101111110: color_data = Z;
		19'b0110010000101111111: color_data = Z;
		19'b0110010000110000000: color_data = Z;
		19'b0110010000110000001: color_data = Z;
		19'b0110010000110000010: color_data = Z;
		19'b0110010000110000011: color_data = Z;
		19'b0110010000110000100: color_data = Z;
		19'b0110010000110000101: color_data = Z;
		19'b0110010000110001100: color_data = Z;
		19'b0110010000110001101: color_data = Z;
		19'b0110010000110001110: color_data = Z;
		19'b0110010000110001111: color_data = Z;
		19'b0110010000110010000: color_data = Z;
		19'b0110010000110010001: color_data = Z;
		19'b0110010000111010001: color_data = Z;
		19'b0110010000111010010: color_data = Z;
		19'b0110010000111010011: color_data = Z;
		19'b0110010000111010100: color_data = Z;
		19'b0110010000111010101: color_data = Z;
		19'b0110010000111010110: color_data = Z;
		19'b0110010000111010111: color_data = Z;
		19'b0110010000111011000: color_data = Z;
		19'b0110010000111011001: color_data = Z;
		19'b0110010000111011010: color_data = Z;
		19'b0110010000111011011: color_data = Z;
		19'b0110010010010100000: color_data = Z;
		19'b0110010010100011010: color_data = Z;
		19'b0110010010100011011: color_data = Z;
		19'b0110010010100011100: color_data = Z;
		19'b0110010010100011101: color_data = Z;
		19'b0110010010100011110: color_data = Z;
		19'b0110010010100011111: color_data = Z;
		19'b0110010010100100000: color_data = Z;
		19'b0110010010100100001: color_data = Z;
		19'b0110010010100100010: color_data = Z;
		19'b0110010010100100011: color_data = Z;
		19'b0110010010100100100: color_data = Z;
		19'b0110010010100100101: color_data = Z;
		19'b0110010010100100110: color_data = Z;
		19'b0110010010100100111: color_data = Z;
		19'b0110010010100101000: color_data = Z;
		19'b0110010010100101001: color_data = Z;
		19'b0110010010100101010: color_data = Z;
		19'b0110010010100101011: color_data = Z;
		19'b0110010010100101100: color_data = Z;
		19'b0110010010100101101: color_data = Z;
		19'b0110010010100101110: color_data = Z;
		19'b0110010010100101111: color_data = Z;
		19'b0110010010100110000: color_data = Z;
		19'b0110010010100110001: color_data = Z;
		19'b0110010010100110010: color_data = Z;
		19'b0110010010100110011: color_data = Z;
		19'b0110010010100110100: color_data = Z;
		19'b0110010010100110101: color_data = Z;
		19'b0110010010100110110: color_data = Z;
		19'b0110010010100110111: color_data = Z;
		19'b0110010010100111000: color_data = Z;
		19'b0110010010100111001: color_data = Z;
		19'b0110010010100111010: color_data = Z;
		19'b0110010010100111011: color_data = Z;
		19'b0110010010100111100: color_data = Z;
		19'b0110010010100111101: color_data = Z;
		19'b0110010010100111110: color_data = Z;
		19'b0110010010100111111: color_data = Z;
		19'b0110010010101000000: color_data = Z;
		19'b0110010010101000001: color_data = Z;
		19'b0110010010101000010: color_data = Z;
		19'b0110010010101000011: color_data = Z;
		19'b0110010010101000100: color_data = Z;
		19'b0110010010101000101: color_data = Z;
		19'b0110010010101000110: color_data = Z;
		19'b0110010010101000111: color_data = Z;
		19'b0110010010101001000: color_data = Z;
		19'b0110010010101001001: color_data = Z;
		19'b0110010010101001010: color_data = Z;
		19'b0110010010101001011: color_data = Z;
		19'b0110010010101001100: color_data = Z;
		19'b0110010010101001101: color_data = Z;
		19'b0110010010101001110: color_data = Z;
		19'b0110010010101001111: color_data = Z;
		19'b0110010010101010000: color_data = Z;
		19'b0110010010101010001: color_data = Z;
		19'b0110010010101010010: color_data = Z;
		19'b0110010010101010011: color_data = Z;
		19'b0110010010101010100: color_data = Z;
		19'b0110010010101010101: color_data = Z;
		19'b0110010010101010110: color_data = Z;
		19'b0110010010101010111: color_data = Z;
		19'b0110010010101011000: color_data = Z;
		19'b0110010010101011001: color_data = Z;
		19'b0110010010101011010: color_data = Z;
		19'b0110010010101011011: color_data = Z;
		19'b0110010010101011100: color_data = Z;
		19'b0110010010101011101: color_data = Z;
		19'b0110010010101011110: color_data = Z;
		19'b0110010010101011111: color_data = Z;
		19'b0110010010101100000: color_data = Z;
		19'b0110010010101100001: color_data = Z;
		19'b0110010010101100010: color_data = Z;
		19'b0110010010101100011: color_data = Z;
		19'b0110010010101100100: color_data = Z;
		19'b0110010010101100101: color_data = Z;
		19'b0110010010101100110: color_data = Z;
		19'b0110010010101100111: color_data = Z;
		19'b0110010010101101000: color_data = Z;
		19'b0110010010101101001: color_data = Z;
		19'b0110010010101101010: color_data = Z;
		19'b0110010010101101011: color_data = Z;
		19'b0110010010101101100: color_data = Z;
		19'b0110010010101101101: color_data = Z;
		19'b0110010010101101110: color_data = Z;
		19'b0110010010101101111: color_data = Z;
		19'b0110010010101110000: color_data = Z;
		19'b0110010010101110001: color_data = Z;
		19'b0110010010101110010: color_data = Z;
		19'b0110010010101110011: color_data = Z;
		19'b0110010010101110100: color_data = Z;
		19'b0110010010101110101: color_data = Z;
		19'b0110010010101110110: color_data = Z;
		19'b0110010010101110111: color_data = Z;
		19'b0110010010101111101: color_data = Z;
		19'b0110010010101111110: color_data = Z;
		19'b0110010010101111111: color_data = Z;
		19'b0110010010110000000: color_data = Z;
		19'b0110010010110000001: color_data = Z;
		19'b0110010010110000010: color_data = Z;
		19'b0110010010110000011: color_data = Z;
		19'b0110010010110000100: color_data = Z;
		19'b0110010010110000101: color_data = Z;
		19'b0110010010110000110: color_data = Z;
		19'b0110010010110001100: color_data = Z;
		19'b0110010010110001101: color_data = Z;
		19'b0110010010110001110: color_data = Z;
		19'b0110010010110001111: color_data = Z;
		19'b0110010010110010000: color_data = Z;
		19'b0110010010110010001: color_data = Z;
		19'b0110010010110010010: color_data = Z;
		19'b0110010010111010001: color_data = Z;
		19'b0110010010111010010: color_data = Z;
		19'b0110010010111010011: color_data = Z;
		19'b0110010010111010100: color_data = Z;
		19'b0110010010111010101: color_data = Z;
		19'b0110010010111010110: color_data = Z;
		19'b0110010010111010111: color_data = Z;
		19'b0110010010111011000: color_data = Z;
		19'b0110010010111011001: color_data = Z;
		19'b0110010010111011010: color_data = Z;
		19'b0110010010111011011: color_data = Z;
		19'b0110010100010100000: color_data = Z;
		19'b0110010100010100001: color_data = Z;
		19'b0110010100100011000: color_data = Z;
		19'b0110010100100011001: color_data = Z;
		19'b0110010100100011010: color_data = Z;
		19'b0110010100100011011: color_data = Z;
		19'b0110010100100011100: color_data = Z;
		19'b0110010100100011101: color_data = Z;
		19'b0110010100100011110: color_data = Z;
		19'b0110010100100011111: color_data = Z;
		19'b0110010100100100000: color_data = Z;
		19'b0110010100100100001: color_data = Z;
		19'b0110010100100100010: color_data = Z;
		19'b0110010100100100011: color_data = Z;
		19'b0110010100100100100: color_data = Z;
		19'b0110010100100100101: color_data = Z;
		19'b0110010100100100110: color_data = Z;
		19'b0110010100100100111: color_data = Z;
		19'b0110010100100101000: color_data = Z;
		19'b0110010100100101001: color_data = Z;
		19'b0110010100100101010: color_data = Z;
		19'b0110010100100101011: color_data = Z;
		19'b0110010100100101100: color_data = Z;
		19'b0110010100100101101: color_data = Z;
		19'b0110010100100101110: color_data = Z;
		19'b0110010100100101111: color_data = Z;
		19'b0110010100100110000: color_data = Z;
		19'b0110010100100110001: color_data = Z;
		19'b0110010100100110010: color_data = Z;
		19'b0110010100100110011: color_data = Z;
		19'b0110010100100110100: color_data = Z;
		19'b0110010100100110101: color_data = Z;
		19'b0110010100100110110: color_data = Z;
		19'b0110010100100110111: color_data = Z;
		19'b0110010100100111000: color_data = Z;
		19'b0110010100100111001: color_data = Z;
		19'b0110010100100111010: color_data = Z;
		19'b0110010100100111011: color_data = Z;
		19'b0110010100100111100: color_data = Z;
		19'b0110010100100111101: color_data = Z;
		19'b0110010100100111110: color_data = Z;
		19'b0110010100100111111: color_data = Z;
		19'b0110010100101000000: color_data = Z;
		19'b0110010100101000001: color_data = Z;
		19'b0110010100101000010: color_data = Z;
		19'b0110010100101000011: color_data = Z;
		19'b0110010100101000100: color_data = Z;
		19'b0110010100101000101: color_data = Z;
		19'b0110010100101000110: color_data = Z;
		19'b0110010100101000111: color_data = Z;
		19'b0110010100101001000: color_data = Z;
		19'b0110010100101001001: color_data = Z;
		19'b0110010100101001010: color_data = Z;
		19'b0110010100101001011: color_data = Z;
		19'b0110010100101001100: color_data = Z;
		19'b0110010100101001101: color_data = Z;
		19'b0110010100101001110: color_data = Z;
		19'b0110010100101001111: color_data = Z;
		19'b0110010100101010000: color_data = Z;
		19'b0110010100101010001: color_data = Z;
		19'b0110010100101010010: color_data = Z;
		19'b0110010100101010011: color_data = Z;
		19'b0110010100101010100: color_data = Z;
		19'b0110010100101010101: color_data = Z;
		19'b0110010100101010110: color_data = Z;
		19'b0110010100101010111: color_data = Z;
		19'b0110010100101011000: color_data = Z;
		19'b0110010100101011001: color_data = Z;
		19'b0110010100101011010: color_data = Z;
		19'b0110010100101011011: color_data = Z;
		19'b0110010100101011100: color_data = Z;
		19'b0110010100101011101: color_data = Z;
		19'b0110010100101011110: color_data = Z;
		19'b0110010100101011111: color_data = Z;
		19'b0110010100101100000: color_data = Z;
		19'b0110010100101100001: color_data = Z;
		19'b0110010100101100010: color_data = Z;
		19'b0110010100101100011: color_data = Z;
		19'b0110010100101100100: color_data = Z;
		19'b0110010100101100101: color_data = Z;
		19'b0110010100101100110: color_data = Z;
		19'b0110010100101100111: color_data = Z;
		19'b0110010100101101000: color_data = Z;
		19'b0110010100101101001: color_data = Z;
		19'b0110010100101101010: color_data = Z;
		19'b0110010100101101011: color_data = Z;
		19'b0110010100101101100: color_data = Z;
		19'b0110010100101101101: color_data = Z;
		19'b0110010100101101110: color_data = Z;
		19'b0110010100101101111: color_data = Z;
		19'b0110010100101110000: color_data = Z;
		19'b0110010100101110001: color_data = Z;
		19'b0110010100101110010: color_data = Z;
		19'b0110010100101110011: color_data = Z;
		19'b0110010100101110100: color_data = Z;
		19'b0110010100101110101: color_data = Z;
		19'b0110010100101110110: color_data = Z;
		19'b0110010100101110111: color_data = Z;
		19'b0110010100101111101: color_data = Z;
		19'b0110010100101111110: color_data = Z;
		19'b0110010100101111111: color_data = Z;
		19'b0110010100110000000: color_data = Z;
		19'b0110010100110000001: color_data = Z;
		19'b0110010100110000010: color_data = Z;
		19'b0110010100110000011: color_data = Z;
		19'b0110010100110000100: color_data = Z;
		19'b0110010100110000101: color_data = Z;
		19'b0110010100110000110: color_data = Z;
		19'b0110010100110001101: color_data = Z;
		19'b0110010100110001110: color_data = Z;
		19'b0110010100110001111: color_data = Z;
		19'b0110010100110010000: color_data = Z;
		19'b0110010100110010001: color_data = Z;
		19'b0110010100110010010: color_data = Z;
		19'b0110010100110010011: color_data = Z;
		19'b0110010100111010001: color_data = Z;
		19'b0110010100111010010: color_data = Z;
		19'b0110010100111010011: color_data = Z;
		19'b0110010100111010100: color_data = Z;
		19'b0110010100111010101: color_data = Z;
		19'b0110010100111010110: color_data = Z;
		19'b0110010100111010111: color_data = Z;
		19'b0110010100111011000: color_data = Z;
		19'b0110010100111011001: color_data = Z;
		19'b0110010100111011010: color_data = Z;
		19'b0110010100111011011: color_data = Z;
		19'b0110010110010100001: color_data = Z;
		19'b0110010110100010111: color_data = Z;
		19'b0110010110100011000: color_data = Z;
		19'b0110010110100011001: color_data = Z;
		19'b0110010110100011010: color_data = Z;
		19'b0110010110100011011: color_data = Z;
		19'b0110010110100011100: color_data = Z;
		19'b0110010110100011101: color_data = Z;
		19'b0110010110100011110: color_data = Z;
		19'b0110010110100011111: color_data = Z;
		19'b0110010110100100000: color_data = Z;
		19'b0110010110100100001: color_data = Z;
		19'b0110010110100100010: color_data = Z;
		19'b0110010110100100011: color_data = Z;
		19'b0110010110100100100: color_data = Z;
		19'b0110010110100100101: color_data = Z;
		19'b0110010110100100110: color_data = Z;
		19'b0110010110100100111: color_data = Z;
		19'b0110010110100101000: color_data = Z;
		19'b0110010110100101001: color_data = Z;
		19'b0110010110100101010: color_data = Z;
		19'b0110010110100101011: color_data = Z;
		19'b0110010110100101100: color_data = Z;
		19'b0110010110100101101: color_data = Z;
		19'b0110010110100101110: color_data = Z;
		19'b0110010110100101111: color_data = Z;
		19'b0110010110100110000: color_data = Z;
		19'b0110010110100110001: color_data = Z;
		19'b0110010110100110010: color_data = Z;
		19'b0110010110100110011: color_data = Z;
		19'b0110010110100110100: color_data = Z;
		19'b0110010110100110101: color_data = Z;
		19'b0110010110100110110: color_data = Z;
		19'b0110010110100110111: color_data = Z;
		19'b0110010110100111000: color_data = Z;
		19'b0110010110100111001: color_data = Z;
		19'b0110010110100111010: color_data = Z;
		19'b0110010110100111011: color_data = Z;
		19'b0110010110100111100: color_data = Z;
		19'b0110010110100111101: color_data = Z;
		19'b0110010110100111110: color_data = Z;
		19'b0110010110100111111: color_data = Z;
		19'b0110010110101000000: color_data = Z;
		19'b0110010110101000001: color_data = Z;
		19'b0110010110101000010: color_data = Z;
		19'b0110010110101000011: color_data = Z;
		19'b0110010110101000100: color_data = Z;
		19'b0110010110101000101: color_data = Z;
		19'b0110010110101000110: color_data = Z;
		19'b0110010110101000111: color_data = Z;
		19'b0110010110101001000: color_data = Z;
		19'b0110010110101001001: color_data = Z;
		19'b0110010110101001010: color_data = Z;
		19'b0110010110101001011: color_data = Z;
		19'b0110010110101001100: color_data = Z;
		19'b0110010110101001101: color_data = Z;
		19'b0110010110101001110: color_data = Z;
		19'b0110010110101001111: color_data = Z;
		19'b0110010110101010000: color_data = Z;
		19'b0110010110101010001: color_data = Z;
		19'b0110010110101010010: color_data = Z;
		19'b0110010110101010011: color_data = Z;
		19'b0110010110101010100: color_data = Z;
		19'b0110010110101010101: color_data = Z;
		19'b0110010110101010110: color_data = Z;
		19'b0110010110101010111: color_data = Z;
		19'b0110010110101011000: color_data = Z;
		19'b0110010110101011001: color_data = Z;
		19'b0110010110101011010: color_data = Z;
		19'b0110010110101011011: color_data = Z;
		19'b0110010110101011100: color_data = Z;
		19'b0110010110101011101: color_data = Z;
		19'b0110010110101011110: color_data = Z;
		19'b0110010110101011111: color_data = Z;
		19'b0110010110101100000: color_data = Z;
		19'b0110010110101100001: color_data = Z;
		19'b0110010110101100010: color_data = Z;
		19'b0110010110101100011: color_data = Z;
		19'b0110010110101100100: color_data = Z;
		19'b0110010110101100101: color_data = Z;
		19'b0110010110101100110: color_data = Z;
		19'b0110010110101100111: color_data = Z;
		19'b0110010110101101001: color_data = Z;
		19'b0110010110101101010: color_data = Z;
		19'b0110010110101101011: color_data = Z;
		19'b0110010110101101100: color_data = Z;
		19'b0110010110101101101: color_data = Z;
		19'b0110010110101101110: color_data = Z;
		19'b0110010110101101111: color_data = Z;
		19'b0110010110101110000: color_data = Z;
		19'b0110010110101110001: color_data = Z;
		19'b0110010110101110010: color_data = Z;
		19'b0110010110101110011: color_data = Z;
		19'b0110010110101110100: color_data = Z;
		19'b0110010110101110101: color_data = Z;
		19'b0110010110101110110: color_data = Z;
		19'b0110010110101110111: color_data = Z;
		19'b0110010110101111101: color_data = Z;
		19'b0110010110101111110: color_data = Z;
		19'b0110010110101111111: color_data = Z;
		19'b0110010110110000000: color_data = Z;
		19'b0110010110110000001: color_data = Z;
		19'b0110010110110000010: color_data = Z;
		19'b0110010110110000011: color_data = Z;
		19'b0110010110110000100: color_data = Z;
		19'b0110010110110000101: color_data = Z;
		19'b0110010110110000110: color_data = Z;
		19'b0110010110110000111: color_data = Z;
		19'b0110010110110001101: color_data = Z;
		19'b0110010110110001110: color_data = Z;
		19'b0110010110110001111: color_data = Z;
		19'b0110010110110010000: color_data = Z;
		19'b0110010110110010001: color_data = Z;
		19'b0110010110110010010: color_data = Z;
		19'b0110010110110010011: color_data = Z;
		19'b0110010110110010100: color_data = Z;
		19'b0110010110111010001: color_data = Z;
		19'b0110010110111010010: color_data = Z;
		19'b0110010110111010011: color_data = Z;
		19'b0110010110111010100: color_data = Z;
		19'b0110010110111010101: color_data = Z;
		19'b0110010110111010110: color_data = Z;
		19'b0110010110111010111: color_data = Z;
		19'b0110010110111011000: color_data = Z;
		19'b0110010110111011001: color_data = Z;
		19'b0110010110111011010: color_data = Z;
		19'b0110010110111011011: color_data = Z;
		19'b0110011000100010110: color_data = Z;
		19'b0110011000100010111: color_data = Z;
		19'b0110011000100011000: color_data = Z;
		19'b0110011000100011001: color_data = Z;
		19'b0110011000100011010: color_data = Z;
		19'b0110011000100011011: color_data = Z;
		19'b0110011000100011100: color_data = Z;
		19'b0110011000100011101: color_data = Z;
		19'b0110011000100011110: color_data = Z;
		19'b0110011000100011111: color_data = Z;
		19'b0110011000100100000: color_data = Z;
		19'b0110011000100100001: color_data = Z;
		19'b0110011000100100010: color_data = Z;
		19'b0110011000100100011: color_data = Z;
		19'b0110011000100100100: color_data = Z;
		19'b0110011000100100101: color_data = Z;
		19'b0110011000100100110: color_data = Z;
		19'b0110011000100100111: color_data = Z;
		19'b0110011000100101000: color_data = Z;
		19'b0110011000100101001: color_data = Z;
		19'b0110011000100101010: color_data = Z;
		19'b0110011000100101011: color_data = Z;
		19'b0110011000100101100: color_data = Z;
		19'b0110011000100101101: color_data = Z;
		19'b0110011000100101110: color_data = Z;
		19'b0110011000100101111: color_data = Z;
		19'b0110011000100110000: color_data = Z;
		19'b0110011000100110001: color_data = Z;
		19'b0110011000100110010: color_data = Z;
		19'b0110011000100110011: color_data = Z;
		19'b0110011000100110100: color_data = Z;
		19'b0110011000100110101: color_data = Z;
		19'b0110011000100110110: color_data = Z;
		19'b0110011000100110111: color_data = Z;
		19'b0110011000100111000: color_data = Z;
		19'b0110011000100111001: color_data = Z;
		19'b0110011000100111010: color_data = Z;
		19'b0110011000100111011: color_data = Z;
		19'b0110011000100111100: color_data = Z;
		19'b0110011000100111101: color_data = Z;
		19'b0110011000100111110: color_data = Z;
		19'b0110011000100111111: color_data = Z;
		19'b0110011000101000000: color_data = Z;
		19'b0110011000101000001: color_data = Z;
		19'b0110011000101000010: color_data = Z;
		19'b0110011000101000011: color_data = Z;
		19'b0110011000101000100: color_data = Z;
		19'b0110011000101000101: color_data = Z;
		19'b0110011000101000110: color_data = Z;
		19'b0110011000101000111: color_data = Z;
		19'b0110011000101001000: color_data = Z;
		19'b0110011000101001001: color_data = Z;
		19'b0110011000101001010: color_data = Z;
		19'b0110011000101001011: color_data = Z;
		19'b0110011000101001100: color_data = Z;
		19'b0110011000101001101: color_data = Z;
		19'b0110011000101001110: color_data = Z;
		19'b0110011000101001111: color_data = Z;
		19'b0110011000101010000: color_data = Z;
		19'b0110011000101010001: color_data = Z;
		19'b0110011000101010010: color_data = Z;
		19'b0110011000101010011: color_data = Z;
		19'b0110011000101010100: color_data = Z;
		19'b0110011000101010101: color_data = Z;
		19'b0110011000101010110: color_data = Z;
		19'b0110011000101010111: color_data = Z;
		19'b0110011000101011000: color_data = Z;
		19'b0110011000101011001: color_data = Z;
		19'b0110011000101011010: color_data = Z;
		19'b0110011000101011011: color_data = Z;
		19'b0110011000101011100: color_data = Z;
		19'b0110011000101011101: color_data = Z;
		19'b0110011000101011110: color_data = Z;
		19'b0110011000101011111: color_data = Z;
		19'b0110011000101100000: color_data = Z;
		19'b0110011000101100001: color_data = Z;
		19'b0110011000101100010: color_data = Z;
		19'b0110011000101100011: color_data = Z;
		19'b0110011000101100100: color_data = Z;
		19'b0110011000101100101: color_data = Z;
		19'b0110011000101100110: color_data = Z;
		19'b0110011000101100111: color_data = Z;
		19'b0110011000101101001: color_data = Z;
		19'b0110011000101101010: color_data = Z;
		19'b0110011000101101011: color_data = Z;
		19'b0110011000101101100: color_data = Z;
		19'b0110011000101101101: color_data = Z;
		19'b0110011000101101110: color_data = Z;
		19'b0110011000101101111: color_data = Z;
		19'b0110011000101110000: color_data = Z;
		19'b0110011000101110001: color_data = Z;
		19'b0110011000101110010: color_data = Z;
		19'b0110011000101110011: color_data = Z;
		19'b0110011000101110100: color_data = Z;
		19'b0110011000101110101: color_data = Z;
		19'b0110011000101110110: color_data = Z;
		19'b0110011000101110111: color_data = Z;
		19'b0110011000101111000: color_data = Z;
		19'b0110011000101111110: color_data = Z;
		19'b0110011000101111111: color_data = Z;
		19'b0110011000110000000: color_data = Z;
		19'b0110011000110000001: color_data = Z;
		19'b0110011000110000010: color_data = Z;
		19'b0110011000110000011: color_data = Z;
		19'b0110011000110000100: color_data = Z;
		19'b0110011000110000101: color_data = Z;
		19'b0110011000110000110: color_data = Z;
		19'b0110011000110000111: color_data = Z;
		19'b0110011000110001000: color_data = Z;
		19'b0110011000110001110: color_data = Z;
		19'b0110011000110001111: color_data = Z;
		19'b0110011000110010000: color_data = Z;
		19'b0110011000110010001: color_data = Z;
		19'b0110011000110010010: color_data = Z;
		19'b0110011000110010011: color_data = Z;
		19'b0110011000110010100: color_data = Z;
		19'b0110011000111010001: color_data = Z;
		19'b0110011000111010010: color_data = Z;
		19'b0110011000111010011: color_data = Z;
		19'b0110011000111010100: color_data = Z;
		19'b0110011000111010101: color_data = Z;
		19'b0110011000111010110: color_data = Z;
		19'b0110011000111010111: color_data = Z;
		19'b0110011000111011000: color_data = Z;
		19'b0110011000111011001: color_data = Z;
		19'b0110011000111011010: color_data = Z;
		19'b0110011000111011011: color_data = Z;
		19'b0110011010100010110: color_data = Z;
		19'b0110011010100010111: color_data = Z;
		19'b0110011010100011000: color_data = Z;
		19'b0110011010100011001: color_data = Z;
		19'b0110011010100011010: color_data = Z;
		19'b0110011010100011011: color_data = Z;
		19'b0110011010100011100: color_data = Z;
		19'b0110011010100011101: color_data = Z;
		19'b0110011010100011110: color_data = Z;
		19'b0110011010100011111: color_data = Z;
		19'b0110011010100100000: color_data = Z;
		19'b0110011010100100001: color_data = Z;
		19'b0110011010100100010: color_data = Z;
		19'b0110011010100100011: color_data = Z;
		19'b0110011010100100100: color_data = Z;
		19'b0110011010100100101: color_data = Z;
		19'b0110011010100100110: color_data = Z;
		19'b0110011010100100111: color_data = Z;
		19'b0110011010100101000: color_data = Z;
		19'b0110011010100101001: color_data = Z;
		19'b0110011010100101010: color_data = Z;
		19'b0110011010100101011: color_data = Z;
		19'b0110011010100101100: color_data = Z;
		19'b0110011010100101101: color_data = Z;
		19'b0110011010100101110: color_data = Z;
		19'b0110011010100101111: color_data = Z;
		19'b0110011010100110000: color_data = Z;
		19'b0110011010100110001: color_data = Z;
		19'b0110011010100110010: color_data = Z;
		19'b0110011010100110011: color_data = Z;
		19'b0110011010100110100: color_data = Z;
		19'b0110011010100110101: color_data = Z;
		19'b0110011010100110110: color_data = Z;
		19'b0110011010100110111: color_data = Z;
		19'b0110011010100111000: color_data = Z;
		19'b0110011010100111001: color_data = Z;
		19'b0110011010100111010: color_data = Z;
		19'b0110011010100111011: color_data = Z;
		19'b0110011010100111100: color_data = Z;
		19'b0110011010100111101: color_data = Z;
		19'b0110011010100111110: color_data = Z;
		19'b0110011010100111111: color_data = Z;
		19'b0110011010101000000: color_data = Z;
		19'b0110011010101000001: color_data = Z;
		19'b0110011010101000010: color_data = Z;
		19'b0110011010101000011: color_data = Z;
		19'b0110011010101000100: color_data = Z;
		19'b0110011010101000101: color_data = Z;
		19'b0110011010101000110: color_data = Z;
		19'b0110011010101000111: color_data = Z;
		19'b0110011010101001000: color_data = Z;
		19'b0110011010101001001: color_data = Z;
		19'b0110011010101001010: color_data = Z;
		19'b0110011010101001011: color_data = Z;
		19'b0110011010101001100: color_data = Z;
		19'b0110011010101001101: color_data = Z;
		19'b0110011010101001110: color_data = Z;
		19'b0110011010101001111: color_data = Z;
		19'b0110011010101010000: color_data = Z;
		19'b0110011010101010001: color_data = Z;
		19'b0110011010101010010: color_data = Z;
		19'b0110011010101010011: color_data = Z;
		19'b0110011010101010100: color_data = Z;
		19'b0110011010101010101: color_data = Z;
		19'b0110011010101010110: color_data = Z;
		19'b0110011010101010111: color_data = Z;
		19'b0110011010101011000: color_data = Z;
		19'b0110011010101011001: color_data = Z;
		19'b0110011010101011010: color_data = Z;
		19'b0110011010101011011: color_data = Z;
		19'b0110011010101011100: color_data = Z;
		19'b0110011010101011101: color_data = Z;
		19'b0110011010101011110: color_data = Z;
		19'b0110011010101011111: color_data = Z;
		19'b0110011010101100000: color_data = Z;
		19'b0110011010101100001: color_data = Z;
		19'b0110011010101100010: color_data = Z;
		19'b0110011010101100011: color_data = Z;
		19'b0110011010101100100: color_data = Z;
		19'b0110011010101100101: color_data = Z;
		19'b0110011010101100110: color_data = Z;
		19'b0110011010101100111: color_data = Z;
		19'b0110011010101101001: color_data = Z;
		19'b0110011010101101010: color_data = Z;
		19'b0110011010101101011: color_data = Z;
		19'b0110011010101101100: color_data = Z;
		19'b0110011010101101101: color_data = Z;
		19'b0110011010101101110: color_data = Z;
		19'b0110011010101101111: color_data = Z;
		19'b0110011010101110000: color_data = Z;
		19'b0110011010101110001: color_data = Z;
		19'b0110011010101110010: color_data = Z;
		19'b0110011010101110011: color_data = Z;
		19'b0110011010101110100: color_data = Z;
		19'b0110011010101110101: color_data = Z;
		19'b0110011010101110110: color_data = Z;
		19'b0110011010101110111: color_data = Z;
		19'b0110011010101111000: color_data = Z;
		19'b0110011010101111110: color_data = Z;
		19'b0110011010101111111: color_data = Z;
		19'b0110011010110000000: color_data = Z;
		19'b0110011010110000001: color_data = Z;
		19'b0110011010110000010: color_data = Z;
		19'b0110011010110000011: color_data = Z;
		19'b0110011010110000100: color_data = Z;
		19'b0110011010110000101: color_data = Z;
		19'b0110011010110000110: color_data = Z;
		19'b0110011010110000111: color_data = Z;
		19'b0110011010110001000: color_data = Z;
		19'b0110011010110001001: color_data = Z;
		19'b0110011010110001111: color_data = Z;
		19'b0110011010110010000: color_data = Z;
		19'b0110011010110010001: color_data = Z;
		19'b0110011010110010010: color_data = Z;
		19'b0110011010110010011: color_data = Z;
		19'b0110011010110010100: color_data = Z;
		19'b0110011010111010010: color_data = Z;
		19'b0110011010111010011: color_data = Z;
		19'b0110011010111010100: color_data = Z;
		19'b0110011010111010101: color_data = Z;
		19'b0110011010111010110: color_data = Z;
		19'b0110011010111010111: color_data = Z;
		19'b0110011010111011000: color_data = Z;
		19'b0110011010111011001: color_data = Z;
		19'b0110011010111011010: color_data = Z;
		19'b0110011010111011011: color_data = Z;
		19'b0110011100010100001: color_data = Z;
		19'b0110011100010100010: color_data = Z;
		19'b0110011100010100100: color_data = Z;
		19'b0110011100010100101: color_data = Z;
		19'b0110011100010100110: color_data = Z;
		19'b0110011100010100111: color_data = Z;
		19'b0110011100010101000: color_data = Z;
		19'b0110011100100010101: color_data = Z;
		19'b0110011100100010110: color_data = Z;
		19'b0110011100100010111: color_data = Z;
		19'b0110011100100011000: color_data = Z;
		19'b0110011100100011001: color_data = Z;
		19'b0110011100100011010: color_data = Z;
		19'b0110011100100011011: color_data = Z;
		19'b0110011100100011100: color_data = Z;
		19'b0110011100100011101: color_data = Z;
		19'b0110011100100011110: color_data = Z;
		19'b0110011100100011111: color_data = Z;
		19'b0110011100100100000: color_data = Z;
		19'b0110011100100100001: color_data = Z;
		19'b0110011100100100010: color_data = Z;
		19'b0110011100100100011: color_data = Z;
		19'b0110011100100100100: color_data = Z;
		19'b0110011100100100101: color_data = Z;
		19'b0110011100100100110: color_data = Z;
		19'b0110011100100100111: color_data = Z;
		19'b0110011100100101000: color_data = Z;
		19'b0110011100100101001: color_data = Z;
		19'b0110011100100101010: color_data = Z;
		19'b0110011100100101011: color_data = Z;
		19'b0110011100100101100: color_data = Z;
		19'b0110011100100101101: color_data = Z;
		19'b0110011100100101110: color_data = Z;
		19'b0110011100100101111: color_data = Z;
		19'b0110011100100110000: color_data = Z;
		19'b0110011100100110001: color_data = Z;
		19'b0110011100100110010: color_data = Z;
		19'b0110011100100110011: color_data = Z;
		19'b0110011100100110100: color_data = Z;
		19'b0110011100100110101: color_data = Z;
		19'b0110011100100110110: color_data = Z;
		19'b0110011100100110111: color_data = Z;
		19'b0110011100100111000: color_data = Z;
		19'b0110011100100111001: color_data = Z;
		19'b0110011100100111010: color_data = Z;
		19'b0110011100100111011: color_data = Z;
		19'b0110011100100111100: color_data = Z;
		19'b0110011100100111101: color_data = Z;
		19'b0110011100100111110: color_data = Z;
		19'b0110011100100111111: color_data = Z;
		19'b0110011100101000000: color_data = Z;
		19'b0110011100101000001: color_data = Z;
		19'b0110011100101000010: color_data = Z;
		19'b0110011100101000011: color_data = Z;
		19'b0110011100101000100: color_data = Z;
		19'b0110011100101000101: color_data = Z;
		19'b0110011100101000110: color_data = Z;
		19'b0110011100101000111: color_data = Z;
		19'b0110011100101001000: color_data = Z;
		19'b0110011100101001001: color_data = Z;
		19'b0110011100101001010: color_data = Z;
		19'b0110011100101001011: color_data = Z;
		19'b0110011100101001100: color_data = Z;
		19'b0110011100101001101: color_data = Z;
		19'b0110011100101001110: color_data = Z;
		19'b0110011100101001111: color_data = Z;
		19'b0110011100101010000: color_data = Z;
		19'b0110011100101010001: color_data = Z;
		19'b0110011100101010010: color_data = Z;
		19'b0110011100101010011: color_data = Z;
		19'b0110011100101010100: color_data = Z;
		19'b0110011100101010101: color_data = Z;
		19'b0110011100101010110: color_data = Z;
		19'b0110011100101010111: color_data = Z;
		19'b0110011100101011000: color_data = Z;
		19'b0110011100101011001: color_data = Z;
		19'b0110011100101011010: color_data = Z;
		19'b0110011100101011011: color_data = Z;
		19'b0110011100101011100: color_data = Z;
		19'b0110011100101011101: color_data = Z;
		19'b0110011100101011110: color_data = Z;
		19'b0110011100101011111: color_data = Z;
		19'b0110011100101100000: color_data = Z;
		19'b0110011100101100001: color_data = Z;
		19'b0110011100101100010: color_data = Z;
		19'b0110011100101100011: color_data = Z;
		19'b0110011100101100100: color_data = Z;
		19'b0110011100101100101: color_data = Z;
		19'b0110011100101100110: color_data = Z;
		19'b0110011100101100111: color_data = Z;
		19'b0110011100101101001: color_data = Z;
		19'b0110011100101101010: color_data = Z;
		19'b0110011100101101011: color_data = Z;
		19'b0110011100101101100: color_data = Z;
		19'b0110011100101101101: color_data = Z;
		19'b0110011100101101110: color_data = Z;
		19'b0110011100101101111: color_data = Z;
		19'b0110011100101110000: color_data = Z;
		19'b0110011100101110001: color_data = Z;
		19'b0110011100101110010: color_data = Z;
		19'b0110011100101110011: color_data = Z;
		19'b0110011100101110100: color_data = Z;
		19'b0110011100101110101: color_data = Z;
		19'b0110011100101110110: color_data = Z;
		19'b0110011100101110111: color_data = Z;
		19'b0110011100101111000: color_data = Z;
		19'b0110011100101111001: color_data = Z;
		19'b0110011100101111101: color_data = Z;
		19'b0110011100101111110: color_data = Z;
		19'b0110011100101111111: color_data = Z;
		19'b0110011100110000000: color_data = Z;
		19'b0110011100110000001: color_data = Z;
		19'b0110011100110000010: color_data = Z;
		19'b0110011100110000011: color_data = Z;
		19'b0110011100110000100: color_data = Z;
		19'b0110011100110000101: color_data = Z;
		19'b0110011100110000110: color_data = Z;
		19'b0110011100110000111: color_data = Z;
		19'b0110011100110001000: color_data = Z;
		19'b0110011100110001001: color_data = Z;
		19'b0110011100110001111: color_data = Z;
		19'b0110011100110010000: color_data = Z;
		19'b0110011100110010001: color_data = Z;
		19'b0110011100110010010: color_data = Z;
		19'b0110011100110010011: color_data = Z;
		19'b0110011100110010100: color_data = Z;
		19'b0110011100111010010: color_data = Z;
		19'b0110011100111010011: color_data = Z;
		19'b0110011100111010100: color_data = Z;
		19'b0110011100111010101: color_data = Z;
		19'b0110011100111010110: color_data = Z;
		19'b0110011100111010111: color_data = Z;
		19'b0110011100111011000: color_data = Z;
		19'b0110011100111011001: color_data = Z;
		19'b0110011100111011010: color_data = Z;
		19'b0110011110010100001: color_data = Z;
		19'b0110011110010100010: color_data = Z;
		19'b0110011110010100011: color_data = Z;
		19'b0110011110010100100: color_data = Z;
		19'b0110011110010100101: color_data = Z;
		19'b0110011110010100110: color_data = Z;
		19'b0110011110010100111: color_data = Z;
		19'b0110011110010101000: color_data = Z;
		19'b0110011110100010011: color_data = Z;
		19'b0110011110100010100: color_data = Z;
		19'b0110011110100010101: color_data = Z;
		19'b0110011110100010110: color_data = Z;
		19'b0110011110100010111: color_data = Z;
		19'b0110011110100011000: color_data = Z;
		19'b0110011110100011001: color_data = Z;
		19'b0110011110100011010: color_data = Z;
		19'b0110011110100011011: color_data = Z;
		19'b0110011110100011100: color_data = Z;
		19'b0110011110100011101: color_data = Z;
		19'b0110011110100011110: color_data = Z;
		19'b0110011110100011111: color_data = Z;
		19'b0110011110100100000: color_data = Z;
		19'b0110011110100100001: color_data = Z;
		19'b0110011110100100010: color_data = Z;
		19'b0110011110100100011: color_data = Z;
		19'b0110011110100100100: color_data = Z;
		19'b0110011110100100101: color_data = Z;
		19'b0110011110100100110: color_data = Z;
		19'b0110011110100100111: color_data = Z;
		19'b0110011110100101000: color_data = Z;
		19'b0110011110100101001: color_data = Z;
		19'b0110011110100101010: color_data = Z;
		19'b0110011110100101011: color_data = Z;
		19'b0110011110100101100: color_data = Z;
		19'b0110011110100101101: color_data = Z;
		19'b0110011110100101110: color_data = Z;
		19'b0110011110100101111: color_data = Z;
		19'b0110011110100110000: color_data = Z;
		19'b0110011110100110001: color_data = Z;
		19'b0110011110100110010: color_data = Z;
		19'b0110011110100110011: color_data = Z;
		19'b0110011110100110100: color_data = Z;
		19'b0110011110100110101: color_data = Z;
		19'b0110011110100110110: color_data = Z;
		19'b0110011110100110111: color_data = Z;
		19'b0110011110100111000: color_data = Z;
		19'b0110011110100111001: color_data = Z;
		19'b0110011110100111010: color_data = Z;
		19'b0110011110100111011: color_data = Z;
		19'b0110011110100111100: color_data = Z;
		19'b0110011110100111101: color_data = Z;
		19'b0110011110100111110: color_data = Z;
		19'b0110011110100111111: color_data = Z;
		19'b0110011110101000000: color_data = Z;
		19'b0110011110101000001: color_data = Z;
		19'b0110011110101000010: color_data = Z;
		19'b0110011110101000011: color_data = Z;
		19'b0110011110101000100: color_data = Z;
		19'b0110011110101000101: color_data = Z;
		19'b0110011110101000110: color_data = Z;
		19'b0110011110101000111: color_data = Z;
		19'b0110011110101001000: color_data = Z;
		19'b0110011110101001001: color_data = Z;
		19'b0110011110101001010: color_data = Z;
		19'b0110011110101001011: color_data = Z;
		19'b0110011110101001100: color_data = Z;
		19'b0110011110101001101: color_data = Z;
		19'b0110011110101001110: color_data = Z;
		19'b0110011110101001111: color_data = Z;
		19'b0110011110101010000: color_data = Z;
		19'b0110011110101010001: color_data = Z;
		19'b0110011110101010010: color_data = Z;
		19'b0110011110101010011: color_data = Z;
		19'b0110011110101010100: color_data = Z;
		19'b0110011110101010101: color_data = Z;
		19'b0110011110101010110: color_data = Z;
		19'b0110011110101010111: color_data = Z;
		19'b0110011110101011000: color_data = Z;
		19'b0110011110101011001: color_data = Z;
		19'b0110011110101011010: color_data = Z;
		19'b0110011110101011011: color_data = Z;
		19'b0110011110101011100: color_data = Z;
		19'b0110011110101011101: color_data = Z;
		19'b0110011110101011110: color_data = Z;
		19'b0110011110101011111: color_data = Z;
		19'b0110011110101100000: color_data = Z;
		19'b0110011110101100001: color_data = Z;
		19'b0110011110101100010: color_data = Z;
		19'b0110011110101100011: color_data = Z;
		19'b0110011110101100100: color_data = Z;
		19'b0110011110101100101: color_data = Z;
		19'b0110011110101100110: color_data = Z;
		19'b0110011110101100111: color_data = Z;
		19'b0110011110101101010: color_data = Z;
		19'b0110011110101101011: color_data = Z;
		19'b0110011110101101100: color_data = Z;
		19'b0110011110101101101: color_data = Z;
		19'b0110011110101101110: color_data = Z;
		19'b0110011110101101111: color_data = Z;
		19'b0110011110101110000: color_data = Z;
		19'b0110011110101110001: color_data = Z;
		19'b0110011110101110010: color_data = Z;
		19'b0110011110101110011: color_data = Z;
		19'b0110011110101110100: color_data = Z;
		19'b0110011110101110101: color_data = Z;
		19'b0110011110101110110: color_data = Z;
		19'b0110011110101110111: color_data = Z;
		19'b0110011110101111000: color_data = Z;
		19'b0110011110101111001: color_data = Z;
		19'b0110011110101111101: color_data = Z;
		19'b0110011110101111110: color_data = Z;
		19'b0110011110101111111: color_data = Z;
		19'b0110011110110000000: color_data = Z;
		19'b0110011110110000001: color_data = Z;
		19'b0110011110110000010: color_data = Z;
		19'b0110011110110000011: color_data = Z;
		19'b0110011110110000100: color_data = Z;
		19'b0110011110110000101: color_data = Z;
		19'b0110011110110000110: color_data = Z;
		19'b0110011110110000111: color_data = Z;
		19'b0110011110110001000: color_data = Z;
		19'b0110011110110001001: color_data = Z;
		19'b0110011110110001010: color_data = Z;
		19'b0110011110110001111: color_data = Z;
		19'b0110011110110010000: color_data = Z;
		19'b0110011110110010001: color_data = Z;
		19'b0110011110110010010: color_data = Z;
		19'b0110011110110010011: color_data = Z;
		19'b0110011110110010100: color_data = Z;
		19'b0110011110110010101: color_data = Z;
		19'b0110011110111010010: color_data = Z;
		19'b0110011110111010011: color_data = Z;
		19'b0110011110111010100: color_data = Z;
		19'b0110011110111010101: color_data = Z;
		19'b0110011110111010110: color_data = Z;
		19'b0110011110111010111: color_data = Z;
		19'b0110011110111011000: color_data = Z;
		19'b0110011110111011001: color_data = Z;
		19'b0110011110111011010: color_data = Z;
		19'b0110100000010100010: color_data = Z;
		19'b0110100000010100011: color_data = Z;
		19'b0110100000010100100: color_data = Z;
		19'b0110100000010100101: color_data = Z;
		19'b0110100000010100110: color_data = Z;
		19'b0110100000010100111: color_data = Z;
		19'b0110100000010101000: color_data = Z;
		19'b0110100000100010010: color_data = Z;
		19'b0110100000100010011: color_data = Z;
		19'b0110100000100010100: color_data = Z;
		19'b0110100000100010101: color_data = Z;
		19'b0110100000100010110: color_data = Z;
		19'b0110100000100010111: color_data = Z;
		19'b0110100000100011000: color_data = Z;
		19'b0110100000100011001: color_data = Z;
		19'b0110100000100011010: color_data = Z;
		19'b0110100000100011011: color_data = Z;
		19'b0110100000100011100: color_data = Z;
		19'b0110100000100011101: color_data = Z;
		19'b0110100000100011110: color_data = Z;
		19'b0110100000100011111: color_data = Z;
		19'b0110100000100100000: color_data = Z;
		19'b0110100000100100001: color_data = Z;
		19'b0110100000100100010: color_data = Z;
		19'b0110100000100100011: color_data = Z;
		19'b0110100000100100100: color_data = Z;
		19'b0110100000100100101: color_data = Z;
		19'b0110100000100100110: color_data = Z;
		19'b0110100000100100111: color_data = Z;
		19'b0110100000100101000: color_data = Z;
		19'b0110100000100101001: color_data = Z;
		19'b0110100000100101010: color_data = Z;
		19'b0110100000100101011: color_data = Z;
		19'b0110100000100101100: color_data = Z;
		19'b0110100000100101101: color_data = Z;
		19'b0110100000100101110: color_data = Z;
		19'b0110100000100101111: color_data = Z;
		19'b0110100000100110000: color_data = Z;
		19'b0110100000100110001: color_data = Z;
		19'b0110100000100110010: color_data = Z;
		19'b0110100000100110011: color_data = Z;
		19'b0110100000100110100: color_data = Z;
		19'b0110100000100110101: color_data = Z;
		19'b0110100000100110110: color_data = Z;
		19'b0110100000100110111: color_data = Z;
		19'b0110100000100111000: color_data = Z;
		19'b0110100000100111001: color_data = Z;
		19'b0110100000100111010: color_data = Z;
		19'b0110100000100111011: color_data = Z;
		19'b0110100000100111100: color_data = Z;
		19'b0110100000100111101: color_data = Z;
		19'b0110100000100111110: color_data = Z;
		19'b0110100000100111111: color_data = Z;
		19'b0110100000101000000: color_data = Z;
		19'b0110100000101000001: color_data = Z;
		19'b0110100000101000010: color_data = Z;
		19'b0110100000101000011: color_data = Z;
		19'b0110100000101000100: color_data = Z;
		19'b0110100000101000101: color_data = Z;
		19'b0110100000101000110: color_data = Z;
		19'b0110100000101000111: color_data = Z;
		19'b0110100000101001000: color_data = Z;
		19'b0110100000101001001: color_data = Z;
		19'b0110100000101001010: color_data = Z;
		19'b0110100000101001011: color_data = Z;
		19'b0110100000101001100: color_data = Z;
		19'b0110100000101001101: color_data = Z;
		19'b0110100000101001110: color_data = Z;
		19'b0110100000101001111: color_data = Z;
		19'b0110100000101010000: color_data = Z;
		19'b0110100000101010001: color_data = Z;
		19'b0110100000101010010: color_data = Z;
		19'b0110100000101010011: color_data = Z;
		19'b0110100000101010100: color_data = Z;
		19'b0110100000101010101: color_data = Z;
		19'b0110100000101010110: color_data = Z;
		19'b0110100000101010111: color_data = Z;
		19'b0110100000101011000: color_data = Z;
		19'b0110100000101011001: color_data = Z;
		19'b0110100000101011010: color_data = Z;
		19'b0110100000101011011: color_data = Z;
		19'b0110100000101011100: color_data = Z;
		19'b0110100000101011101: color_data = Z;
		19'b0110100000101011110: color_data = Z;
		19'b0110100000101011111: color_data = Z;
		19'b0110100000101100000: color_data = Z;
		19'b0110100000101100001: color_data = Z;
		19'b0110100000101100010: color_data = Z;
		19'b0110100000101100011: color_data = Z;
		19'b0110100000101100100: color_data = Z;
		19'b0110100000101100101: color_data = Z;
		19'b0110100000101100110: color_data = Z;
		19'b0110100000101100111: color_data = Z;
		19'b0110100000101101010: color_data = Z;
		19'b0110100000101101011: color_data = Z;
		19'b0110100000101101100: color_data = Z;
		19'b0110100000101101101: color_data = Z;
		19'b0110100000101101110: color_data = Z;
		19'b0110100000101101111: color_data = Z;
		19'b0110100000101110000: color_data = Z;
		19'b0110100000101110001: color_data = Z;
		19'b0110100000101110010: color_data = Z;
		19'b0110100000101110011: color_data = Z;
		19'b0110100000101110100: color_data = Z;
		19'b0110100000101110101: color_data = Z;
		19'b0110100000101110110: color_data = Z;
		19'b0110100000101110111: color_data = Z;
		19'b0110100000101111000: color_data = Z;
		19'b0110100000101111001: color_data = Z;
		19'b0110100000101111101: color_data = Z;
		19'b0110100000101111110: color_data = Z;
		19'b0110100000101111111: color_data = Z;
		19'b0110100000110000000: color_data = Z;
		19'b0110100000110000001: color_data = Z;
		19'b0110100000110000010: color_data = Z;
		19'b0110100000110000011: color_data = Z;
		19'b0110100000110000100: color_data = Z;
		19'b0110100000110000101: color_data = Z;
		19'b0110100000110000110: color_data = Z;
		19'b0110100000110000111: color_data = Z;
		19'b0110100000110001000: color_data = Z;
		19'b0110100000110001001: color_data = Z;
		19'b0110100000110001010: color_data = Z;
		19'b0110100000110001011: color_data = Z;
		19'b0110100000110001110: color_data = Z;
		19'b0110100000110001111: color_data = Z;
		19'b0110100000110010000: color_data = Z;
		19'b0110100000110010001: color_data = Z;
		19'b0110100000110010010: color_data = Z;
		19'b0110100000110010011: color_data = Z;
		19'b0110100000110010100: color_data = Z;
		19'b0110100000110010101: color_data = Z;
		19'b0110100000111010001: color_data = Z;
		19'b0110100000111010010: color_data = Z;
		19'b0110100000111010011: color_data = Z;
		19'b0110100000111010100: color_data = Z;
		19'b0110100000111010101: color_data = Z;
		19'b0110100000111010110: color_data = Z;
		19'b0110100000111010111: color_data = Z;
		19'b0110100000111011000: color_data = Z;
		19'b0110100000111011001: color_data = Z;
		19'b0110100000111011010: color_data = Z;
		19'b0110100010010100010: color_data = Z;
		19'b0110100010010100011: color_data = Z;
		19'b0110100010010100100: color_data = Z;
		19'b0110100010010100101: color_data = Z;
		19'b0110100010010100110: color_data = Z;
		19'b0110100010010100111: color_data = Z;
		19'b0110100010010101000: color_data = Z;
		19'b0110100010100010001: color_data = Z;
		19'b0110100010100010010: color_data = Z;
		19'b0110100010100010011: color_data = Z;
		19'b0110100010100010100: color_data = Z;
		19'b0110100010100010101: color_data = Z;
		19'b0110100010100010110: color_data = Z;
		19'b0110100010100010111: color_data = Z;
		19'b0110100010100011000: color_data = Z;
		19'b0110100010100011001: color_data = Z;
		19'b0110100010100011010: color_data = Z;
		19'b0110100010100011100: color_data = Z;
		19'b0110100010100011101: color_data = Z;
		19'b0110100010100011110: color_data = Z;
		19'b0110100010100011111: color_data = Z;
		19'b0110100010100100000: color_data = Z;
		19'b0110100010100100001: color_data = Z;
		19'b0110100010100100010: color_data = Z;
		19'b0110100010100100011: color_data = Z;
		19'b0110100010100100100: color_data = Z;
		19'b0110100010100100101: color_data = Z;
		19'b0110100010100100110: color_data = Z;
		19'b0110100010100100111: color_data = Z;
		19'b0110100010100101000: color_data = Z;
		19'b0110100010100101001: color_data = Z;
		19'b0110100010100101010: color_data = Z;
		19'b0110100010100101011: color_data = Z;
		19'b0110100010100101100: color_data = Z;
		19'b0110100010100101101: color_data = Z;
		19'b0110100010100101110: color_data = Z;
		19'b0110100010100101111: color_data = Z;
		19'b0110100010100110000: color_data = Z;
		19'b0110100010100110001: color_data = Z;
		19'b0110100010100110010: color_data = Z;
		19'b0110100010100110011: color_data = Z;
		19'b0110100010100110100: color_data = Z;
		19'b0110100010100110101: color_data = Z;
		19'b0110100010100110110: color_data = Z;
		19'b0110100010100110111: color_data = Z;
		19'b0110100010100111000: color_data = Z;
		19'b0110100010100111001: color_data = Z;
		19'b0110100010100111010: color_data = Z;
		19'b0110100010100111011: color_data = Z;
		19'b0110100010100111100: color_data = Z;
		19'b0110100010100111101: color_data = Z;
		19'b0110100010100111110: color_data = Z;
		19'b0110100010100111111: color_data = Z;
		19'b0110100010101000000: color_data = Z;
		19'b0110100010101000001: color_data = Z;
		19'b0110100010101000010: color_data = Z;
		19'b0110100010101000011: color_data = Z;
		19'b0110100010101000100: color_data = Z;
		19'b0110100010101000101: color_data = Z;
		19'b0110100010101000110: color_data = Z;
		19'b0110100010101000111: color_data = Z;
		19'b0110100010101001000: color_data = Z;
		19'b0110100010101001001: color_data = Z;
		19'b0110100010101001010: color_data = Z;
		19'b0110100010101001011: color_data = Z;
		19'b0110100010101001100: color_data = Z;
		19'b0110100010101001101: color_data = Z;
		19'b0110100010101001110: color_data = Z;
		19'b0110100010101001111: color_data = Z;
		19'b0110100010101010000: color_data = Z;
		19'b0110100010101010001: color_data = Z;
		19'b0110100010101010010: color_data = Z;
		19'b0110100010101010011: color_data = Z;
		19'b0110100010101010100: color_data = Z;
		19'b0110100010101010101: color_data = Z;
		19'b0110100010101010110: color_data = Z;
		19'b0110100010101010111: color_data = Z;
		19'b0110100010101011000: color_data = Z;
		19'b0110100010101011001: color_data = Z;
		19'b0110100010101011010: color_data = Z;
		19'b0110100010101011011: color_data = Z;
		19'b0110100010101011100: color_data = Z;
		19'b0110100010101011101: color_data = Z;
		19'b0110100010101011110: color_data = Z;
		19'b0110100010101011111: color_data = Z;
		19'b0110100010101100000: color_data = Z;
		19'b0110100010101100001: color_data = Z;
		19'b0110100010101100010: color_data = Z;
		19'b0110100010101100011: color_data = Z;
		19'b0110100010101100100: color_data = Z;
		19'b0110100010101100101: color_data = Z;
		19'b0110100010101100110: color_data = Z;
		19'b0110100010101100111: color_data = Z;
		19'b0110100010101101011: color_data = Z;
		19'b0110100010101101100: color_data = Z;
		19'b0110100010101101101: color_data = Z;
		19'b0110100010101101110: color_data = Z;
		19'b0110100010101101111: color_data = Z;
		19'b0110100010101110000: color_data = Z;
		19'b0110100010101110001: color_data = Z;
		19'b0110100010101110010: color_data = Z;
		19'b0110100010101110011: color_data = Z;
		19'b0110100010101110100: color_data = Z;
		19'b0110100010101110101: color_data = Z;
		19'b0110100010101110110: color_data = Z;
		19'b0110100010101110111: color_data = Z;
		19'b0110100010101111000: color_data = Z;
		19'b0110100010101111001: color_data = Z;
		19'b0110100010101111110: color_data = Z;
		19'b0110100010101111111: color_data = Z;
		19'b0110100010110000000: color_data = Z;
		19'b0110100010110000001: color_data = Z;
		19'b0110100010110000010: color_data = Z;
		19'b0110100010110000011: color_data = Z;
		19'b0110100010110000100: color_data = Z;
		19'b0110100010110000101: color_data = Z;
		19'b0110100010110000110: color_data = Z;
		19'b0110100010110000111: color_data = Z;
		19'b0110100010110001000: color_data = Z;
		19'b0110100010110001001: color_data = Z;
		19'b0110100010110001010: color_data = Z;
		19'b0110100010110001011: color_data = Z;
		19'b0110100010110001100: color_data = Z;
		19'b0110100010110001111: color_data = Z;
		19'b0110100010110010000: color_data = Z;
		19'b0110100010110010001: color_data = Z;
		19'b0110100010110010010: color_data = Z;
		19'b0110100010110010011: color_data = Z;
		19'b0110100010110010100: color_data = Z;
		19'b0110100010110010101: color_data = Z;
		19'b0110100010111010001: color_data = Z;
		19'b0110100010111010010: color_data = Z;
		19'b0110100010111010011: color_data = Z;
		19'b0110100010111010100: color_data = Z;
		19'b0110100010111010101: color_data = Z;
		19'b0110100010111010110: color_data = Z;
		19'b0110100010111010111: color_data = Z;
		19'b0110100010111011000: color_data = Z;
		19'b0110100010111011001: color_data = Z;
		19'b0110100010111011010: color_data = Z;
		19'b0110100100010100011: color_data = Z;
		19'b0110100100010100100: color_data = Z;
		19'b0110100100010100101: color_data = Z;
		19'b0110100100010100110: color_data = Z;
		19'b0110100100010100111: color_data = Z;
		19'b0110100100010101000: color_data = Z;
		19'b0110100100100001110: color_data = Z;
		19'b0110100100100001111: color_data = Z;
		19'b0110100100100010000: color_data = Z;
		19'b0110100100100010001: color_data = Z;
		19'b0110100100100010010: color_data = Z;
		19'b0110100100100010011: color_data = Z;
		19'b0110100100100010100: color_data = Z;
		19'b0110100100100010101: color_data = Z;
		19'b0110100100100010110: color_data = Z;
		19'b0110100100100010111: color_data = Z;
		19'b0110100100100011000: color_data = Z;
		19'b0110100100100011001: color_data = Z;
		19'b0110100100100011010: color_data = Z;
		19'b0110100100100011100: color_data = Z;
		19'b0110100100100011101: color_data = Z;
		19'b0110100100100011110: color_data = Z;
		19'b0110100100100011111: color_data = Z;
		19'b0110100100100100000: color_data = Z;
		19'b0110100100100100001: color_data = Z;
		19'b0110100100100100010: color_data = Z;
		19'b0110100100100100011: color_data = Z;
		19'b0110100100100100100: color_data = Z;
		19'b0110100100100100101: color_data = Z;
		19'b0110100100100100110: color_data = Z;
		19'b0110100100100100111: color_data = Z;
		19'b0110100100100101000: color_data = Z;
		19'b0110100100100101001: color_data = Z;
		19'b0110100100100101010: color_data = Z;
		19'b0110100100100101011: color_data = Z;
		19'b0110100100100101100: color_data = Z;
		19'b0110100100100101101: color_data = Z;
		19'b0110100100100101110: color_data = Z;
		19'b0110100100100101111: color_data = Z;
		19'b0110100100100110000: color_data = Z;
		19'b0110100100100110001: color_data = Z;
		19'b0110100100100110010: color_data = Z;
		19'b0110100100100110011: color_data = Z;
		19'b0110100100100110100: color_data = Z;
		19'b0110100100100110101: color_data = Z;
		19'b0110100100100110110: color_data = Z;
		19'b0110100100100110111: color_data = Z;
		19'b0110100100100111000: color_data = Z;
		19'b0110100100100111001: color_data = Z;
		19'b0110100100100111010: color_data = Z;
		19'b0110100100100111011: color_data = Z;
		19'b0110100100100111100: color_data = Z;
		19'b0110100100100111101: color_data = Z;
		19'b0110100100100111110: color_data = Z;
		19'b0110100100100111111: color_data = Z;
		19'b0110100100101000000: color_data = Z;
		19'b0110100100101000001: color_data = Z;
		19'b0110100100101000010: color_data = Z;
		19'b0110100100101000011: color_data = Z;
		19'b0110100100101000100: color_data = Z;
		19'b0110100100101000101: color_data = Z;
		19'b0110100100101000110: color_data = Z;
		19'b0110100100101000111: color_data = Z;
		19'b0110100100101001000: color_data = Z;
		19'b0110100100101001001: color_data = Z;
		19'b0110100100101001010: color_data = Z;
		19'b0110100100101001011: color_data = Z;
		19'b0110100100101001100: color_data = Z;
		19'b0110100100101001101: color_data = Z;
		19'b0110100100101001110: color_data = Z;
		19'b0110100100101001111: color_data = Z;
		19'b0110100100101010000: color_data = Z;
		19'b0110100100101010001: color_data = Z;
		19'b0110100100101010010: color_data = Z;
		19'b0110100100101010011: color_data = Z;
		19'b0110100100101010100: color_data = Z;
		19'b0110100100101010101: color_data = Z;
		19'b0110100100101010110: color_data = Z;
		19'b0110100100101010111: color_data = Z;
		19'b0110100100101011000: color_data = Z;
		19'b0110100100101011001: color_data = Z;
		19'b0110100100101011010: color_data = Z;
		19'b0110100100101011011: color_data = Z;
		19'b0110100100101011100: color_data = Z;
		19'b0110100100101011101: color_data = Z;
		19'b0110100100101011110: color_data = Z;
		19'b0110100100101011111: color_data = Z;
		19'b0110100100101100000: color_data = Z;
		19'b0110100100101100001: color_data = Z;
		19'b0110100100101100010: color_data = Z;
		19'b0110100100101100011: color_data = Z;
		19'b0110100100101100100: color_data = Z;
		19'b0110100100101100101: color_data = Z;
		19'b0110100100101100110: color_data = Z;
		19'b0110100100101100111: color_data = Z;
		19'b0110100100101101011: color_data = Z;
		19'b0110100100101101100: color_data = Z;
		19'b0110100100101101101: color_data = Z;
		19'b0110100100101101110: color_data = Z;
		19'b0110100100101101111: color_data = Z;
		19'b0110100100101110000: color_data = Z;
		19'b0110100100101110001: color_data = Z;
		19'b0110100100101110010: color_data = Z;
		19'b0110100100101110011: color_data = Z;
		19'b0110100100101110100: color_data = Z;
		19'b0110100100101110101: color_data = Z;
		19'b0110100100101110110: color_data = Z;
		19'b0110100100101110111: color_data = Z;
		19'b0110100100101111000: color_data = Z;
		19'b0110100100101111001: color_data = Z;
		19'b0110100100101111110: color_data = Z;
		19'b0110100100101111111: color_data = Z;
		19'b0110100100110000000: color_data = Z;
		19'b0110100100110000001: color_data = Z;
		19'b0110100100110000010: color_data = Z;
		19'b0110100100110000011: color_data = Z;
		19'b0110100100110000100: color_data = Z;
		19'b0110100100110000101: color_data = Z;
		19'b0110100100110000110: color_data = Z;
		19'b0110100100110000111: color_data = Z;
		19'b0110100100110001000: color_data = Z;
		19'b0110100100110001001: color_data = Z;
		19'b0110100100110001010: color_data = Z;
		19'b0110100100110001011: color_data = Z;
		19'b0110100100110001100: color_data = Z;
		19'b0110100100110001101: color_data = Z;
		19'b0110100100110001110: color_data = Z;
		19'b0110100100110001111: color_data = Z;
		19'b0110100100110010000: color_data = Z;
		19'b0110100100110010001: color_data = Z;
		19'b0110100100110010010: color_data = Z;
		19'b0110100100110010011: color_data = Z;
		19'b0110100100110010100: color_data = Z;
		19'b0110100100110010101: color_data = Z;
		19'b0110100100111010001: color_data = Z;
		19'b0110100100111010010: color_data = Z;
		19'b0110100100111010011: color_data = Z;
		19'b0110100100111010100: color_data = Z;
		19'b0110100100111010101: color_data = Z;
		19'b0110100100111010110: color_data = Z;
		19'b0110100100111010111: color_data = Z;
		19'b0110100100111011000: color_data = Z;
		19'b0110100100111011001: color_data = Z;
		19'b0110100100111011010: color_data = Z;
		19'b0110100110010100011: color_data = Z;
		19'b0110100110010100100: color_data = Z;
		19'b0110100110010100101: color_data = Z;
		19'b0110100110010100110: color_data = Z;
		19'b0110100110010100111: color_data = Z;
		19'b0110100110010101000: color_data = Z;
		19'b0110100110010101001: color_data = Z;
		19'b0110100110100001101: color_data = Z;
		19'b0110100110100001110: color_data = Z;
		19'b0110100110100001111: color_data = Z;
		19'b0110100110100010000: color_data = Z;
		19'b0110100110100010001: color_data = Z;
		19'b0110100110100010010: color_data = Z;
		19'b0110100110100010011: color_data = Z;
		19'b0110100110100010100: color_data = Z;
		19'b0110100110100010101: color_data = Z;
		19'b0110100110100010110: color_data = Z;
		19'b0110100110100010111: color_data = Z;
		19'b0110100110100011000: color_data = Z;
		19'b0110100110100011001: color_data = Z;
		19'b0110100110100011011: color_data = Z;
		19'b0110100110100011100: color_data = Z;
		19'b0110100110100011101: color_data = Z;
		19'b0110100110100011110: color_data = Z;
		19'b0110100110100011111: color_data = Z;
		19'b0110100110100100000: color_data = Z;
		19'b0110100110100100001: color_data = Z;
		19'b0110100110100100010: color_data = Z;
		19'b0110100110100100011: color_data = Z;
		19'b0110100110100100100: color_data = Z;
		19'b0110100110100100101: color_data = Z;
		19'b0110100110100100110: color_data = Z;
		19'b0110100110100100111: color_data = Z;
		19'b0110100110100101000: color_data = Z;
		19'b0110100110100101001: color_data = Z;
		19'b0110100110100101010: color_data = Z;
		19'b0110100110100101011: color_data = Z;
		19'b0110100110100101100: color_data = Z;
		19'b0110100110100101101: color_data = Z;
		19'b0110100110100101110: color_data = Z;
		19'b0110100110100101111: color_data = Z;
		19'b0110100110100110000: color_data = Z;
		19'b0110100110100110001: color_data = Z;
		19'b0110100110100110010: color_data = Z;
		19'b0110100110100110011: color_data = Z;
		19'b0110100110100110100: color_data = Z;
		19'b0110100110100110101: color_data = Z;
		19'b0110100110100110110: color_data = Z;
		19'b0110100110100110111: color_data = Z;
		19'b0110100110100111000: color_data = Z;
		19'b0110100110100111001: color_data = Z;
		19'b0110100110100111010: color_data = Z;
		19'b0110100110100111011: color_data = Z;
		19'b0110100110100111100: color_data = Z;
		19'b0110100110100111101: color_data = Z;
		19'b0110100110100111110: color_data = Z;
		19'b0110100110100111111: color_data = Z;
		19'b0110100110101000000: color_data = Z;
		19'b0110100110101000001: color_data = Z;
		19'b0110100110101000010: color_data = Z;
		19'b0110100110101000011: color_data = Z;
		19'b0110100110101000100: color_data = Z;
		19'b0110100110101000101: color_data = Z;
		19'b0110100110101000110: color_data = Z;
		19'b0110100110101000111: color_data = Z;
		19'b0110100110101001000: color_data = Z;
		19'b0110100110101001001: color_data = Z;
		19'b0110100110101001010: color_data = Z;
		19'b0110100110101001011: color_data = Z;
		19'b0110100110101001100: color_data = Z;
		19'b0110100110101001101: color_data = Z;
		19'b0110100110101001110: color_data = Z;
		19'b0110100110101001111: color_data = Z;
		19'b0110100110101010000: color_data = Z;
		19'b0110100110101010001: color_data = Z;
		19'b0110100110101010010: color_data = Z;
		19'b0110100110101010011: color_data = Z;
		19'b0110100110101010100: color_data = Z;
		19'b0110100110101010101: color_data = Z;
		19'b0110100110101010110: color_data = Z;
		19'b0110100110101010111: color_data = Z;
		19'b0110100110101011000: color_data = Z;
		19'b0110100110101011001: color_data = Z;
		19'b0110100110101011010: color_data = Z;
		19'b0110100110101011011: color_data = Z;
		19'b0110100110101011100: color_data = Z;
		19'b0110100110101011101: color_data = Z;
		19'b0110100110101011110: color_data = Z;
		19'b0110100110101011111: color_data = Z;
		19'b0110100110101100000: color_data = Z;
		19'b0110100110101100001: color_data = Z;
		19'b0110100110101100010: color_data = Z;
		19'b0110100110101100011: color_data = Z;
		19'b0110100110101100100: color_data = Z;
		19'b0110100110101100101: color_data = Z;
		19'b0110100110101100110: color_data = Z;
		19'b0110100110101100111: color_data = Z;
		19'b0110100110101101011: color_data = Z;
		19'b0110100110101101100: color_data = Z;
		19'b0110100110101101101: color_data = Z;
		19'b0110100110101101110: color_data = Z;
		19'b0110100110101101111: color_data = Z;
		19'b0110100110101110000: color_data = Z;
		19'b0110100110101110001: color_data = Z;
		19'b0110100110101110010: color_data = Z;
		19'b0110100110101110011: color_data = Z;
		19'b0110100110101110100: color_data = Z;
		19'b0110100110101110101: color_data = Z;
		19'b0110100110101110110: color_data = Z;
		19'b0110100110101110111: color_data = Z;
		19'b0110100110101111000: color_data = Z;
		19'b0110100110101111001: color_data = Z;
		19'b0110100110101111010: color_data = Z;
		19'b0110100110101111110: color_data = Z;
		19'b0110100110101111111: color_data = Z;
		19'b0110100110110000000: color_data = Z;
		19'b0110100110110000001: color_data = Z;
		19'b0110100110110000010: color_data = Z;
		19'b0110100110110000011: color_data = Z;
		19'b0110100110110000100: color_data = Z;
		19'b0110100110110000101: color_data = Z;
		19'b0110100110110000110: color_data = Z;
		19'b0110100110110000111: color_data = Z;
		19'b0110100110110001000: color_data = Z;
		19'b0110100110110001001: color_data = Z;
		19'b0110100110110001010: color_data = Z;
		19'b0110100110110001011: color_data = Z;
		19'b0110100110110001100: color_data = Z;
		19'b0110100110110001101: color_data = Z;
		19'b0110100110110001110: color_data = Z;
		19'b0110100110110001111: color_data = Z;
		19'b0110100110110010000: color_data = Z;
		19'b0110100110110010001: color_data = Z;
		19'b0110100110110010010: color_data = Z;
		19'b0110100110111010001: color_data = Z;
		19'b0110100110111010010: color_data = Z;
		19'b0110100110111010011: color_data = Z;
		19'b0110100110111010100: color_data = Z;
		19'b0110100110111010101: color_data = Z;
		19'b0110100110111010110: color_data = Z;
		19'b0110100110111010111: color_data = Z;
		19'b0110100110111011000: color_data = Z;
		19'b0110100110111011001: color_data = Z;
		19'b0110100110111011010: color_data = Z;
		19'b0110101000010100011: color_data = Z;
		19'b0110101000010100100: color_data = Z;
		19'b0110101000010100101: color_data = Z;
		19'b0110101000010100110: color_data = Z;
		19'b0110101000010100111: color_data = Z;
		19'b0110101000010101000: color_data = Z;
		19'b0110101000010101001: color_data = Z;
		19'b0110101000100001101: color_data = Z;
		19'b0110101000100001110: color_data = Z;
		19'b0110101000100001111: color_data = Z;
		19'b0110101000100010000: color_data = Z;
		19'b0110101000100010001: color_data = Z;
		19'b0110101000100010010: color_data = Z;
		19'b0110101000100010011: color_data = Z;
		19'b0110101000100010100: color_data = Z;
		19'b0110101000100010101: color_data = Z;
		19'b0110101000100010110: color_data = Z;
		19'b0110101000100010111: color_data = Z;
		19'b0110101000100011000: color_data = Z;
		19'b0110101000100011001: color_data = Z;
		19'b0110101000100011011: color_data = Z;
		19'b0110101000100011100: color_data = Z;
		19'b0110101000100011101: color_data = Z;
		19'b0110101000100011110: color_data = Z;
		19'b0110101000100011111: color_data = Z;
		19'b0110101000100100000: color_data = Z;
		19'b0110101000100100001: color_data = Z;
		19'b0110101000100100010: color_data = Z;
		19'b0110101000100100011: color_data = Z;
		19'b0110101000100100100: color_data = Z;
		19'b0110101000100100101: color_data = Z;
		19'b0110101000100100110: color_data = Z;
		19'b0110101000100100111: color_data = Z;
		19'b0110101000100101000: color_data = Z;
		19'b0110101000100101001: color_data = Z;
		19'b0110101000100101010: color_data = Z;
		19'b0110101000100101011: color_data = Z;
		19'b0110101000100101100: color_data = Z;
		19'b0110101000100101101: color_data = Z;
		19'b0110101000100101110: color_data = Z;
		19'b0110101000100101111: color_data = Z;
		19'b0110101000100110000: color_data = Z;
		19'b0110101000100110001: color_data = Z;
		19'b0110101000100110010: color_data = Z;
		19'b0110101000100110011: color_data = Z;
		19'b0110101000100110100: color_data = Z;
		19'b0110101000100110101: color_data = Z;
		19'b0110101000100110110: color_data = Z;
		19'b0110101000100110111: color_data = Z;
		19'b0110101000100111000: color_data = Z;
		19'b0110101000100111001: color_data = Z;
		19'b0110101000100111010: color_data = Z;
		19'b0110101000100111011: color_data = Z;
		19'b0110101000100111100: color_data = Z;
		19'b0110101000100111101: color_data = Z;
		19'b0110101000100111110: color_data = Z;
		19'b0110101000100111111: color_data = Z;
		19'b0110101000101000000: color_data = Z;
		19'b0110101000101000001: color_data = Z;
		19'b0110101000101000010: color_data = Z;
		19'b0110101000101000011: color_data = Z;
		19'b0110101000101000100: color_data = Z;
		19'b0110101000101000101: color_data = Z;
		19'b0110101000101000110: color_data = Z;
		19'b0110101000101000111: color_data = Z;
		19'b0110101000101001000: color_data = Z;
		19'b0110101000101001001: color_data = Z;
		19'b0110101000101001010: color_data = Z;
		19'b0110101000101001011: color_data = Z;
		19'b0110101000101001100: color_data = Z;
		19'b0110101000101001101: color_data = Z;
		19'b0110101000101001110: color_data = Z;
		19'b0110101000101001111: color_data = Z;
		19'b0110101000101010000: color_data = Z;
		19'b0110101000101010001: color_data = Z;
		19'b0110101000101010010: color_data = Z;
		19'b0110101000101010011: color_data = Z;
		19'b0110101000101010100: color_data = Z;
		19'b0110101000101010101: color_data = Z;
		19'b0110101000101010110: color_data = Z;
		19'b0110101000101010111: color_data = Z;
		19'b0110101000101011000: color_data = Z;
		19'b0110101000101011001: color_data = Z;
		19'b0110101000101011010: color_data = Z;
		19'b0110101000101011011: color_data = Z;
		19'b0110101000101011100: color_data = Z;
		19'b0110101000101011101: color_data = Z;
		19'b0110101000101011110: color_data = Z;
		19'b0110101000101011111: color_data = Z;
		19'b0110101000101100000: color_data = Z;
		19'b0110101000101100001: color_data = Z;
		19'b0110101000101100010: color_data = Z;
		19'b0110101000101100011: color_data = Z;
		19'b0110101000101100100: color_data = Z;
		19'b0110101000101100101: color_data = Z;
		19'b0110101000101100110: color_data = Z;
		19'b0110101000101100111: color_data = Z;
		19'b0110101000101101000: color_data = Z;
		19'b0110101000101101011: color_data = Z;
		19'b0110101000101101100: color_data = Z;
		19'b0110101000101101101: color_data = Z;
		19'b0110101000101101110: color_data = Z;
		19'b0110101000101101111: color_data = Z;
		19'b0110101000101110000: color_data = Z;
		19'b0110101000101110001: color_data = Z;
		19'b0110101000101110010: color_data = Z;
		19'b0110101000101110011: color_data = Z;
		19'b0110101000101110100: color_data = Z;
		19'b0110101000101110101: color_data = Z;
		19'b0110101000101110110: color_data = Z;
		19'b0110101000101110111: color_data = Z;
		19'b0110101000101111000: color_data = Z;
		19'b0110101000101111001: color_data = Z;
		19'b0110101000101111010: color_data = Z;
		19'b0110101000101111111: color_data = Z;
		19'b0110101000110000000: color_data = Z;
		19'b0110101000110000001: color_data = Z;
		19'b0110101000110000010: color_data = Z;
		19'b0110101000110000011: color_data = Z;
		19'b0110101000110000100: color_data = Z;
		19'b0110101000110000101: color_data = Z;
		19'b0110101000110000110: color_data = Z;
		19'b0110101000110000111: color_data = Z;
		19'b0110101000110001000: color_data = Z;
		19'b0110101000110001001: color_data = Z;
		19'b0110101000110001010: color_data = Z;
		19'b0110101000110001011: color_data = Z;
		19'b0110101000110001100: color_data = Z;
		19'b0110101000110001101: color_data = Z;
		19'b0110101000110001110: color_data = Z;
		19'b0110101000110001111: color_data = Z;
		19'b0110101000110010000: color_data = Z;
		19'b0110101000110010001: color_data = Z;
		19'b0110101000111010001: color_data = Z;
		19'b0110101000111010010: color_data = Z;
		19'b0110101000111010011: color_data = Z;
		19'b0110101000111010100: color_data = Z;
		19'b0110101000111010101: color_data = Z;
		19'b0110101000111010110: color_data = Z;
		19'b0110101000111010111: color_data = Z;
		19'b0110101000111011000: color_data = Z;
		19'b0110101000111011001: color_data = Z;
		19'b0110101000111011010: color_data = Z;
		19'b0110101010010100011: color_data = Z;
		19'b0110101010010100100: color_data = Z;
		19'b0110101010010100101: color_data = Z;
		19'b0110101010010100110: color_data = Z;
		19'b0110101010010100111: color_data = Z;
		19'b0110101010010101000: color_data = Z;
		19'b0110101010010101001: color_data = Z;
		19'b0110101010100001100: color_data = Z;
		19'b0110101010100001101: color_data = Z;
		19'b0110101010100001110: color_data = Z;
		19'b0110101010100001111: color_data = Z;
		19'b0110101010100010000: color_data = Z;
		19'b0110101010100010001: color_data = Z;
		19'b0110101010100010010: color_data = Z;
		19'b0110101010100010011: color_data = Z;
		19'b0110101010100010100: color_data = Z;
		19'b0110101010100010101: color_data = Z;
		19'b0110101010100010110: color_data = Z;
		19'b0110101010100010111: color_data = Z;
		19'b0110101010100011000: color_data = Z;
		19'b0110101010100011001: color_data = Z;
		19'b0110101010100011010: color_data = Z;
		19'b0110101010100011011: color_data = Z;
		19'b0110101010100011100: color_data = Z;
		19'b0110101010100011101: color_data = Z;
		19'b0110101010100011110: color_data = Z;
		19'b0110101010100011111: color_data = Z;
		19'b0110101010100100000: color_data = Z;
		19'b0110101010100100001: color_data = Z;
		19'b0110101010100100010: color_data = Z;
		19'b0110101010100100011: color_data = Z;
		19'b0110101010100100100: color_data = Z;
		19'b0110101010100100101: color_data = Z;
		19'b0110101010100100110: color_data = Z;
		19'b0110101010100100111: color_data = Z;
		19'b0110101010100101000: color_data = Z;
		19'b0110101010100101001: color_data = Z;
		19'b0110101010100101010: color_data = Z;
		19'b0110101010100101011: color_data = Z;
		19'b0110101010100101100: color_data = Z;
		19'b0110101010100101101: color_data = Z;
		19'b0110101010100101111: color_data = Z;
		19'b0110101010100110000: color_data = Z;
		19'b0110101010100110001: color_data = Z;
		19'b0110101010100110010: color_data = Z;
		19'b0110101010100110011: color_data = Z;
		19'b0110101010100110100: color_data = Z;
		19'b0110101010100110101: color_data = Z;
		19'b0110101010100110110: color_data = Z;
		19'b0110101010100110111: color_data = Z;
		19'b0110101010100111000: color_data = Z;
		19'b0110101010100111001: color_data = Z;
		19'b0110101010100111010: color_data = Z;
		19'b0110101010100111011: color_data = Z;
		19'b0110101010100111100: color_data = Z;
		19'b0110101010100111101: color_data = Z;
		19'b0110101010100111110: color_data = Z;
		19'b0110101010100111111: color_data = Z;
		19'b0110101010101000000: color_data = Z;
		19'b0110101010101000001: color_data = Z;
		19'b0110101010101000010: color_data = Z;
		19'b0110101010101000011: color_data = Z;
		19'b0110101010101000100: color_data = Z;
		19'b0110101010101000101: color_data = Z;
		19'b0110101010101000110: color_data = Z;
		19'b0110101010101000111: color_data = Z;
		19'b0110101010101001000: color_data = Z;
		19'b0110101010101001001: color_data = Z;
		19'b0110101010101001010: color_data = Z;
		19'b0110101010101001011: color_data = Z;
		19'b0110101010101001100: color_data = Z;
		19'b0110101010101001101: color_data = Z;
		19'b0110101010101001110: color_data = Z;
		19'b0110101010101001111: color_data = Z;
		19'b0110101010101010000: color_data = Z;
		19'b0110101010101010001: color_data = Z;
		19'b0110101010101010010: color_data = Z;
		19'b0110101010101010011: color_data = Z;
		19'b0110101010101010100: color_data = Z;
		19'b0110101010101010101: color_data = Z;
		19'b0110101010101010110: color_data = Z;
		19'b0110101010101010111: color_data = Z;
		19'b0110101010101011000: color_data = Z;
		19'b0110101010101011001: color_data = Z;
		19'b0110101010101011010: color_data = Z;
		19'b0110101010101011011: color_data = Z;
		19'b0110101010101011100: color_data = Z;
		19'b0110101010101011101: color_data = Z;
		19'b0110101010101011110: color_data = Z;
		19'b0110101010101011111: color_data = Z;
		19'b0110101010101100000: color_data = Z;
		19'b0110101010101100001: color_data = Z;
		19'b0110101010101100010: color_data = Z;
		19'b0110101010101100011: color_data = Z;
		19'b0110101010101100100: color_data = Z;
		19'b0110101010101100101: color_data = Z;
		19'b0110101010101100110: color_data = Z;
		19'b0110101010101100111: color_data = Z;
		19'b0110101010101101000: color_data = Z;
		19'b0110101010101101100: color_data = Z;
		19'b0110101010101101101: color_data = Z;
		19'b0110101010101101110: color_data = Z;
		19'b0110101010101101111: color_data = Z;
		19'b0110101010101110000: color_data = Z;
		19'b0110101010101110001: color_data = Z;
		19'b0110101010101110010: color_data = Z;
		19'b0110101010101110011: color_data = Z;
		19'b0110101010101110100: color_data = Z;
		19'b0110101010101110101: color_data = Z;
		19'b0110101010101110110: color_data = Z;
		19'b0110101010101110111: color_data = Z;
		19'b0110101010101111000: color_data = Z;
		19'b0110101010101111001: color_data = Z;
		19'b0110101010101111010: color_data = Z;
		19'b0110101010101111111: color_data = Z;
		19'b0110101010110000000: color_data = Z;
		19'b0110101010110000001: color_data = Z;
		19'b0110101010110000010: color_data = Z;
		19'b0110101010110000011: color_data = Z;
		19'b0110101010110000100: color_data = Z;
		19'b0110101010110000101: color_data = Z;
		19'b0110101010110000110: color_data = Z;
		19'b0110101010110000111: color_data = Z;
		19'b0110101010110001000: color_data = Z;
		19'b0110101010110001001: color_data = Z;
		19'b0110101010110001010: color_data = Z;
		19'b0110101010110001011: color_data = Z;
		19'b0110101010110001100: color_data = Z;
		19'b0110101010110001101: color_data = Z;
		19'b0110101010110001110: color_data = Z;
		19'b0110101010110001111: color_data = Z;
		19'b0110101010110010000: color_data = Z;
		19'b0110101010110010001: color_data = Z;
		19'b0110101010111010010: color_data = Z;
		19'b0110101010111010011: color_data = Z;
		19'b0110101010111010100: color_data = Z;
		19'b0110101010111010101: color_data = Z;
		19'b0110101010111010110: color_data = Z;
		19'b0110101010111010111: color_data = Z;
		19'b0110101010111011000: color_data = Z;
		19'b0110101010111011001: color_data = Z;
		19'b0110101010111011010: color_data = Z;
		19'b0110101100010100100: color_data = Z;
		19'b0110101100010100101: color_data = Z;
		19'b0110101100010100110: color_data = Z;
		19'b0110101100010100111: color_data = Z;
		19'b0110101100010101000: color_data = Z;
		19'b0110101100010101001: color_data = Z;
		19'b0110101100010101010: color_data = Z;
		19'b0110101100010110001: color_data = Z;
		19'b0110101100010110010: color_data = Z;
		19'b0110101100100001100: color_data = Z;
		19'b0110101100100001101: color_data = Z;
		19'b0110101100100001110: color_data = Z;
		19'b0110101100100001111: color_data = Z;
		19'b0110101100100010000: color_data = Z;
		19'b0110101100100010001: color_data = Z;
		19'b0110101100100010010: color_data = Z;
		19'b0110101100100010011: color_data = Z;
		19'b0110101100100010100: color_data = Z;
		19'b0110101100100010101: color_data = Z;
		19'b0110101100100010110: color_data = Z;
		19'b0110101100100010111: color_data = Z;
		19'b0110101100100011010: color_data = Z;
		19'b0110101100100011011: color_data = Z;
		19'b0110101100100011100: color_data = Z;
		19'b0110101100100011101: color_data = Z;
		19'b0110101100100011110: color_data = Z;
		19'b0110101100100011111: color_data = Z;
		19'b0110101100100100000: color_data = Z;
		19'b0110101100100100001: color_data = Z;
		19'b0110101100100100010: color_data = Z;
		19'b0110101100100100011: color_data = Z;
		19'b0110101100100100100: color_data = Z;
		19'b0110101100100100101: color_data = Z;
		19'b0110101100100100110: color_data = Z;
		19'b0110101100100100111: color_data = Z;
		19'b0110101100100101000: color_data = Z;
		19'b0110101100100101001: color_data = Z;
		19'b0110101100100101010: color_data = Z;
		19'b0110101100100101011: color_data = Z;
		19'b0110101100100101100: color_data = Z;
		19'b0110101100100101111: color_data = Z;
		19'b0110101100100110000: color_data = Z;
		19'b0110101100100110001: color_data = Z;
		19'b0110101100100110010: color_data = Z;
		19'b0110101100100110011: color_data = Z;
		19'b0110101100100110100: color_data = Z;
		19'b0110101100100110101: color_data = Z;
		19'b0110101100100110110: color_data = Z;
		19'b0110101100100110111: color_data = Z;
		19'b0110101100100111000: color_data = Z;
		19'b0110101100100111001: color_data = Z;
		19'b0110101100100111010: color_data = Z;
		19'b0110101100100111011: color_data = Z;
		19'b0110101100100111100: color_data = Z;
		19'b0110101100100111101: color_data = Z;
		19'b0110101100100111110: color_data = Z;
		19'b0110101100100111111: color_data = Z;
		19'b0110101100101000000: color_data = Z;
		19'b0110101100101000001: color_data = Z;
		19'b0110101100101000010: color_data = Z;
		19'b0110101100101000011: color_data = Z;
		19'b0110101100101000100: color_data = Z;
		19'b0110101100101000101: color_data = Z;
		19'b0110101100101000110: color_data = Z;
		19'b0110101100101000111: color_data = Z;
		19'b0110101100101001000: color_data = Z;
		19'b0110101100101001001: color_data = Z;
		19'b0110101100101001010: color_data = Z;
		19'b0110101100101001011: color_data = Z;
		19'b0110101100101001100: color_data = Z;
		19'b0110101100101001101: color_data = Z;
		19'b0110101100101001110: color_data = Z;
		19'b0110101100101001111: color_data = Z;
		19'b0110101100101010000: color_data = Z;
		19'b0110101100101010001: color_data = Z;
		19'b0110101100101010010: color_data = Z;
		19'b0110101100101010011: color_data = Z;
		19'b0110101100101010100: color_data = Z;
		19'b0110101100101010101: color_data = Z;
		19'b0110101100101010110: color_data = Z;
		19'b0110101100101010111: color_data = Z;
		19'b0110101100101011000: color_data = Z;
		19'b0110101100101011001: color_data = Z;
		19'b0110101100101011010: color_data = Z;
		19'b0110101100101011011: color_data = Z;
		19'b0110101100101011100: color_data = Z;
		19'b0110101100101011101: color_data = Z;
		19'b0110101100101011110: color_data = Z;
		19'b0110101100101011111: color_data = Z;
		19'b0110101100101100000: color_data = Z;
		19'b0110101100101100001: color_data = Z;
		19'b0110101100101100010: color_data = Z;
		19'b0110101100101100011: color_data = Z;
		19'b0110101100101100100: color_data = Z;
		19'b0110101100101100101: color_data = Z;
		19'b0110101100101100110: color_data = Z;
		19'b0110101100101100111: color_data = Z;
		19'b0110101100101101000: color_data = Z;
		19'b0110101100101101101: color_data = Z;
		19'b0110101100101101110: color_data = Z;
		19'b0110101100101101111: color_data = Z;
		19'b0110101100101110000: color_data = Z;
		19'b0110101100101110001: color_data = Z;
		19'b0110101100101110010: color_data = Z;
		19'b0110101100101110011: color_data = Z;
		19'b0110101100101110100: color_data = Z;
		19'b0110101100101110101: color_data = Z;
		19'b0110101100101110110: color_data = Z;
		19'b0110101100101110111: color_data = Z;
		19'b0110101100101111000: color_data = Z;
		19'b0110101100101111001: color_data = Z;
		19'b0110101100101111010: color_data = Z;
		19'b0110101100110000000: color_data = Z;
		19'b0110101100110000001: color_data = Z;
		19'b0110101100110000010: color_data = Z;
		19'b0110101100110000011: color_data = Z;
		19'b0110101100110000100: color_data = Z;
		19'b0110101100110000101: color_data = Z;
		19'b0110101100110000110: color_data = Z;
		19'b0110101100110000111: color_data = Z;
		19'b0110101100110001000: color_data = Z;
		19'b0110101100110001001: color_data = Z;
		19'b0110101100110001010: color_data = Z;
		19'b0110101100110001011: color_data = Z;
		19'b0110101100110001100: color_data = Z;
		19'b0110101100110001101: color_data = Z;
		19'b0110101100110001110: color_data = Z;
		19'b0110101100110001111: color_data = Z;
		19'b0110101100110010000: color_data = Z;
		19'b0110101100110010001: color_data = Z;
		19'b0110101100110010010: color_data = Z;
		19'b0110101100111010010: color_data = Z;
		19'b0110101100111010011: color_data = Z;
		19'b0110101100111010100: color_data = Z;
		19'b0110101100111010101: color_data = Z;
		19'b0110101100111010110: color_data = Z;
		19'b0110101100111010111: color_data = Z;
		19'b0110101100111011000: color_data = Z;
		19'b0110101100111011001: color_data = Z;
		19'b0110101110010100100: color_data = Z;
		19'b0110101110010100101: color_data = Z;
		19'b0110101110010100110: color_data = Z;
		19'b0110101110010100111: color_data = Z;
		19'b0110101110010101000: color_data = Z;
		19'b0110101110010101001: color_data = Z;
		19'b0110101110010101010: color_data = Z;
		19'b0110101110010110010: color_data = Z;
		19'b0110101110010110011: color_data = Z;
		19'b0110101110100001100: color_data = Z;
		19'b0110101110100001101: color_data = Z;
		19'b0110101110100001110: color_data = Z;
		19'b0110101110100001111: color_data = Z;
		19'b0110101110100010000: color_data = Z;
		19'b0110101110100010001: color_data = Z;
		19'b0110101110100010010: color_data = Z;
		19'b0110101110100010011: color_data = Z;
		19'b0110101110100010100: color_data = Z;
		19'b0110101110100010101: color_data = Z;
		19'b0110101110100010110: color_data = Z;
		19'b0110101110100011001: color_data = Z;
		19'b0110101110100011010: color_data = Z;
		19'b0110101110100011011: color_data = Z;
		19'b0110101110100011100: color_data = Z;
		19'b0110101110100011101: color_data = Z;
		19'b0110101110100011110: color_data = Z;
		19'b0110101110100011111: color_data = Z;
		19'b0110101110100100000: color_data = Z;
		19'b0110101110100100001: color_data = Z;
		19'b0110101110100100010: color_data = Z;
		19'b0110101110100100011: color_data = Z;
		19'b0110101110100100100: color_data = Z;
		19'b0110101110100100101: color_data = Z;
		19'b0110101110100100110: color_data = Z;
		19'b0110101110100100111: color_data = Z;
		19'b0110101110100101000: color_data = Z;
		19'b0110101110100101001: color_data = Z;
		19'b0110101110100101010: color_data = Z;
		19'b0110101110100101011: color_data = Z;
		19'b0110101110100101100: color_data = Z;
		19'b0110101110100101111: color_data = Z;
		19'b0110101110100110000: color_data = Z;
		19'b0110101110100110001: color_data = Z;
		19'b0110101110100110010: color_data = Z;
		19'b0110101110100110011: color_data = Z;
		19'b0110101110100110100: color_data = Z;
		19'b0110101110100110101: color_data = Z;
		19'b0110101110100110110: color_data = Z;
		19'b0110101110100110111: color_data = Z;
		19'b0110101110100111000: color_data = Z;
		19'b0110101110100111001: color_data = Z;
		19'b0110101110100111010: color_data = Z;
		19'b0110101110100111011: color_data = Z;
		19'b0110101110100111100: color_data = Z;
		19'b0110101110100111101: color_data = Z;
		19'b0110101110100111110: color_data = Z;
		19'b0110101110100111111: color_data = Z;
		19'b0110101110101000000: color_data = Z;
		19'b0110101110101000001: color_data = Z;
		19'b0110101110101000010: color_data = Z;
		19'b0110101110101000011: color_data = Z;
		19'b0110101110101000100: color_data = Z;
		19'b0110101110101000101: color_data = Z;
		19'b0110101110101000110: color_data = Z;
		19'b0110101110101000111: color_data = Z;
		19'b0110101110101001000: color_data = Z;
		19'b0110101110101001001: color_data = Z;
		19'b0110101110101001010: color_data = Z;
		19'b0110101110101001011: color_data = Z;
		19'b0110101110101001100: color_data = Z;
		19'b0110101110101001101: color_data = Z;
		19'b0110101110101001110: color_data = Z;
		19'b0110101110101001111: color_data = Z;
		19'b0110101110101010000: color_data = Z;
		19'b0110101110101010001: color_data = Z;
		19'b0110101110101010010: color_data = Z;
		19'b0110101110101010011: color_data = Z;
		19'b0110101110101010100: color_data = Z;
		19'b0110101110101010101: color_data = Z;
		19'b0110101110101010110: color_data = Z;
		19'b0110101110101010111: color_data = Z;
		19'b0110101110101011000: color_data = Z;
		19'b0110101110101011001: color_data = Z;
		19'b0110101110101011010: color_data = Z;
		19'b0110101110101011011: color_data = Z;
		19'b0110101110101011100: color_data = Z;
		19'b0110101110101011101: color_data = Z;
		19'b0110101110101011110: color_data = Z;
		19'b0110101110101011111: color_data = Z;
		19'b0110101110101100000: color_data = Z;
		19'b0110101110101100001: color_data = Z;
		19'b0110101110101100010: color_data = Z;
		19'b0110101110101100011: color_data = Z;
		19'b0110101110101100100: color_data = Z;
		19'b0110101110101100101: color_data = Z;
		19'b0110101110101100110: color_data = Z;
		19'b0110101110101100111: color_data = Z;
		19'b0110101110101101000: color_data = Z;
		19'b0110101110101101101: color_data = Z;
		19'b0110101110101101110: color_data = Z;
		19'b0110101110101101111: color_data = Z;
		19'b0110101110101110000: color_data = Z;
		19'b0110101110101110001: color_data = Z;
		19'b0110101110101110010: color_data = Z;
		19'b0110101110101110011: color_data = Z;
		19'b0110101110101110100: color_data = Z;
		19'b0110101110101110101: color_data = Z;
		19'b0110101110101110110: color_data = Z;
		19'b0110101110101110111: color_data = Z;
		19'b0110101110101111000: color_data = Z;
		19'b0110101110101111001: color_data = Z;
		19'b0110101110101111010: color_data = Z;
		19'b0110101110110000000: color_data = Z;
		19'b0110101110110000001: color_data = Z;
		19'b0110101110110000010: color_data = Z;
		19'b0110101110110000011: color_data = Z;
		19'b0110101110110000100: color_data = Z;
		19'b0110101110110000101: color_data = Z;
		19'b0110101110110000110: color_data = Z;
		19'b0110101110110000111: color_data = Z;
		19'b0110101110110001000: color_data = Z;
		19'b0110101110110001001: color_data = Z;
		19'b0110101110110001010: color_data = Z;
		19'b0110101110110001011: color_data = Z;
		19'b0110101110110001100: color_data = Z;
		19'b0110101110110001101: color_data = Z;
		19'b0110101110110001110: color_data = Z;
		19'b0110101110110001111: color_data = Z;
		19'b0110101110110010000: color_data = Z;
		19'b0110101110110010001: color_data = Z;
		19'b0110101110110010010: color_data = Z;
		19'b0110101110110010011: color_data = Z;
		19'b0110101110111010001: color_data = Z;
		19'b0110101110111010010: color_data = Z;
		19'b0110101110111010011: color_data = Z;
		19'b0110101110111010100: color_data = Z;
		19'b0110101110111010101: color_data = Z;
		19'b0110101110111010110: color_data = Z;
		19'b0110101110111010111: color_data = Z;
		19'b0110101110111011000: color_data = Z;
		19'b0110101110111011001: color_data = Z;
		19'b0110110000010100101: color_data = Z;
		19'b0110110000010100110: color_data = Z;
		19'b0110110000010100111: color_data = Z;
		19'b0110110000010101000: color_data = Z;
		19'b0110110000010101001: color_data = Z;
		19'b0110110000010101010: color_data = Z;
		19'b0110110000010110010: color_data = Z;
		19'b0110110000010110011: color_data = Z;
		19'b0110110000010110100: color_data = Z;
		19'b0110110000100001101: color_data = Z;
		19'b0110110000100001110: color_data = Z;
		19'b0110110000100001111: color_data = Z;
		19'b0110110000100010000: color_data = Z;
		19'b0110110000100010001: color_data = Z;
		19'b0110110000100010010: color_data = Z;
		19'b0110110000100010011: color_data = Z;
		19'b0110110000100010100: color_data = Z;
		19'b0110110000100010101: color_data = Z;
		19'b0110110000100011001: color_data = Z;
		19'b0110110000100011010: color_data = Z;
		19'b0110110000100011011: color_data = Z;
		19'b0110110000100011100: color_data = Z;
		19'b0110110000100011101: color_data = Z;
		19'b0110110000100011110: color_data = Z;
		19'b0110110000100011111: color_data = Z;
		19'b0110110000100100000: color_data = Z;
		19'b0110110000100100001: color_data = Z;
		19'b0110110000100100010: color_data = Z;
		19'b0110110000100100011: color_data = Z;
		19'b0110110000100100100: color_data = Z;
		19'b0110110000100100101: color_data = Z;
		19'b0110110000100100110: color_data = Z;
		19'b0110110000100100111: color_data = Z;
		19'b0110110000100101000: color_data = Z;
		19'b0110110000100101001: color_data = Z;
		19'b0110110000100101010: color_data = Z;
		19'b0110110000100101011: color_data = Z;
		19'b0110110000100101100: color_data = Z;
		19'b0110110000100101110: color_data = Z;
		19'b0110110000100101111: color_data = Z;
		19'b0110110000100110000: color_data = Z;
		19'b0110110000100110001: color_data = Z;
		19'b0110110000100110010: color_data = Z;
		19'b0110110000100110011: color_data = Z;
		19'b0110110000100110100: color_data = Z;
		19'b0110110000100110101: color_data = Z;
		19'b0110110000100110110: color_data = Z;
		19'b0110110000100110111: color_data = Z;
		19'b0110110000100111000: color_data = Z;
		19'b0110110000100111001: color_data = Z;
		19'b0110110000100111010: color_data = Z;
		19'b0110110000100111011: color_data = Z;
		19'b0110110000100111100: color_data = Z;
		19'b0110110000100111101: color_data = Z;
		19'b0110110000100111110: color_data = Z;
		19'b0110110000100111111: color_data = Z;
		19'b0110110000101000000: color_data = Z;
		19'b0110110000101000001: color_data = Z;
		19'b0110110000101000010: color_data = Z;
		19'b0110110000101000011: color_data = Z;
		19'b0110110000101000100: color_data = Z;
		19'b0110110000101000101: color_data = Z;
		19'b0110110000101000110: color_data = Z;
		19'b0110110000101000111: color_data = Z;
		19'b0110110000101001000: color_data = Z;
		19'b0110110000101001001: color_data = Z;
		19'b0110110000101001010: color_data = Z;
		19'b0110110000101001011: color_data = Z;
		19'b0110110000101001100: color_data = Z;
		19'b0110110000101001101: color_data = Z;
		19'b0110110000101001110: color_data = Z;
		19'b0110110000101001111: color_data = Z;
		19'b0110110000101010000: color_data = Z;
		19'b0110110000101010001: color_data = Z;
		19'b0110110000101010010: color_data = Z;
		19'b0110110000101010011: color_data = Z;
		19'b0110110000101010100: color_data = Z;
		19'b0110110000101010101: color_data = Z;
		19'b0110110000101010110: color_data = Z;
		19'b0110110000101010111: color_data = Z;
		19'b0110110000101011000: color_data = Z;
		19'b0110110000101011001: color_data = Z;
		19'b0110110000101011010: color_data = Z;
		19'b0110110000101011011: color_data = Z;
		19'b0110110000101011100: color_data = Z;
		19'b0110110000101011101: color_data = Z;
		19'b0110110000101011110: color_data = Z;
		19'b0110110000101011111: color_data = Z;
		19'b0110110000101100000: color_data = Z;
		19'b0110110000101100001: color_data = Z;
		19'b0110110000101100010: color_data = Z;
		19'b0110110000101100011: color_data = Z;
		19'b0110110000101100100: color_data = Z;
		19'b0110110000101100101: color_data = Z;
		19'b0110110000101100110: color_data = Z;
		19'b0110110000101100111: color_data = Z;
		19'b0110110000101101000: color_data = Z;
		19'b0110110000101101110: color_data = Z;
		19'b0110110000101101111: color_data = Z;
		19'b0110110000101110000: color_data = Z;
		19'b0110110000101110001: color_data = Z;
		19'b0110110000101110010: color_data = Z;
		19'b0110110000101110011: color_data = Z;
		19'b0110110000101110100: color_data = Z;
		19'b0110110000101110101: color_data = Z;
		19'b0110110000101110110: color_data = Z;
		19'b0110110000101110111: color_data = Z;
		19'b0110110000101111000: color_data = Z;
		19'b0110110000101111001: color_data = Z;
		19'b0110110000101111010: color_data = Z;
		19'b0110110000101111011: color_data = Z;
		19'b0110110000110000001: color_data = Z;
		19'b0110110000110000010: color_data = Z;
		19'b0110110000110000011: color_data = Z;
		19'b0110110000110000100: color_data = Z;
		19'b0110110000110000101: color_data = Z;
		19'b0110110000110000110: color_data = Z;
		19'b0110110000110000111: color_data = Z;
		19'b0110110000110001000: color_data = Z;
		19'b0110110000110001001: color_data = Z;
		19'b0110110000110001010: color_data = Z;
		19'b0110110000110001011: color_data = Z;
		19'b0110110000110001100: color_data = Z;
		19'b0110110000110001101: color_data = Z;
		19'b0110110000110001110: color_data = Z;
		19'b0110110000110001111: color_data = Z;
		19'b0110110000110010000: color_data = Z;
		19'b0110110000110010001: color_data = Z;
		19'b0110110000110010010: color_data = Z;
		19'b0110110000111010000: color_data = Z;
		19'b0110110000111010001: color_data = Z;
		19'b0110110000111010010: color_data = Z;
		19'b0110110000111010011: color_data = Z;
		19'b0110110000111010100: color_data = Z;
		19'b0110110000111010101: color_data = Z;
		19'b0110110000111010110: color_data = Z;
		19'b0110110000111010111: color_data = Z;
		19'b0110110000111011000: color_data = Z;
		19'b0110110000111011001: color_data = Z;
		19'b0110110010010100101: color_data = Z;
		19'b0110110010010100110: color_data = Z;
		19'b0110110010010100111: color_data = Z;
		19'b0110110010010101000: color_data = Z;
		19'b0110110010010101001: color_data = Z;
		19'b0110110010010101010: color_data = Z;
		19'b0110110010010101011: color_data = Z;
		19'b0110110010010110011: color_data = Z;
		19'b0110110010010110100: color_data = Z;
		19'b0110110010100001101: color_data = Z;
		19'b0110110010100001110: color_data = Z;
		19'b0110110010100001111: color_data = Z;
		19'b0110110010100010000: color_data = Z;
		19'b0110110010100010001: color_data = Z;
		19'b0110110010100010010: color_data = Z;
		19'b0110110010100010011: color_data = Z;
		19'b0110110010100011001: color_data = Z;
		19'b0110110010100011010: color_data = Z;
		19'b0110110010100011011: color_data = Z;
		19'b0110110010100011100: color_data = Z;
		19'b0110110010100011101: color_data = Z;
		19'b0110110010100011110: color_data = Z;
		19'b0110110010100011111: color_data = Z;
		19'b0110110010100100000: color_data = Z;
		19'b0110110010100100001: color_data = Z;
		19'b0110110010100100010: color_data = Z;
		19'b0110110010100100011: color_data = Z;
		19'b0110110010100100100: color_data = Z;
		19'b0110110010100100101: color_data = Z;
		19'b0110110010100100110: color_data = Z;
		19'b0110110010100100111: color_data = Z;
		19'b0110110010100101000: color_data = Z;
		19'b0110110010100101001: color_data = Z;
		19'b0110110010100101010: color_data = Z;
		19'b0110110010100101011: color_data = Z;
		19'b0110110010100101100: color_data = Z;
		19'b0110110010100101110: color_data = Z;
		19'b0110110010100101111: color_data = Z;
		19'b0110110010100110000: color_data = Z;
		19'b0110110010100110001: color_data = Z;
		19'b0110110010100110010: color_data = Z;
		19'b0110110010100110011: color_data = Z;
		19'b0110110010100110100: color_data = Z;
		19'b0110110010100110101: color_data = Z;
		19'b0110110010100110110: color_data = Z;
		19'b0110110010100110111: color_data = Z;
		19'b0110110010100111000: color_data = Z;
		19'b0110110010100111001: color_data = Z;
		19'b0110110010100111010: color_data = Z;
		19'b0110110010100111011: color_data = Z;
		19'b0110110010100111100: color_data = Z;
		19'b0110110010100111101: color_data = Z;
		19'b0110110010100111110: color_data = Z;
		19'b0110110010100111111: color_data = Z;
		19'b0110110010101000000: color_data = Z;
		19'b0110110010101000001: color_data = Z;
		19'b0110110010101000010: color_data = Z;
		19'b0110110010101000011: color_data = Z;
		19'b0110110010101000100: color_data = Z;
		19'b0110110010101000101: color_data = Z;
		19'b0110110010101000110: color_data = Z;
		19'b0110110010101000111: color_data = Z;
		19'b0110110010101001000: color_data = Z;
		19'b0110110010101001001: color_data = Z;
		19'b0110110010101001010: color_data = Z;
		19'b0110110010101001011: color_data = Z;
		19'b0110110010101001100: color_data = Z;
		19'b0110110010101001101: color_data = Z;
		19'b0110110010101001110: color_data = Z;
		19'b0110110010101001111: color_data = Z;
		19'b0110110010101010000: color_data = Z;
		19'b0110110010101010001: color_data = Z;
		19'b0110110010101010010: color_data = Z;
		19'b0110110010101010011: color_data = Z;
		19'b0110110010101010100: color_data = Z;
		19'b0110110010101010101: color_data = Z;
		19'b0110110010101010110: color_data = Z;
		19'b0110110010101010111: color_data = Z;
		19'b0110110010101011000: color_data = Z;
		19'b0110110010101011001: color_data = Z;
		19'b0110110010101011010: color_data = Z;
		19'b0110110010101011011: color_data = Z;
		19'b0110110010101011100: color_data = Z;
		19'b0110110010101011101: color_data = Z;
		19'b0110110010101011110: color_data = Z;
		19'b0110110010101011111: color_data = Z;
		19'b0110110010101100000: color_data = Z;
		19'b0110110010101100001: color_data = Z;
		19'b0110110010101100010: color_data = Z;
		19'b0110110010101100011: color_data = Z;
		19'b0110110010101100100: color_data = Z;
		19'b0110110010101100101: color_data = Z;
		19'b0110110010101100110: color_data = Z;
		19'b0110110010101100111: color_data = Z;
		19'b0110110010101101000: color_data = Z;
		19'b0110110010101101101: color_data = Z;
		19'b0110110010101101110: color_data = Z;
		19'b0110110010101101111: color_data = Z;
		19'b0110110010101110000: color_data = Z;
		19'b0110110010101110001: color_data = Z;
		19'b0110110010101110010: color_data = Z;
		19'b0110110010101110011: color_data = Z;
		19'b0110110010101110100: color_data = Z;
		19'b0110110010101110101: color_data = Z;
		19'b0110110010101110110: color_data = Z;
		19'b0110110010101110111: color_data = Z;
		19'b0110110010101111000: color_data = Z;
		19'b0110110010101111001: color_data = Z;
		19'b0110110010101111010: color_data = Z;
		19'b0110110010101111011: color_data = Z;
		19'b0110110010110000001: color_data = Z;
		19'b0110110010110000010: color_data = Z;
		19'b0110110010110000011: color_data = Z;
		19'b0110110010110000100: color_data = Z;
		19'b0110110010110000101: color_data = Z;
		19'b0110110010110000110: color_data = Z;
		19'b0110110010110000111: color_data = Z;
		19'b0110110010110001000: color_data = Z;
		19'b0110110010110001001: color_data = Z;
		19'b0110110010110001010: color_data = Z;
		19'b0110110010110001011: color_data = Z;
		19'b0110110010110001100: color_data = Z;
		19'b0110110010110001101: color_data = Z;
		19'b0110110010110001110: color_data = Z;
		19'b0110110010110001111: color_data = Z;
		19'b0110110010110010000: color_data = Z;
		19'b0110110010110010001: color_data = Z;
		19'b0110110010110010010: color_data = Z;
		19'b0110110010110010011: color_data = Z;
		19'b0110110010111010000: color_data = Z;
		19'b0110110010111010001: color_data = Z;
		19'b0110110010111010010: color_data = Z;
		19'b0110110010111010011: color_data = Z;
		19'b0110110010111010100: color_data = Z;
		19'b0110110010111010101: color_data = Z;
		19'b0110110010111010110: color_data = Z;
		19'b0110110010111010111: color_data = Z;
		19'b0110110010111011000: color_data = Z;
		19'b0110110100010100110: color_data = Z;
		19'b0110110100010100111: color_data = Z;
		19'b0110110100010101000: color_data = Z;
		19'b0110110100010101001: color_data = Z;
		19'b0110110100010101010: color_data = Z;
		19'b0110110100010101011: color_data = Z;
		19'b0110110100010110011: color_data = Z;
		19'b0110110100010110100: color_data = Z;
		19'b0110110100100001110: color_data = Z;
		19'b0110110100100001111: color_data = Z;
		19'b0110110100100010000: color_data = Z;
		19'b0110110100100010001: color_data = Z;
		19'b0110110100100010010: color_data = Z;
		19'b0110110100100011001: color_data = Z;
		19'b0110110100100011010: color_data = Z;
		19'b0110110100100011011: color_data = Z;
		19'b0110110100100011100: color_data = Z;
		19'b0110110100100011101: color_data = Z;
		19'b0110110100100011110: color_data = Z;
		19'b0110110100100011111: color_data = Z;
		19'b0110110100100100000: color_data = Z;
		19'b0110110100100100001: color_data = Z;
		19'b0110110100100100010: color_data = Z;
		19'b0110110100100100011: color_data = Z;
		19'b0110110100100100100: color_data = Z;
		19'b0110110100100100101: color_data = Z;
		19'b0110110100100100110: color_data = Z;
		19'b0110110100100100111: color_data = Z;
		19'b0110110100100101000: color_data = Z;
		19'b0110110100100101001: color_data = Z;
		19'b0110110100100101010: color_data = Z;
		19'b0110110100100101011: color_data = Z;
		19'b0110110100100101100: color_data = Z;
		19'b0110110100100101110: color_data = Z;
		19'b0110110100100101111: color_data = Z;
		19'b0110110100100110000: color_data = Z;
		19'b0110110100100110001: color_data = Z;
		19'b0110110100100110010: color_data = Z;
		19'b0110110100100110011: color_data = Z;
		19'b0110110100100110100: color_data = Z;
		19'b0110110100100110101: color_data = Z;
		19'b0110110100100110110: color_data = Z;
		19'b0110110100100110111: color_data = Z;
		19'b0110110100100111000: color_data = Z;
		19'b0110110100100111001: color_data = Z;
		19'b0110110100100111010: color_data = Z;
		19'b0110110100100111011: color_data = Z;
		19'b0110110100100111100: color_data = Z;
		19'b0110110100100111101: color_data = Z;
		19'b0110110100100111110: color_data = Z;
		19'b0110110100100111111: color_data = Z;
		19'b0110110100101000000: color_data = Z;
		19'b0110110100101000001: color_data = Z;
		19'b0110110100101000010: color_data = Z;
		19'b0110110100101000011: color_data = Z;
		19'b0110110100101000100: color_data = Z;
		19'b0110110100101000101: color_data = Z;
		19'b0110110100101000110: color_data = Z;
		19'b0110110100101000111: color_data = Z;
		19'b0110110100101001000: color_data = Z;
		19'b0110110100101001001: color_data = Z;
		19'b0110110100101001010: color_data = Z;
		19'b0110110100101001011: color_data = Z;
		19'b0110110100101001100: color_data = Z;
		19'b0110110100101001101: color_data = Z;
		19'b0110110100101001110: color_data = Z;
		19'b0110110100101001111: color_data = Z;
		19'b0110110100101010000: color_data = Z;
		19'b0110110100101010001: color_data = Z;
		19'b0110110100101010010: color_data = Z;
		19'b0110110100101010011: color_data = Z;
		19'b0110110100101010100: color_data = Z;
		19'b0110110100101010101: color_data = Z;
		19'b0110110100101010110: color_data = Z;
		19'b0110110100101010111: color_data = Z;
		19'b0110110100101011000: color_data = Z;
		19'b0110110100101011001: color_data = Z;
		19'b0110110100101011010: color_data = Z;
		19'b0110110100101011011: color_data = Z;
		19'b0110110100101011100: color_data = Z;
		19'b0110110100101011101: color_data = Z;
		19'b0110110100101011110: color_data = Z;
		19'b0110110100101011111: color_data = Z;
		19'b0110110100101100000: color_data = Z;
		19'b0110110100101100001: color_data = Z;
		19'b0110110100101100010: color_data = Z;
		19'b0110110100101100011: color_data = Z;
		19'b0110110100101100100: color_data = Z;
		19'b0110110100101100101: color_data = Z;
		19'b0110110100101100110: color_data = Z;
		19'b0110110100101100111: color_data = Z;
		19'b0110110100101101000: color_data = Z;
		19'b0110110100101101001: color_data = Z;
		19'b0110110100101101101: color_data = Z;
		19'b0110110100101101110: color_data = Z;
		19'b0110110100101101111: color_data = Z;
		19'b0110110100101110000: color_data = Z;
		19'b0110110100101110001: color_data = Z;
		19'b0110110100101110010: color_data = Z;
		19'b0110110100101110011: color_data = Z;
		19'b0110110100101110100: color_data = Z;
		19'b0110110100101110101: color_data = Z;
		19'b0110110100101110110: color_data = Z;
		19'b0110110100101110111: color_data = Z;
		19'b0110110100101111000: color_data = Z;
		19'b0110110100101111001: color_data = Z;
		19'b0110110100101111010: color_data = Z;
		19'b0110110100101111011: color_data = Z;
		19'b0110110100101111100: color_data = Z;
		19'b0110110100110000010: color_data = Z;
		19'b0110110100110000011: color_data = Z;
		19'b0110110100110000100: color_data = Z;
		19'b0110110100110000101: color_data = Z;
		19'b0110110100110000110: color_data = Z;
		19'b0110110100110000111: color_data = Z;
		19'b0110110100110001000: color_data = Z;
		19'b0110110100110001001: color_data = Z;
		19'b0110110100110001010: color_data = Z;
		19'b0110110100110001011: color_data = Z;
		19'b0110110100110001100: color_data = Z;
		19'b0110110100110001101: color_data = Z;
		19'b0110110100110001110: color_data = Z;
		19'b0110110100110001111: color_data = Z;
		19'b0110110100110010000: color_data = Z;
		19'b0110110100110010001: color_data = Z;
		19'b0110110100110010010: color_data = Z;
		19'b0110110100110010011: color_data = Z;
		19'b0110110100110010100: color_data = Z;
		19'b0110110100111010000: color_data = Z;
		19'b0110110100111010001: color_data = Z;
		19'b0110110100111010010: color_data = Z;
		19'b0110110100111010011: color_data = Z;
		19'b0110110100111010100: color_data = Z;
		19'b0110110100111010101: color_data = Z;
		19'b0110110100111010110: color_data = Z;
		19'b0110110100111010111: color_data = Z;
		19'b0110110110010100110: color_data = Z;
		19'b0110110110010100111: color_data = Z;
		19'b0110110110010101000: color_data = Z;
		19'b0110110110010101001: color_data = Z;
		19'b0110110110010101010: color_data = Z;
		19'b0110110110010101011: color_data = Z;
		19'b0110110110010101100: color_data = Z;
		19'b0110110110010110100: color_data = Z;
		19'b0110110110010110101: color_data = Z;
		19'b0110110110100011001: color_data = Z;
		19'b0110110110100011010: color_data = Z;
		19'b0110110110100011011: color_data = Z;
		19'b0110110110100011100: color_data = Z;
		19'b0110110110100011101: color_data = Z;
		19'b0110110110100011110: color_data = Z;
		19'b0110110110100011111: color_data = Z;
		19'b0110110110100100000: color_data = Z;
		19'b0110110110100100001: color_data = Z;
		19'b0110110110100100010: color_data = Z;
		19'b0110110110100100011: color_data = Z;
		19'b0110110110100100100: color_data = Z;
		19'b0110110110100100101: color_data = Z;
		19'b0110110110100100110: color_data = Z;
		19'b0110110110100100111: color_data = Z;
		19'b0110110110100101000: color_data = Z;
		19'b0110110110100101001: color_data = Z;
		19'b0110110110100101010: color_data = Z;
		19'b0110110110100101011: color_data = Z;
		19'b0110110110100101101: color_data = Z;
		19'b0110110110100101110: color_data = Z;
		19'b0110110110100101111: color_data = Z;
		19'b0110110110100110000: color_data = Z;
		19'b0110110110100110001: color_data = Z;
		19'b0110110110100110010: color_data = Z;
		19'b0110110110100110011: color_data = Z;
		19'b0110110110100110100: color_data = Z;
		19'b0110110110100110101: color_data = Z;
		19'b0110110110100110110: color_data = Z;
		19'b0110110110100110111: color_data = Z;
		19'b0110110110100111000: color_data = Z;
		19'b0110110110100111001: color_data = Z;
		19'b0110110110100111010: color_data = Z;
		19'b0110110110100111011: color_data = Z;
		19'b0110110110100111100: color_data = Z;
		19'b0110110110100111101: color_data = Z;
		19'b0110110110100111110: color_data = Z;
		19'b0110110110100111111: color_data = Z;
		19'b0110110110101000000: color_data = Z;
		19'b0110110110101000001: color_data = Z;
		19'b0110110110101000010: color_data = Z;
		19'b0110110110101000011: color_data = Z;
		19'b0110110110101000100: color_data = Z;
		19'b0110110110101000101: color_data = Z;
		19'b0110110110101000110: color_data = Z;
		19'b0110110110101000111: color_data = Z;
		19'b0110110110101001000: color_data = Z;
		19'b0110110110101001001: color_data = Z;
		19'b0110110110101001010: color_data = Z;
		19'b0110110110101001011: color_data = Z;
		19'b0110110110101001100: color_data = Z;
		19'b0110110110101001101: color_data = Z;
		19'b0110110110101001110: color_data = Z;
		19'b0110110110101001111: color_data = Z;
		19'b0110110110101010000: color_data = Z;
		19'b0110110110101010001: color_data = Z;
		19'b0110110110101010010: color_data = Z;
		19'b0110110110101010011: color_data = Z;
		19'b0110110110101010100: color_data = Z;
		19'b0110110110101010101: color_data = Z;
		19'b0110110110101010110: color_data = Z;
		19'b0110110110101010111: color_data = Z;
		19'b0110110110101011000: color_data = Z;
		19'b0110110110101011001: color_data = Z;
		19'b0110110110101011010: color_data = Z;
		19'b0110110110101011011: color_data = Z;
		19'b0110110110101011100: color_data = Z;
		19'b0110110110101011101: color_data = Z;
		19'b0110110110101011110: color_data = Z;
		19'b0110110110101011111: color_data = Z;
		19'b0110110110101100000: color_data = Z;
		19'b0110110110101100001: color_data = Z;
		19'b0110110110101100010: color_data = Z;
		19'b0110110110101100011: color_data = Z;
		19'b0110110110101100100: color_data = Z;
		19'b0110110110101100101: color_data = Z;
		19'b0110110110101100110: color_data = Z;
		19'b0110110110101100111: color_data = Z;
		19'b0110110110101101000: color_data = Z;
		19'b0110110110101101001: color_data = Z;
		19'b0110110110101101101: color_data = Z;
		19'b0110110110101101110: color_data = Z;
		19'b0110110110101101111: color_data = Z;
		19'b0110110110101110000: color_data = Z;
		19'b0110110110101110001: color_data = Z;
		19'b0110110110101110010: color_data = Z;
		19'b0110110110101110011: color_data = Z;
		19'b0110110110101110100: color_data = Z;
		19'b0110110110101110101: color_data = Z;
		19'b0110110110101110110: color_data = Z;
		19'b0110110110101110111: color_data = Z;
		19'b0110110110101111000: color_data = Z;
		19'b0110110110101111001: color_data = Z;
		19'b0110110110101111010: color_data = Z;
		19'b0110110110101111011: color_data = Z;
		19'b0110110110101111100: color_data = Z;
		19'b0110110110110000011: color_data = Z;
		19'b0110110110110000100: color_data = Z;
		19'b0110110110110000101: color_data = Z;
		19'b0110110110110000110: color_data = Z;
		19'b0110110110110000111: color_data = Z;
		19'b0110110110110001000: color_data = Z;
		19'b0110110110110001001: color_data = Z;
		19'b0110110110110001010: color_data = Z;
		19'b0110110110110001011: color_data = Z;
		19'b0110110110110001100: color_data = Z;
		19'b0110110110110001101: color_data = Z;
		19'b0110110110110001110: color_data = Z;
		19'b0110110110110001111: color_data = Z;
		19'b0110110110110010000: color_data = Z;
		19'b0110110110110010001: color_data = Z;
		19'b0110110110110010010: color_data = Z;
		19'b0110110110110010011: color_data = Z;
		19'b0110110110110010100: color_data = Z;
		19'b0110110110110010101: color_data = Z;
		19'b0110110110110010110: color_data = Z;
		19'b0110110110111010000: color_data = Z;
		19'b0110110110111010001: color_data = Z;
		19'b0110110110111010010: color_data = Z;
		19'b0110110110111010011: color_data = Z;
		19'b0110110110111010100: color_data = Z;
		19'b0110110110111010101: color_data = Z;
		19'b0110110110111010110: color_data = Z;
		19'b0110110110111010111: color_data = Z;
		19'b0110111000010100111: color_data = Z;
		19'b0110111000010101000: color_data = Z;
		19'b0110111000010101001: color_data = Z;
		19'b0110111000010101010: color_data = Z;
		19'b0110111000010101011: color_data = Z;
		19'b0110111000010101100: color_data = Z;
		19'b0110111000010101101: color_data = Z;
		19'b0110111000010110101: color_data = Z;
		19'b0110111000010110110: color_data = Z;
		19'b0110111000100011001: color_data = Z;
		19'b0110111000100011010: color_data = Z;
		19'b0110111000100011011: color_data = Z;
		19'b0110111000100011100: color_data = Z;
		19'b0110111000100011101: color_data = Z;
		19'b0110111000100011110: color_data = Z;
		19'b0110111000100011111: color_data = Z;
		19'b0110111000100100000: color_data = Z;
		19'b0110111000100100001: color_data = Z;
		19'b0110111000100100010: color_data = Z;
		19'b0110111000100100011: color_data = Z;
		19'b0110111000100100100: color_data = Z;
		19'b0110111000100100101: color_data = Z;
		19'b0110111000100100110: color_data = Z;
		19'b0110111000100100111: color_data = Z;
		19'b0110111000100101000: color_data = Z;
		19'b0110111000100101001: color_data = Z;
		19'b0110111000100101010: color_data = Z;
		19'b0110111000100101011: color_data = Z;
		19'b0110111000100101101: color_data = Z;
		19'b0110111000100101110: color_data = Z;
		19'b0110111000100101111: color_data = Z;
		19'b0110111000100110000: color_data = Z;
		19'b0110111000100110001: color_data = Z;
		19'b0110111000100110010: color_data = Z;
		19'b0110111000100110011: color_data = Z;
		19'b0110111000100110100: color_data = Z;
		19'b0110111000100110101: color_data = Z;
		19'b0110111000100110110: color_data = Z;
		19'b0110111000100110111: color_data = Z;
		19'b0110111000100111000: color_data = Z;
		19'b0110111000100111001: color_data = Z;
		19'b0110111000100111010: color_data = Z;
		19'b0110111000100111011: color_data = Z;
		19'b0110111000100111100: color_data = Z;
		19'b0110111000100111101: color_data = Z;
		19'b0110111000100111110: color_data = Z;
		19'b0110111000100111111: color_data = Z;
		19'b0110111000101000000: color_data = Z;
		19'b0110111000101000001: color_data = Z;
		19'b0110111000101000010: color_data = Z;
		19'b0110111000101000011: color_data = Z;
		19'b0110111000101000100: color_data = Z;
		19'b0110111000101000101: color_data = Z;
		19'b0110111000101000110: color_data = Z;
		19'b0110111000101000111: color_data = Z;
		19'b0110111000101001000: color_data = Z;
		19'b0110111000101001001: color_data = Z;
		19'b0110111000101001010: color_data = Z;
		19'b0110111000101001011: color_data = Z;
		19'b0110111000101001100: color_data = Z;
		19'b0110111000101001101: color_data = Z;
		19'b0110111000101001110: color_data = Z;
		19'b0110111000101001111: color_data = Z;
		19'b0110111000101010000: color_data = Z;
		19'b0110111000101010001: color_data = Z;
		19'b0110111000101010010: color_data = Z;
		19'b0110111000101010011: color_data = Z;
		19'b0110111000101010100: color_data = Z;
		19'b0110111000101010101: color_data = Z;
		19'b0110111000101010110: color_data = Z;
		19'b0110111000101010111: color_data = Z;
		19'b0110111000101011000: color_data = Z;
		19'b0110111000101011001: color_data = Z;
		19'b0110111000101011010: color_data = Z;
		19'b0110111000101011011: color_data = Z;
		19'b0110111000101011100: color_data = Z;
		19'b0110111000101011101: color_data = Z;
		19'b0110111000101011110: color_data = Z;
		19'b0110111000101011111: color_data = Z;
		19'b0110111000101100000: color_data = Z;
		19'b0110111000101100001: color_data = Z;
		19'b0110111000101100010: color_data = Z;
		19'b0110111000101100011: color_data = Z;
		19'b0110111000101100100: color_data = Z;
		19'b0110111000101100101: color_data = Z;
		19'b0110111000101100110: color_data = Z;
		19'b0110111000101100111: color_data = Z;
		19'b0110111000101101000: color_data = Z;
		19'b0110111000101101001: color_data = Z;
		19'b0110111000101101010: color_data = Z;
		19'b0110111000101101101: color_data = Z;
		19'b0110111000101101110: color_data = Z;
		19'b0110111000101101111: color_data = Z;
		19'b0110111000101110000: color_data = Z;
		19'b0110111000101110001: color_data = Z;
		19'b0110111000101110010: color_data = Z;
		19'b0110111000101110011: color_data = Z;
		19'b0110111000101110100: color_data = Z;
		19'b0110111000101110101: color_data = Z;
		19'b0110111000101110110: color_data = Z;
		19'b0110111000101110111: color_data = Z;
		19'b0110111000101111000: color_data = Z;
		19'b0110111000101111001: color_data = Z;
		19'b0110111000101111010: color_data = Z;
		19'b0110111000101111011: color_data = Z;
		19'b0110111000101111100: color_data = Z;
		19'b0110111000101111101: color_data = Z;
		19'b0110111000110000011: color_data = Z;
		19'b0110111000110000100: color_data = Z;
		19'b0110111000110000101: color_data = Z;
		19'b0110111000110000110: color_data = Z;
		19'b0110111000110000111: color_data = Z;
		19'b0110111000110001000: color_data = Z;
		19'b0110111000110001001: color_data = Z;
		19'b0110111000110001010: color_data = Z;
		19'b0110111000110001011: color_data = Z;
		19'b0110111000110001100: color_data = Z;
		19'b0110111000110001101: color_data = Z;
		19'b0110111000110001110: color_data = Z;
		19'b0110111000110001111: color_data = Z;
		19'b0110111000110010000: color_data = Z;
		19'b0110111000110010001: color_data = Z;
		19'b0110111000110010010: color_data = Z;
		19'b0110111000110010011: color_data = Z;
		19'b0110111000110010100: color_data = Z;
		19'b0110111000110010101: color_data = Z;
		19'b0110111000110010110: color_data = Z;
		19'b0110111000110010111: color_data = Z;
		19'b0110111000110011000: color_data = Z;
		19'b0110111000110101111: color_data = Z;
		19'b0110111000110110000: color_data = Z;
		19'b0110111000110110001: color_data = Z;
		19'b0110111000110110010: color_data = Z;
		19'b0110111000111010001: color_data = Z;
		19'b0110111000111010010: color_data = Z;
		19'b0110111000111010011: color_data = Z;
		19'b0110111000111010100: color_data = Z;
		19'b0110111000111010101: color_data = Z;
		19'b0110111000111010110: color_data = Z;
		19'b0110111000111010111: color_data = Z;
		19'b0110111010010100111: color_data = Z;
		19'b0110111010010101000: color_data = Z;
		19'b0110111010010101001: color_data = Z;
		19'b0110111010010101010: color_data = Z;
		19'b0110111010010101011: color_data = Z;
		19'b0110111010010101100: color_data = Z;
		19'b0110111010010101101: color_data = Z;
		19'b0110111010010110101: color_data = Z;
		19'b0110111010010110110: color_data = Z;
		19'b0110111010010111011: color_data = Z;
		19'b0110111010100010011: color_data = Z;
		19'b0110111010100010100: color_data = Z;
		19'b0110111010100010101: color_data = Z;
		19'b0110111010100011001: color_data = Z;
		19'b0110111010100011010: color_data = Z;
		19'b0110111010100011011: color_data = Z;
		19'b0110111010100011100: color_data = Z;
		19'b0110111010100011101: color_data = Z;
		19'b0110111010100011110: color_data = Z;
		19'b0110111010100011111: color_data = Z;
		19'b0110111010100100000: color_data = Z;
		19'b0110111010100100001: color_data = Z;
		19'b0110111010100100010: color_data = Z;
		19'b0110111010100100100: color_data = Z;
		19'b0110111010100100101: color_data = Z;
		19'b0110111010100100110: color_data = Z;
		19'b0110111010100100111: color_data = Z;
		19'b0110111010100101000: color_data = Z;
		19'b0110111010100101001: color_data = Z;
		19'b0110111010100101010: color_data = Z;
		19'b0110111010100101011: color_data = Z;
		19'b0110111010100101101: color_data = Z;
		19'b0110111010100101110: color_data = Z;
		19'b0110111010100101111: color_data = Z;
		19'b0110111010100110000: color_data = Z;
		19'b0110111010100110001: color_data = Z;
		19'b0110111010100110010: color_data = Z;
		19'b0110111010100110011: color_data = Z;
		19'b0110111010100110100: color_data = Z;
		19'b0110111010100110101: color_data = Z;
		19'b0110111010100110110: color_data = Z;
		19'b0110111010100110111: color_data = Z;
		19'b0110111010100111000: color_data = Z;
		19'b0110111010100111001: color_data = Z;
		19'b0110111010100111010: color_data = Z;
		19'b0110111010100111011: color_data = Z;
		19'b0110111010100111100: color_data = Z;
		19'b0110111010100111101: color_data = Z;
		19'b0110111010100111110: color_data = Z;
		19'b0110111010100111111: color_data = Z;
		19'b0110111010101000000: color_data = Z;
		19'b0110111010101000001: color_data = Z;
		19'b0110111010101000010: color_data = Z;
		19'b0110111010101000011: color_data = Z;
		19'b0110111010101000100: color_data = Z;
		19'b0110111010101000101: color_data = Z;
		19'b0110111010101000110: color_data = Z;
		19'b0110111010101000111: color_data = Z;
		19'b0110111010101001000: color_data = Z;
		19'b0110111010101001001: color_data = Z;
		19'b0110111010101001010: color_data = Z;
		19'b0110111010101001011: color_data = Z;
		19'b0110111010101001100: color_data = Z;
		19'b0110111010101001101: color_data = Z;
		19'b0110111010101001110: color_data = Z;
		19'b0110111010101001111: color_data = Z;
		19'b0110111010101010000: color_data = Z;
		19'b0110111010101010001: color_data = Z;
		19'b0110111010101010010: color_data = Z;
		19'b0110111010101010011: color_data = Z;
		19'b0110111010101010100: color_data = Z;
		19'b0110111010101010101: color_data = Z;
		19'b0110111010101010110: color_data = Z;
		19'b0110111010101010111: color_data = Z;
		19'b0110111010101011000: color_data = Z;
		19'b0110111010101011001: color_data = Z;
		19'b0110111010101011010: color_data = Z;
		19'b0110111010101011011: color_data = Z;
		19'b0110111010101011100: color_data = Z;
		19'b0110111010101011101: color_data = Z;
		19'b0110111010101011110: color_data = Z;
		19'b0110111010101011111: color_data = Z;
		19'b0110111010101100000: color_data = Z;
		19'b0110111010101100001: color_data = Z;
		19'b0110111010101100010: color_data = Z;
		19'b0110111010101100011: color_data = Z;
		19'b0110111010101100100: color_data = Z;
		19'b0110111010101100101: color_data = Z;
		19'b0110111010101100110: color_data = Z;
		19'b0110111010101100111: color_data = Z;
		19'b0110111010101101000: color_data = Z;
		19'b0110111010101101001: color_data = Z;
		19'b0110111010101101010: color_data = Z;
		19'b0110111010101101101: color_data = Z;
		19'b0110111010101101110: color_data = Z;
		19'b0110111010101101111: color_data = Z;
		19'b0110111010101110000: color_data = Z;
		19'b0110111010101110001: color_data = Z;
		19'b0110111010101110010: color_data = Z;
		19'b0110111010101110011: color_data = Z;
		19'b0110111010101110100: color_data = Z;
		19'b0110111010101110101: color_data = Z;
		19'b0110111010101110110: color_data = Z;
		19'b0110111010101110111: color_data = Z;
		19'b0110111010101111000: color_data = Z;
		19'b0110111010101111001: color_data = Z;
		19'b0110111010101111010: color_data = Z;
		19'b0110111010101111011: color_data = Z;
		19'b0110111010101111100: color_data = Z;
		19'b0110111010101111101: color_data = Z;
		19'b0110111010101111110: color_data = Z;
		19'b0110111010110000100: color_data = Z;
		19'b0110111010110000101: color_data = Z;
		19'b0110111010110000110: color_data = Z;
		19'b0110111010110000111: color_data = Z;
		19'b0110111010110001000: color_data = Z;
		19'b0110111010110001001: color_data = Z;
		19'b0110111010110001010: color_data = Z;
		19'b0110111010110001011: color_data = Z;
		19'b0110111010110001100: color_data = Z;
		19'b0110111010110001101: color_data = Z;
		19'b0110111010110001110: color_data = Z;
		19'b0110111010110001111: color_data = Z;
		19'b0110111010110010000: color_data = Z;
		19'b0110111010110010001: color_data = Z;
		19'b0110111010110010010: color_data = Z;
		19'b0110111010110010011: color_data = Z;
		19'b0110111010110010100: color_data = Z;
		19'b0110111010110010101: color_data = Z;
		19'b0110111010110010110: color_data = Z;
		19'b0110111010110010111: color_data = Z;
		19'b0110111010110011000: color_data = Z;
		19'b0110111010110011001: color_data = Z;
		19'b0110111010110011010: color_data = Z;
		19'b0110111010110011011: color_data = Z;
		19'b0110111010110011100: color_data = Z;
		19'b0110111010110101111: color_data = Z;
		19'b0110111010110110000: color_data = Z;
		19'b0110111010110110001: color_data = Z;
		19'b0110111010110110010: color_data = Z;
		19'b0110111010110111100: color_data = Z;
		19'b0110111010110111101: color_data = Z;
		19'b0110111010110111110: color_data = Z;
		19'b0110111010111010010: color_data = Z;
		19'b0110111010111010011: color_data = Z;
		19'b0110111010111010100: color_data = Z;
		19'b0110111010111010101: color_data = Z;
		19'b0110111010111010110: color_data = Z;
		19'b0110111010111010111: color_data = Z;
		19'b0110111100010101000: color_data = Z;
		19'b0110111100010101001: color_data = Z;
		19'b0110111100010101010: color_data = Z;
		19'b0110111100010101011: color_data = Z;
		19'b0110111100010101100: color_data = Z;
		19'b0110111100010101101: color_data = Z;
		19'b0110111100010110101: color_data = Z;
		19'b0110111100010110110: color_data = Z;
		19'b0110111100010110111: color_data = Z;
		19'b0110111100010111000: color_data = Z;
		19'b0110111100010111001: color_data = Z;
		19'b0110111100010111010: color_data = Z;
		19'b0110111100010111011: color_data = Z;
		19'b0110111100010111100: color_data = Z;
		19'b0110111100100010011: color_data = Z;
		19'b0110111100100010100: color_data = Z;
		19'b0110111100100010101: color_data = Z;
		19'b0110111100100010110: color_data = Z;
		19'b0110111100100011001: color_data = Z;
		19'b0110111100100011010: color_data = Z;
		19'b0110111100100011011: color_data = Z;
		19'b0110111100100011100: color_data = Z;
		19'b0110111100100011101: color_data = Z;
		19'b0110111100100011110: color_data = Z;
		19'b0110111100100011111: color_data = Z;
		19'b0110111100100100000: color_data = Z;
		19'b0110111100100100001: color_data = Z;
		19'b0110111100100100011: color_data = Z;
		19'b0110111100100100100: color_data = Z;
		19'b0110111100100100101: color_data = Z;
		19'b0110111100100100110: color_data = Z;
		19'b0110111100100100111: color_data = Z;
		19'b0110111100100101000: color_data = Z;
		19'b0110111100100101001: color_data = Z;
		19'b0110111100100101010: color_data = Z;
		19'b0110111100100101100: color_data = Z;
		19'b0110111100100101101: color_data = Z;
		19'b0110111100100101110: color_data = Z;
		19'b0110111100100101111: color_data = Z;
		19'b0110111100100110000: color_data = Z;
		19'b0110111100100110001: color_data = Z;
		19'b0110111100100110010: color_data = Z;
		19'b0110111100100110011: color_data = Z;
		19'b0110111100100110100: color_data = Z;
		19'b0110111100100110101: color_data = Z;
		19'b0110111100100110110: color_data = Z;
		19'b0110111100100110111: color_data = Z;
		19'b0110111100100111000: color_data = Z;
		19'b0110111100100111001: color_data = Z;
		19'b0110111100100111010: color_data = Z;
		19'b0110111100100111011: color_data = Z;
		19'b0110111100100111100: color_data = Z;
		19'b0110111100100111101: color_data = Z;
		19'b0110111100100111110: color_data = Z;
		19'b0110111100100111111: color_data = Z;
		19'b0110111100101000000: color_data = Z;
		19'b0110111100101000001: color_data = Z;
		19'b0110111100101000010: color_data = Z;
		19'b0110111100101000011: color_data = Z;
		19'b0110111100101000100: color_data = Z;
		19'b0110111100101000101: color_data = Z;
		19'b0110111100101000110: color_data = Z;
		19'b0110111100101000111: color_data = Z;
		19'b0110111100101001000: color_data = Z;
		19'b0110111100101001001: color_data = Z;
		19'b0110111100101001010: color_data = Z;
		19'b0110111100101001011: color_data = Z;
		19'b0110111100101001100: color_data = Z;
		19'b0110111100101001101: color_data = Z;
		19'b0110111100101001110: color_data = Z;
		19'b0110111100101001111: color_data = Z;
		19'b0110111100101010000: color_data = Z;
		19'b0110111100101010001: color_data = Z;
		19'b0110111100101010010: color_data = Z;
		19'b0110111100101010011: color_data = Z;
		19'b0110111100101010100: color_data = Z;
		19'b0110111100101010101: color_data = Z;
		19'b0110111100101010110: color_data = Z;
		19'b0110111100101010111: color_data = Z;
		19'b0110111100101011000: color_data = Z;
		19'b0110111100101011001: color_data = Z;
		19'b0110111100101011010: color_data = Z;
		19'b0110111100101011011: color_data = Z;
		19'b0110111100101011100: color_data = Z;
		19'b0110111100101011101: color_data = Z;
		19'b0110111100101011110: color_data = Z;
		19'b0110111100101011111: color_data = Z;
		19'b0110111100101100000: color_data = Z;
		19'b0110111100101100001: color_data = Z;
		19'b0110111100101100010: color_data = Z;
		19'b0110111100101100011: color_data = Z;
		19'b0110111100101100100: color_data = Z;
		19'b0110111100101100101: color_data = Z;
		19'b0110111100101100110: color_data = Z;
		19'b0110111100101100111: color_data = Z;
		19'b0110111100101101000: color_data = Z;
		19'b0110111100101101001: color_data = Z;
		19'b0110111100101101010: color_data = Z;
		19'b0110111100101101101: color_data = Z;
		19'b0110111100101101110: color_data = Z;
		19'b0110111100101101111: color_data = Z;
		19'b0110111100101110000: color_data = Z;
		19'b0110111100101110001: color_data = Z;
		19'b0110111100101110010: color_data = Z;
		19'b0110111100101110011: color_data = Z;
		19'b0110111100101110100: color_data = Z;
		19'b0110111100101110101: color_data = Z;
		19'b0110111100101110110: color_data = Z;
		19'b0110111100101110111: color_data = Z;
		19'b0110111100101111000: color_data = Z;
		19'b0110111100101111001: color_data = Z;
		19'b0110111100101111010: color_data = Z;
		19'b0110111100101111011: color_data = Z;
		19'b0110111100101111100: color_data = Z;
		19'b0110111100101111101: color_data = Z;
		19'b0110111100101111110: color_data = Z;
		19'b0110111100101111111: color_data = Z;
		19'b0110111100110000101: color_data = Z;
		19'b0110111100110000110: color_data = Z;
		19'b0110111100110000111: color_data = Z;
		19'b0110111100110001000: color_data = Z;
		19'b0110111100110001001: color_data = Z;
		19'b0110111100110001010: color_data = Z;
		19'b0110111100110001011: color_data = Z;
		19'b0110111100110001100: color_data = Z;
		19'b0110111100110001101: color_data = Z;
		19'b0110111100110001110: color_data = Z;
		19'b0110111100110001111: color_data = Z;
		19'b0110111100110010000: color_data = Z;
		19'b0110111100110010001: color_data = Z;
		19'b0110111100110010010: color_data = Z;
		19'b0110111100110010011: color_data = Z;
		19'b0110111100110010100: color_data = Z;
		19'b0110111100110010101: color_data = Z;
		19'b0110111100110010110: color_data = Z;
		19'b0110111100110010111: color_data = Z;
		19'b0110111100110011000: color_data = Z;
		19'b0110111100110011001: color_data = Z;
		19'b0110111100110011010: color_data = Z;
		19'b0110111100110011011: color_data = Z;
		19'b0110111100110011100: color_data = Z;
		19'b0110111100110011101: color_data = Z;
		19'b0110111100110011110: color_data = Z;
		19'b0110111100110111010: color_data = Z;
		19'b0110111100110111011: color_data = Z;
		19'b0110111100110111100: color_data = Z;
		19'b0110111100110111101: color_data = Z;
		19'b0110111100111010011: color_data = Z;
		19'b0110111100111010100: color_data = Z;
		19'b0110111100111010101: color_data = Z;
		19'b0110111100111010110: color_data = Z;
		19'b0110111100111010111: color_data = Z;
		19'b0110111110010101000: color_data = Z;
		19'b0110111110010101001: color_data = Z;
		19'b0110111110010101010: color_data = Z;
		19'b0110111110010101011: color_data = Z;
		19'b0110111110010101100: color_data = Z;
		19'b0110111110010101101: color_data = Z;
		19'b0110111110010101110: color_data = Z;
		19'b0110111110010110101: color_data = Z;
		19'b0110111110010110110: color_data = Z;
		19'b0110111110010110111: color_data = Z;
		19'b0110111110010111000: color_data = Z;
		19'b0110111110010111001: color_data = Z;
		19'b0110111110010111010: color_data = Z;
		19'b0110111110010111011: color_data = Z;
		19'b0110111110010111100: color_data = Z;
		19'b0110111110010111101: color_data = Z;
		19'b0110111110100010011: color_data = Z;
		19'b0110111110100010100: color_data = Z;
		19'b0110111110100010101: color_data = Z;
		19'b0110111110100010110: color_data = Z;
		19'b0110111110100011001: color_data = Z;
		19'b0110111110100011010: color_data = Z;
		19'b0110111110100011011: color_data = Z;
		19'b0110111110100011100: color_data = Z;
		19'b0110111110100011101: color_data = Z;
		19'b0110111110100011110: color_data = Z;
		19'b0110111110100011111: color_data = Z;
		19'b0110111110100100000: color_data = Z;
		19'b0110111110100100001: color_data = Z;
		19'b0110111110100100011: color_data = Z;
		19'b0110111110100100100: color_data = Z;
		19'b0110111110100100101: color_data = Z;
		19'b0110111110100100110: color_data = Z;
		19'b0110111110100100111: color_data = Z;
		19'b0110111110100101000: color_data = Z;
		19'b0110111110100101001: color_data = Z;
		19'b0110111110100101010: color_data = Z;
		19'b0110111110100101100: color_data = Z;
		19'b0110111110100101101: color_data = Z;
		19'b0110111110100101110: color_data = Z;
		19'b0110111110100101111: color_data = Z;
		19'b0110111110100110000: color_data = Z;
		19'b0110111110100110001: color_data = Z;
		19'b0110111110100110010: color_data = Z;
		19'b0110111110100110011: color_data = Z;
		19'b0110111110100110100: color_data = Z;
		19'b0110111110100110101: color_data = Z;
		19'b0110111110100110110: color_data = Z;
		19'b0110111110100110111: color_data = Z;
		19'b0110111110100111000: color_data = Z;
		19'b0110111110100111001: color_data = Z;
		19'b0110111110100111010: color_data = Z;
		19'b0110111110100111011: color_data = Z;
		19'b0110111110100111100: color_data = Z;
		19'b0110111110100111101: color_data = Z;
		19'b0110111110100111110: color_data = Z;
		19'b0110111110100111111: color_data = Z;
		19'b0110111110101000000: color_data = Z;
		19'b0110111110101000001: color_data = Z;
		19'b0110111110101000010: color_data = Z;
		19'b0110111110101000011: color_data = Z;
		19'b0110111110101000100: color_data = Z;
		19'b0110111110101000101: color_data = Z;
		19'b0110111110101000110: color_data = Z;
		19'b0110111110101000111: color_data = Z;
		19'b0110111110101001000: color_data = Z;
		19'b0110111110101001001: color_data = Z;
		19'b0110111110101001010: color_data = Z;
		19'b0110111110101001011: color_data = Z;
		19'b0110111110101001100: color_data = Z;
		19'b0110111110101001101: color_data = Z;
		19'b0110111110101001110: color_data = Z;
		19'b0110111110101001111: color_data = Z;
		19'b0110111110101010000: color_data = Z;
		19'b0110111110101010001: color_data = Z;
		19'b0110111110101010010: color_data = Z;
		19'b0110111110101010011: color_data = Z;
		19'b0110111110101010100: color_data = Z;
		19'b0110111110101010101: color_data = Z;
		19'b0110111110101010110: color_data = Z;
		19'b0110111110101010111: color_data = Z;
		19'b0110111110101011000: color_data = Z;
		19'b0110111110101011001: color_data = Z;
		19'b0110111110101011010: color_data = Z;
		19'b0110111110101011011: color_data = Z;
		19'b0110111110101011100: color_data = Z;
		19'b0110111110101011101: color_data = Z;
		19'b0110111110101011110: color_data = Z;
		19'b0110111110101011111: color_data = Z;
		19'b0110111110101100000: color_data = Z;
		19'b0110111110101100001: color_data = Z;
		19'b0110111110101100010: color_data = Z;
		19'b0110111110101100011: color_data = Z;
		19'b0110111110101100100: color_data = Z;
		19'b0110111110101100101: color_data = Z;
		19'b0110111110101100110: color_data = Z;
		19'b0110111110101100111: color_data = Z;
		19'b0110111110101101000: color_data = Z;
		19'b0110111110101101001: color_data = Z;
		19'b0110111110101101010: color_data = Z;
		19'b0110111110101101101: color_data = Z;
		19'b0110111110101101110: color_data = Z;
		19'b0110111110101101111: color_data = Z;
		19'b0110111110101110000: color_data = Z;
		19'b0110111110101110001: color_data = Z;
		19'b0110111110101110010: color_data = Z;
		19'b0110111110101110011: color_data = Z;
		19'b0110111110101110100: color_data = Z;
		19'b0110111110101110101: color_data = Z;
		19'b0110111110101110110: color_data = Z;
		19'b0110111110101110111: color_data = Z;
		19'b0110111110101111000: color_data = Z;
		19'b0110111110101111001: color_data = Z;
		19'b0110111110101111010: color_data = Z;
		19'b0110111110101111011: color_data = Z;
		19'b0110111110101111100: color_data = Z;
		19'b0110111110101111101: color_data = Z;
		19'b0110111110101111110: color_data = Z;
		19'b0110111110101111111: color_data = Z;
		19'b0110111110110000000: color_data = Z;
		19'b0110111110110000101: color_data = Z;
		19'b0110111110110000110: color_data = Z;
		19'b0110111110110000111: color_data = Z;
		19'b0110111110110001000: color_data = Z;
		19'b0110111110110001001: color_data = Z;
		19'b0110111110110001010: color_data = Z;
		19'b0110111110110001011: color_data = Z;
		19'b0110111110110001100: color_data = Z;
		19'b0110111110110001101: color_data = Z;
		19'b0110111110110001110: color_data = Z;
		19'b0110111110110001111: color_data = Z;
		19'b0110111110110010000: color_data = Z;
		19'b0110111110110010001: color_data = Z;
		19'b0110111110110010010: color_data = Z;
		19'b0110111110110010011: color_data = Z;
		19'b0110111110110010100: color_data = Z;
		19'b0110111110110010101: color_data = Z;
		19'b0110111110110010110: color_data = Z;
		19'b0110111110110010111: color_data = Z;
		19'b0110111110110011000: color_data = Z;
		19'b0110111110110011001: color_data = Z;
		19'b0110111110110011010: color_data = Z;
		19'b0110111110110011011: color_data = Z;
		19'b0110111110110011100: color_data = Z;
		19'b0110111110110011101: color_data = Z;
		19'b0110111110110011110: color_data = Z;
		19'b0110111110110011111: color_data = Z;
		19'b0110111110110100000: color_data = Z;
		19'b0110111110110111000: color_data = Z;
		19'b0110111110110111001: color_data = Z;
		19'b0110111110110111010: color_data = Z;
		19'b0110111110110111011: color_data = Z;
		19'b0110111110110111100: color_data = Z;
		19'b0110111110110111101: color_data = Z;
		19'b0110111110110111110: color_data = Z;
		19'b0110111110111010100: color_data = Z;
		19'b0110111110111010101: color_data = Z;
		19'b0110111110111010110: color_data = Z;
		19'b0110111110111010111: color_data = Z;
		19'b0111000000010101000: color_data = Z;
		19'b0111000000010101001: color_data = Z;
		19'b0111000000010101010: color_data = Z;
		19'b0111000000010101011: color_data = Z;
		19'b0111000000010101100: color_data = Z;
		19'b0111000000010101101: color_data = Z;
		19'b0111000000010101110: color_data = Z;
		19'b0111000000010110010: color_data = Z;
		19'b0111000000010110011: color_data = Z;
		19'b0111000000010110101: color_data = Z;
		19'b0111000000010110110: color_data = Z;
		19'b0111000000010110111: color_data = Z;
		19'b0111000000010111000: color_data = Z;
		19'b0111000000010111001: color_data = Z;
		19'b0111000000010111010: color_data = Z;
		19'b0111000000010111011: color_data = Z;
		19'b0111000000010111100: color_data = Z;
		19'b0111000000010111101: color_data = Z;
		19'b0111000000100010011: color_data = Z;
		19'b0111000000100010100: color_data = Z;
		19'b0111000000100010101: color_data = Z;
		19'b0111000000100010110: color_data = Z;
		19'b0111000000100011001: color_data = Z;
		19'b0111000000100011010: color_data = Z;
		19'b0111000000100011011: color_data = Z;
		19'b0111000000100011100: color_data = Z;
		19'b0111000000100011101: color_data = Z;
		19'b0111000000100011110: color_data = Z;
		19'b0111000000100011111: color_data = Z;
		19'b0111000000100100000: color_data = Z;
		19'b0111000000100100001: color_data = Z;
		19'b0111000000100100010: color_data = Z;
		19'b0111000000100100011: color_data = Z;
		19'b0111000000100100100: color_data = Z;
		19'b0111000000100100101: color_data = Z;
		19'b0111000000100100110: color_data = Z;
		19'b0111000000100100111: color_data = Z;
		19'b0111000000100101000: color_data = Z;
		19'b0111000000100101001: color_data = Z;
		19'b0111000000100101100: color_data = Z;
		19'b0111000000100101101: color_data = Z;
		19'b0111000000100101110: color_data = Z;
		19'b0111000000100101111: color_data = Z;
		19'b0111000000100110000: color_data = Z;
		19'b0111000000100110001: color_data = Z;
		19'b0111000000100110010: color_data = Z;
		19'b0111000000100110011: color_data = Z;
		19'b0111000000100110100: color_data = Z;
		19'b0111000000100110101: color_data = Z;
		19'b0111000000100110110: color_data = Z;
		19'b0111000000100110111: color_data = Z;
		19'b0111000000100111000: color_data = Z;
		19'b0111000000100111001: color_data = Z;
		19'b0111000000100111010: color_data = Z;
		19'b0111000000100111011: color_data = Z;
		19'b0111000000100111100: color_data = Z;
		19'b0111000000100111101: color_data = Z;
		19'b0111000000100111110: color_data = Z;
		19'b0111000000100111111: color_data = Z;
		19'b0111000000101000000: color_data = Z;
		19'b0111000000101000001: color_data = Z;
		19'b0111000000101000010: color_data = Z;
		19'b0111000000101000011: color_data = Z;
		19'b0111000000101000100: color_data = Z;
		19'b0111000000101000101: color_data = Z;
		19'b0111000000101000110: color_data = Z;
		19'b0111000000101000111: color_data = Z;
		19'b0111000000101001000: color_data = Z;
		19'b0111000000101001001: color_data = Z;
		19'b0111000000101001010: color_data = Z;
		19'b0111000000101001011: color_data = Z;
		19'b0111000000101001100: color_data = Z;
		19'b0111000000101001101: color_data = Z;
		19'b0111000000101001110: color_data = Z;
		19'b0111000000101001111: color_data = Z;
		19'b0111000000101010000: color_data = Z;
		19'b0111000000101010001: color_data = Z;
		19'b0111000000101010010: color_data = Z;
		19'b0111000000101010011: color_data = Z;
		19'b0111000000101010100: color_data = Z;
		19'b0111000000101010101: color_data = Z;
		19'b0111000000101010110: color_data = Z;
		19'b0111000000101010111: color_data = Z;
		19'b0111000000101011000: color_data = Z;
		19'b0111000000101011001: color_data = Z;
		19'b0111000000101011010: color_data = Z;
		19'b0111000000101011011: color_data = Z;
		19'b0111000000101011100: color_data = Z;
		19'b0111000000101011101: color_data = Z;
		19'b0111000000101011110: color_data = Z;
		19'b0111000000101011111: color_data = Z;
		19'b0111000000101100000: color_data = Z;
		19'b0111000000101100001: color_data = Z;
		19'b0111000000101100010: color_data = Z;
		19'b0111000000101100011: color_data = Z;
		19'b0111000000101100100: color_data = Z;
		19'b0111000000101100101: color_data = Z;
		19'b0111000000101100110: color_data = Z;
		19'b0111000000101100111: color_data = Z;
		19'b0111000000101101000: color_data = Z;
		19'b0111000000101101001: color_data = Z;
		19'b0111000000101101010: color_data = Z;
		19'b0111000000101101011: color_data = Z;
		19'b0111000000101101101: color_data = Z;
		19'b0111000000101101110: color_data = Z;
		19'b0111000000101101111: color_data = Z;
		19'b0111000000101110000: color_data = Z;
		19'b0111000000101110001: color_data = Z;
		19'b0111000000101110010: color_data = Z;
		19'b0111000000101110011: color_data = Z;
		19'b0111000000101110100: color_data = Z;
		19'b0111000000101110101: color_data = Z;
		19'b0111000000101110110: color_data = Z;
		19'b0111000000101110111: color_data = Z;
		19'b0111000000101111000: color_data = Z;
		19'b0111000000101111001: color_data = Z;
		19'b0111000000101111010: color_data = Z;
		19'b0111000000101111011: color_data = Z;
		19'b0111000000101111100: color_data = Z;
		19'b0111000000101111101: color_data = Z;
		19'b0111000000101111110: color_data = Z;
		19'b0111000000101111111: color_data = Z;
		19'b0111000000110000000: color_data = Z;
		19'b0111000000110000001: color_data = Z;
		19'b0111000000110000110: color_data = Z;
		19'b0111000000110000111: color_data = Z;
		19'b0111000000110001000: color_data = Z;
		19'b0111000000110001001: color_data = Z;
		19'b0111000000110001010: color_data = Z;
		19'b0111000000110001011: color_data = Z;
		19'b0111000000110001100: color_data = Z;
		19'b0111000000110001101: color_data = Z;
		19'b0111000000110001110: color_data = Z;
		19'b0111000000110001111: color_data = Z;
		19'b0111000000110010000: color_data = Z;
		19'b0111000000110010001: color_data = Z;
		19'b0111000000110010010: color_data = Z;
		19'b0111000000110010011: color_data = Z;
		19'b0111000000110010100: color_data = Z;
		19'b0111000000110010101: color_data = Z;
		19'b0111000000110010110: color_data = Z;
		19'b0111000000110010111: color_data = Z;
		19'b0111000000110011000: color_data = Z;
		19'b0111000000110011001: color_data = Z;
		19'b0111000000110011010: color_data = Z;
		19'b0111000000110011011: color_data = Z;
		19'b0111000000110011100: color_data = Z;
		19'b0111000000110011101: color_data = Z;
		19'b0111000000110011110: color_data = Z;
		19'b0111000000110011111: color_data = Z;
		19'b0111000000110100000: color_data = Z;
		19'b0111000000110100001: color_data = Z;
		19'b0111000000110100010: color_data = Z;
		19'b0111000000110100011: color_data = Z;
		19'b0111000000110110111: color_data = Z;
		19'b0111000000110111000: color_data = Z;
		19'b0111000000110111001: color_data = Z;
		19'b0111000000110111010: color_data = Z;
		19'b0111000000110111011: color_data = Z;
		19'b0111000000110111100: color_data = Z;
		19'b0111000000110111101: color_data = Z;
		19'b0111000000110111110: color_data = Z;
		19'b0111000000111010101: color_data = Z;
		19'b0111000000111010110: color_data = Z;
		19'b0111000000111010111: color_data = Z;
		19'b0111000010010101000: color_data = Z;
		19'b0111000010010101001: color_data = Z;
		19'b0111000010010101010: color_data = Z;
		19'b0111000010010101011: color_data = Z;
		19'b0111000010010101100: color_data = Z;
		19'b0111000010010101101: color_data = Z;
		19'b0111000010010101110: color_data = Z;
		19'b0111000010010101111: color_data = Z;
		19'b0111000010010110010: color_data = Z;
		19'b0111000010010110011: color_data = Z;
		19'b0111000010010110101: color_data = Z;
		19'b0111000010010110110: color_data = Z;
		19'b0111000010010110111: color_data = Z;
		19'b0111000010010111000: color_data = Z;
		19'b0111000010010111001: color_data = Z;
		19'b0111000010010111010: color_data = Z;
		19'b0111000010010111011: color_data = Z;
		19'b0111000010010111100: color_data = Z;
		19'b0111000010010111101: color_data = Z;
		19'b0111000010010111110: color_data = Z;
		19'b0111000010100010011: color_data = Z;
		19'b0111000010100010100: color_data = Z;
		19'b0111000010100010101: color_data = Z;
		19'b0111000010100011000: color_data = Z;
		19'b0111000010100011001: color_data = Z;
		19'b0111000010100011010: color_data = Z;
		19'b0111000010100011011: color_data = Z;
		19'b0111000010100011100: color_data = Z;
		19'b0111000010100011101: color_data = Z;
		19'b0111000010100011110: color_data = Z;
		19'b0111000010100011111: color_data = Z;
		19'b0111000010100100000: color_data = Z;
		19'b0111000010100100001: color_data = Z;
		19'b0111000010100100010: color_data = Z;
		19'b0111000010100100011: color_data = Z;
		19'b0111000010100100100: color_data = Z;
		19'b0111000010100100101: color_data = Z;
		19'b0111000010100100110: color_data = Z;
		19'b0111000010100100111: color_data = Z;
		19'b0111000010100101000: color_data = Z;
		19'b0111000010100101001: color_data = Z;
		19'b0111000010100101100: color_data = Z;
		19'b0111000010100101101: color_data = Z;
		19'b0111000010100101110: color_data = Z;
		19'b0111000010100101111: color_data = Z;
		19'b0111000010100110000: color_data = Z;
		19'b0111000010100110001: color_data = Z;
		19'b0111000010100110010: color_data = Z;
		19'b0111000010100110011: color_data = Z;
		19'b0111000010100110100: color_data = Z;
		19'b0111000010100110101: color_data = Z;
		19'b0111000010100110110: color_data = Z;
		19'b0111000010100110111: color_data = Z;
		19'b0111000010100111000: color_data = Z;
		19'b0111000010100111001: color_data = Z;
		19'b0111000010100111010: color_data = Z;
		19'b0111000010100111011: color_data = Z;
		19'b0111000010100111100: color_data = Z;
		19'b0111000010100111101: color_data = Z;
		19'b0111000010100111110: color_data = Z;
		19'b0111000010100111111: color_data = Z;
		19'b0111000010101000000: color_data = Z;
		19'b0111000010101000001: color_data = Z;
		19'b0111000010101000010: color_data = Z;
		19'b0111000010101000011: color_data = Z;
		19'b0111000010101000100: color_data = Z;
		19'b0111000010101000101: color_data = Z;
		19'b0111000010101000110: color_data = Z;
		19'b0111000010101000111: color_data = Z;
		19'b0111000010101001000: color_data = Z;
		19'b0111000010101001001: color_data = Z;
		19'b0111000010101001010: color_data = Z;
		19'b0111000010101001011: color_data = Z;
		19'b0111000010101001100: color_data = Z;
		19'b0111000010101001101: color_data = Z;
		19'b0111000010101001110: color_data = Z;
		19'b0111000010101001111: color_data = Z;
		19'b0111000010101010000: color_data = Z;
		19'b0111000010101010001: color_data = Z;
		19'b0111000010101010010: color_data = Z;
		19'b0111000010101010011: color_data = Z;
		19'b0111000010101010100: color_data = Z;
		19'b0111000010101010101: color_data = Z;
		19'b0111000010101010110: color_data = Z;
		19'b0111000010101010111: color_data = Z;
		19'b0111000010101011000: color_data = Z;
		19'b0111000010101011001: color_data = Z;
		19'b0111000010101011010: color_data = Z;
		19'b0111000010101011011: color_data = Z;
		19'b0111000010101011100: color_data = Z;
		19'b0111000010101011101: color_data = Z;
		19'b0111000010101011110: color_data = Z;
		19'b0111000010101011111: color_data = Z;
		19'b0111000010101100000: color_data = Z;
		19'b0111000010101100001: color_data = Z;
		19'b0111000010101100010: color_data = Z;
		19'b0111000010101100011: color_data = Z;
		19'b0111000010101100100: color_data = Z;
		19'b0111000010101100101: color_data = Z;
		19'b0111000010101100110: color_data = Z;
		19'b0111000010101100111: color_data = Z;
		19'b0111000010101101000: color_data = Z;
		19'b0111000010101101001: color_data = Z;
		19'b0111000010101101010: color_data = Z;
		19'b0111000010101101101: color_data = Z;
		19'b0111000010101101110: color_data = Z;
		19'b0111000010101101111: color_data = Z;
		19'b0111000010101110000: color_data = Z;
		19'b0111000010101110001: color_data = Z;
		19'b0111000010101110010: color_data = Z;
		19'b0111000010101110011: color_data = Z;
		19'b0111000010101110100: color_data = Z;
		19'b0111000010101110101: color_data = Z;
		19'b0111000010101110110: color_data = Z;
		19'b0111000010101110111: color_data = Z;
		19'b0111000010101111000: color_data = Z;
		19'b0111000010101111001: color_data = Z;
		19'b0111000010101111010: color_data = Z;
		19'b0111000010101111011: color_data = Z;
		19'b0111000010101111100: color_data = Z;
		19'b0111000010101111101: color_data = Z;
		19'b0111000010101111110: color_data = Z;
		19'b0111000010101111111: color_data = Z;
		19'b0111000010110000000: color_data = Z;
		19'b0111000010110000001: color_data = Z;
		19'b0111000010110000010: color_data = Z;
		19'b0111000010110000111: color_data = Z;
		19'b0111000010110001000: color_data = Z;
		19'b0111000010110001001: color_data = Z;
		19'b0111000010110001010: color_data = Z;
		19'b0111000010110001011: color_data = Z;
		19'b0111000010110001100: color_data = Z;
		19'b0111000010110001101: color_data = Z;
		19'b0111000010110001110: color_data = Z;
		19'b0111000010110001111: color_data = Z;
		19'b0111000010110010000: color_data = Z;
		19'b0111000010110010001: color_data = Z;
		19'b0111000010110010010: color_data = Z;
		19'b0111000010110010011: color_data = Z;
		19'b0111000010110010100: color_data = Z;
		19'b0111000010110010101: color_data = Z;
		19'b0111000010110010110: color_data = Z;
		19'b0111000010110010111: color_data = Z;
		19'b0111000010110011000: color_data = Z;
		19'b0111000010110011001: color_data = Z;
		19'b0111000010110011010: color_data = Z;
		19'b0111000010110011011: color_data = Z;
		19'b0111000010110011100: color_data = Z;
		19'b0111000010110011101: color_data = Z;
		19'b0111000010110011110: color_data = Z;
		19'b0111000010110011111: color_data = Z;
		19'b0111000010110100000: color_data = Z;
		19'b0111000010110100001: color_data = Z;
		19'b0111000010110100010: color_data = Z;
		19'b0111000010110100011: color_data = Z;
		19'b0111000010110100100: color_data = Z;
		19'b0111000010110100101: color_data = Z;
		19'b0111000010110100110: color_data = Z;
		19'b0111000010110110111: color_data = Z;
		19'b0111000010110111000: color_data = Z;
		19'b0111000010110111001: color_data = Z;
		19'b0111000010110111010: color_data = Z;
		19'b0111000010110111011: color_data = Z;
		19'b0111000010110111100: color_data = Z;
		19'b0111000010110111101: color_data = Z;
		19'b0111000010110111110: color_data = Z;
		19'b0111000010111010110: color_data = Z;
		19'b0111000010111010111: color_data = Z;
		19'b0111000100010101001: color_data = Z;
		19'b0111000100010101010: color_data = Z;
		19'b0111000100010101011: color_data = Z;
		19'b0111000100010101100: color_data = Z;
		19'b0111000100010101101: color_data = Z;
		19'b0111000100010101110: color_data = Z;
		19'b0111000100010101111: color_data = Z;
		19'b0111000100010110010: color_data = Z;
		19'b0111000100010110011: color_data = Z;
		19'b0111000100010110100: color_data = Z;
		19'b0111000100010110110: color_data = Z;
		19'b0111000100010110111: color_data = Z;
		19'b0111000100010111000: color_data = Z;
		19'b0111000100010111001: color_data = Z;
		19'b0111000100010111010: color_data = Z;
		19'b0111000100010111011: color_data = Z;
		19'b0111000100010111100: color_data = Z;
		19'b0111000100010111101: color_data = Z;
		19'b0111000100010111110: color_data = Z;
		19'b0111000100010111111: color_data = Z;
		19'b0111000100100010011: color_data = Z;
		19'b0111000100100010100: color_data = Z;
		19'b0111000100100010111: color_data = Z;
		19'b0111000100100011000: color_data = Z;
		19'b0111000100100011001: color_data = Z;
		19'b0111000100100011010: color_data = Z;
		19'b0111000100100011011: color_data = Z;
		19'b0111000100100011100: color_data = Z;
		19'b0111000100100011101: color_data = Z;
		19'b0111000100100011110: color_data = Z;
		19'b0111000100100011111: color_data = Z;
		19'b0111000100100100000: color_data = Z;
		19'b0111000100100100001: color_data = Z;
		19'b0111000100100100010: color_data = Z;
		19'b0111000100100100011: color_data = Z;
		19'b0111000100100100100: color_data = Z;
		19'b0111000100100100101: color_data = Z;
		19'b0111000100100100110: color_data = Z;
		19'b0111000100100100111: color_data = Z;
		19'b0111000100100101000: color_data = Z;
		19'b0111000100100101100: color_data = Z;
		19'b0111000100100101101: color_data = Z;
		19'b0111000100100101110: color_data = Z;
		19'b0111000100100101111: color_data = Z;
		19'b0111000100100110000: color_data = Z;
		19'b0111000100100110001: color_data = Z;
		19'b0111000100100110010: color_data = Z;
		19'b0111000100100110011: color_data = Z;
		19'b0111000100100110100: color_data = Z;
		19'b0111000100100110101: color_data = Z;
		19'b0111000100100110110: color_data = Z;
		19'b0111000100100110111: color_data = Z;
		19'b0111000100100111000: color_data = Z;
		19'b0111000100100111001: color_data = Z;
		19'b0111000100100111010: color_data = Z;
		19'b0111000100100111011: color_data = Z;
		19'b0111000100100111100: color_data = Z;
		19'b0111000100100111101: color_data = Z;
		19'b0111000100100111110: color_data = Z;
		19'b0111000100100111111: color_data = Z;
		19'b0111000100101000000: color_data = Z;
		19'b0111000100101000001: color_data = Z;
		19'b0111000100101000010: color_data = Z;
		19'b0111000100101000011: color_data = Z;
		19'b0111000100101000100: color_data = Z;
		19'b0111000100101000101: color_data = Z;
		19'b0111000100101000110: color_data = Z;
		19'b0111000100101000111: color_data = Z;
		19'b0111000100101001000: color_data = Z;
		19'b0111000100101001001: color_data = Z;
		19'b0111000100101001010: color_data = Z;
		19'b0111000100101001011: color_data = Z;
		19'b0111000100101001100: color_data = Z;
		19'b0111000100101001101: color_data = Z;
		19'b0111000100101001110: color_data = Z;
		19'b0111000100101001111: color_data = Z;
		19'b0111000100101010000: color_data = Z;
		19'b0111000100101010001: color_data = Z;
		19'b0111000100101010010: color_data = Z;
		19'b0111000100101010011: color_data = Z;
		19'b0111000100101010100: color_data = Z;
		19'b0111000100101010101: color_data = Z;
		19'b0111000100101010110: color_data = Z;
		19'b0111000100101010111: color_data = Z;
		19'b0111000100101011000: color_data = Z;
		19'b0111000100101011001: color_data = Z;
		19'b0111000100101011010: color_data = Z;
		19'b0111000100101011011: color_data = Z;
		19'b0111000100101011100: color_data = Z;
		19'b0111000100101011101: color_data = Z;
		19'b0111000100101011110: color_data = Z;
		19'b0111000100101011111: color_data = Z;
		19'b0111000100101100000: color_data = Z;
		19'b0111000100101100001: color_data = Z;
		19'b0111000100101100010: color_data = Z;
		19'b0111000100101100011: color_data = Z;
		19'b0111000100101100100: color_data = Z;
		19'b0111000100101100101: color_data = Z;
		19'b0111000100101100110: color_data = Z;
		19'b0111000100101100111: color_data = Z;
		19'b0111000100101101000: color_data = Z;
		19'b0111000100101101001: color_data = Z;
		19'b0111000100101101010: color_data = Z;
		19'b0111000100101101011: color_data = Z;
		19'b0111000100101101110: color_data = Z;
		19'b0111000100101101111: color_data = Z;
		19'b0111000100101110000: color_data = Z;
		19'b0111000100101110001: color_data = Z;
		19'b0111000100101110010: color_data = Z;
		19'b0111000100101110011: color_data = Z;
		19'b0111000100101110100: color_data = Z;
		19'b0111000100101110101: color_data = Z;
		19'b0111000100101110110: color_data = Z;
		19'b0111000100101110111: color_data = Z;
		19'b0111000100101111000: color_data = Z;
		19'b0111000100101111001: color_data = Z;
		19'b0111000100101111010: color_data = Z;
		19'b0111000100101111011: color_data = Z;
		19'b0111000100101111100: color_data = Z;
		19'b0111000100101111101: color_data = Z;
		19'b0111000100101111110: color_data = Z;
		19'b0111000100101111111: color_data = Z;
		19'b0111000100110000000: color_data = Z;
		19'b0111000100110000001: color_data = Z;
		19'b0111000100110000010: color_data = Z;
		19'b0111000100110000011: color_data = Z;
		19'b0111000100110001000: color_data = Z;
		19'b0111000100110001001: color_data = Z;
		19'b0111000100110001010: color_data = Z;
		19'b0111000100110001011: color_data = Z;
		19'b0111000100110001100: color_data = Z;
		19'b0111000100110001101: color_data = Z;
		19'b0111000100110001110: color_data = Z;
		19'b0111000100110001111: color_data = Z;
		19'b0111000100110010000: color_data = Z;
		19'b0111000100110010001: color_data = Z;
		19'b0111000100110010010: color_data = Z;
		19'b0111000100110010011: color_data = Z;
		19'b0111000100110010100: color_data = Z;
		19'b0111000100110010101: color_data = Z;
		19'b0111000100110010110: color_data = Z;
		19'b0111000100110010111: color_data = Z;
		19'b0111000100110011000: color_data = Z;
		19'b0111000100110011001: color_data = Z;
		19'b0111000100110011010: color_data = Z;
		19'b0111000100110011011: color_data = Z;
		19'b0111000100110011100: color_data = Z;
		19'b0111000100110011101: color_data = Z;
		19'b0111000100110011110: color_data = Z;
		19'b0111000100110011111: color_data = Z;
		19'b0111000100110100000: color_data = Z;
		19'b0111000100110100001: color_data = Z;
		19'b0111000100110100010: color_data = Z;
		19'b0111000100110100011: color_data = Z;
		19'b0111000100110100100: color_data = Z;
		19'b0111000100110100101: color_data = Z;
		19'b0111000100110100110: color_data = Z;
		19'b0111000100110100111: color_data = Z;
		19'b0111000100110101000: color_data = Z;
		19'b0111000100110110110: color_data = Z;
		19'b0111000100110110111: color_data = Z;
		19'b0111000100110111000: color_data = Z;
		19'b0111000100110111001: color_data = Z;
		19'b0111000100110111010: color_data = Z;
		19'b0111000100110111011: color_data = Z;
		19'b0111000100110111100: color_data = Z;
		19'b0111000100110111101: color_data = Z;
		19'b0111000100110111110: color_data = Z;
		19'b0111000110010101001: color_data = Z;
		19'b0111000110010101010: color_data = Z;
		19'b0111000110010101011: color_data = Z;
		19'b0111000110010101100: color_data = Z;
		19'b0111000110010101101: color_data = Z;
		19'b0111000110010101110: color_data = Z;
		19'b0111000110010101111: color_data = Z;
		19'b0111000110010110000: color_data = Z;
		19'b0111000110010110001: color_data = Z;
		19'b0111000110010110010: color_data = Z;
		19'b0111000110010110011: color_data = Z;
		19'b0111000110010110100: color_data = Z;
		19'b0111000110010110111: color_data = Z;
		19'b0111000110010111000: color_data = Z;
		19'b0111000110010111001: color_data = Z;
		19'b0111000110010111010: color_data = Z;
		19'b0111000110010111011: color_data = Z;
		19'b0111000110010111100: color_data = Z;
		19'b0111000110010111101: color_data = Z;
		19'b0111000110010111110: color_data = Z;
		19'b0111000110010111111: color_data = Z;
		19'b0111000110100010010: color_data = Z;
		19'b0111000110100010011: color_data = Z;
		19'b0111000110100010111: color_data = Z;
		19'b0111000110100011000: color_data = Z;
		19'b0111000110100011001: color_data = Z;
		19'b0111000110100011010: color_data = Z;
		19'b0111000110100011011: color_data = Z;
		19'b0111000110100011100: color_data = Z;
		19'b0111000110100011101: color_data = Z;
		19'b0111000110100011110: color_data = Z;
		19'b0111000110100011111: color_data = Z;
		19'b0111000110100100000: color_data = Z;
		19'b0111000110100100001: color_data = Z;
		19'b0111000110100100010: color_data = Z;
		19'b0111000110100100011: color_data = Z;
		19'b0111000110100100100: color_data = Z;
		19'b0111000110100100101: color_data = Z;
		19'b0111000110100100110: color_data = Z;
		19'b0111000110100100111: color_data = Z;
		19'b0111000110100101000: color_data = Z;
		19'b0111000110100101011: color_data = Z;
		19'b0111000110100101100: color_data = Z;
		19'b0111000110100101101: color_data = Z;
		19'b0111000110100101110: color_data = Z;
		19'b0111000110100101111: color_data = Z;
		19'b0111000110100110000: color_data = Z;
		19'b0111000110100110001: color_data = Z;
		19'b0111000110100110010: color_data = Z;
		19'b0111000110100110011: color_data = Z;
		19'b0111000110100110100: color_data = Z;
		19'b0111000110100110101: color_data = Z;
		19'b0111000110100110110: color_data = Z;
		19'b0111000110100110111: color_data = Z;
		19'b0111000110100111000: color_data = Z;
		19'b0111000110100111001: color_data = Z;
		19'b0111000110100111010: color_data = Z;
		19'b0111000110100111011: color_data = Z;
		19'b0111000110100111100: color_data = Z;
		19'b0111000110100111101: color_data = Z;
		19'b0111000110100111110: color_data = Z;
		19'b0111000110100111111: color_data = Z;
		19'b0111000110101000000: color_data = Z;
		19'b0111000110101000001: color_data = Z;
		19'b0111000110101000010: color_data = Z;
		19'b0111000110101000011: color_data = Z;
		19'b0111000110101000100: color_data = Z;
		19'b0111000110101000101: color_data = Z;
		19'b0111000110101000110: color_data = Z;
		19'b0111000110101000111: color_data = Z;
		19'b0111000110101001000: color_data = Z;
		19'b0111000110101001001: color_data = Z;
		19'b0111000110101001010: color_data = Z;
		19'b0111000110101001011: color_data = Z;
		19'b0111000110101001100: color_data = Z;
		19'b0111000110101001101: color_data = Z;
		19'b0111000110101001110: color_data = Z;
		19'b0111000110101001111: color_data = Z;
		19'b0111000110101010000: color_data = Z;
		19'b0111000110101010001: color_data = Z;
		19'b0111000110101010010: color_data = Z;
		19'b0111000110101010011: color_data = Z;
		19'b0111000110101010100: color_data = Z;
		19'b0111000110101010101: color_data = Z;
		19'b0111000110101010110: color_data = Z;
		19'b0111000110101010111: color_data = Z;
		19'b0111000110101011000: color_data = Z;
		19'b0111000110101011001: color_data = Z;
		19'b0111000110101011010: color_data = Z;
		19'b0111000110101011011: color_data = Z;
		19'b0111000110101011100: color_data = Z;
		19'b0111000110101011101: color_data = Z;
		19'b0111000110101011110: color_data = Z;
		19'b0111000110101011111: color_data = Z;
		19'b0111000110101100000: color_data = Z;
		19'b0111000110101100001: color_data = Z;
		19'b0111000110101100010: color_data = Z;
		19'b0111000110101100011: color_data = Z;
		19'b0111000110101100100: color_data = Z;
		19'b0111000110101100101: color_data = Z;
		19'b0111000110101100110: color_data = Z;
		19'b0111000110101100111: color_data = Z;
		19'b0111000110101101000: color_data = Z;
		19'b0111000110101101001: color_data = Z;
		19'b0111000110101101010: color_data = Z;
		19'b0111000110101101011: color_data = Z;
		19'b0111000110101101110: color_data = Z;
		19'b0111000110101101111: color_data = Z;
		19'b0111000110101110000: color_data = Z;
		19'b0111000110101110001: color_data = Z;
		19'b0111000110101110010: color_data = Z;
		19'b0111000110101110011: color_data = Z;
		19'b0111000110101110100: color_data = Z;
		19'b0111000110101110101: color_data = Z;
		19'b0111000110101110110: color_data = Z;
		19'b0111000110101110111: color_data = Z;
		19'b0111000110101111000: color_data = Z;
		19'b0111000110101111001: color_data = Z;
		19'b0111000110101111010: color_data = Z;
		19'b0111000110101111011: color_data = Z;
		19'b0111000110101111100: color_data = Z;
		19'b0111000110101111101: color_data = Z;
		19'b0111000110101111110: color_data = Z;
		19'b0111000110101111111: color_data = Z;
		19'b0111000110110000000: color_data = Z;
		19'b0111000110110000001: color_data = Z;
		19'b0111000110110000010: color_data = Z;
		19'b0111000110110000011: color_data = Z;
		19'b0111000110110000100: color_data = Z;
		19'b0111000110110001000: color_data = Z;
		19'b0111000110110001001: color_data = Z;
		19'b0111000110110001010: color_data = Z;
		19'b0111000110110001011: color_data = Z;
		19'b0111000110110001100: color_data = Z;
		19'b0111000110110001101: color_data = Z;
		19'b0111000110110001110: color_data = Z;
		19'b0111000110110001111: color_data = Z;
		19'b0111000110110010000: color_data = Z;
		19'b0111000110110010001: color_data = Z;
		19'b0111000110110010010: color_data = Z;
		19'b0111000110110010011: color_data = Z;
		19'b0111000110110010100: color_data = Z;
		19'b0111000110110010101: color_data = Z;
		19'b0111000110110010110: color_data = Z;
		19'b0111000110110010111: color_data = Z;
		19'b0111000110110011000: color_data = Z;
		19'b0111000110110011001: color_data = Z;
		19'b0111000110110011010: color_data = Z;
		19'b0111000110110011011: color_data = Z;
		19'b0111000110110011100: color_data = Z;
		19'b0111000110110011101: color_data = Z;
		19'b0111000110110011110: color_data = Z;
		19'b0111000110110011111: color_data = Z;
		19'b0111000110110100000: color_data = Z;
		19'b0111000110110100001: color_data = Z;
		19'b0111000110110100010: color_data = Z;
		19'b0111000110110100011: color_data = Z;
		19'b0111000110110100100: color_data = Z;
		19'b0111000110110100101: color_data = Z;
		19'b0111000110110100110: color_data = Z;
		19'b0111000110110100111: color_data = Z;
		19'b0111000110110101000: color_data = Z;
		19'b0111000110110101001: color_data = Z;
		19'b0111000110110110100: color_data = Z;
		19'b0111000110110110101: color_data = Z;
		19'b0111000110110110110: color_data = Z;
		19'b0111000110110110111: color_data = Z;
		19'b0111000110110111000: color_data = Z;
		19'b0111000110110111001: color_data = Z;
		19'b0111000110110111010: color_data = Z;
		19'b0111000110110111011: color_data = Z;
		19'b0111000110110111100: color_data = Z;
		19'b0111000110110111101: color_data = Z;
		19'b0111000110110111110: color_data = Z;
		19'b0111001000010101001: color_data = Z;
		19'b0111001000010101010: color_data = Z;
		19'b0111001000010101011: color_data = Z;
		19'b0111001000010101100: color_data = Z;
		19'b0111001000010101101: color_data = Z;
		19'b0111001000010101110: color_data = Z;
		19'b0111001000010101111: color_data = Z;
		19'b0111001000010110000: color_data = Z;
		19'b0111001000010110010: color_data = Z;
		19'b0111001000010110011: color_data = Z;
		19'b0111001000010110100: color_data = Z;
		19'b0111001000010110101: color_data = Z;
		19'b0111001000010111001: color_data = Z;
		19'b0111001000010111010: color_data = Z;
		19'b0111001000010111011: color_data = Z;
		19'b0111001000010111100: color_data = Z;
		19'b0111001000010111101: color_data = Z;
		19'b0111001000010111110: color_data = Z;
		19'b0111001000010111111: color_data = Z;
		19'b0111001000011000000: color_data = Z;
		19'b0111001000100010111: color_data = Z;
		19'b0111001000100011000: color_data = Z;
		19'b0111001000100011001: color_data = Z;
		19'b0111001000100011010: color_data = Z;
		19'b0111001000100011011: color_data = Z;
		19'b0111001000100011100: color_data = Z;
		19'b0111001000100011101: color_data = Z;
		19'b0111001000100011110: color_data = Z;
		19'b0111001000100011111: color_data = Z;
		19'b0111001000100100000: color_data = Z;
		19'b0111001000100100001: color_data = Z;
		19'b0111001000100100010: color_data = Z;
		19'b0111001000100100011: color_data = Z;
		19'b0111001000100100100: color_data = Z;
		19'b0111001000100100101: color_data = Z;
		19'b0111001000100100110: color_data = Z;
		19'b0111001000100100111: color_data = Z;
		19'b0111001000100101011: color_data = Z;
		19'b0111001000100101100: color_data = Z;
		19'b0111001000100101101: color_data = Z;
		19'b0111001000100101110: color_data = Z;
		19'b0111001000100101111: color_data = Z;
		19'b0111001000100110000: color_data = Z;
		19'b0111001000100110001: color_data = Z;
		19'b0111001000100110010: color_data = Z;
		19'b0111001000100110011: color_data = Z;
		19'b0111001000100110100: color_data = Z;
		19'b0111001000100110101: color_data = Z;
		19'b0111001000100110110: color_data = Z;
		19'b0111001000100110111: color_data = Z;
		19'b0111001000100111000: color_data = Z;
		19'b0111001000100111001: color_data = Z;
		19'b0111001000100111010: color_data = Z;
		19'b0111001000100111100: color_data = Z;
		19'b0111001000100111101: color_data = Z;
		19'b0111001000100111110: color_data = Z;
		19'b0111001000100111111: color_data = Z;
		19'b0111001000101000000: color_data = Z;
		19'b0111001000101000001: color_data = Z;
		19'b0111001000101000010: color_data = Z;
		19'b0111001000101000011: color_data = Z;
		19'b0111001000101000100: color_data = Z;
		19'b0111001000101000101: color_data = Z;
		19'b0111001000101000110: color_data = Z;
		19'b0111001000101000111: color_data = Z;
		19'b0111001000101001000: color_data = Z;
		19'b0111001000101001001: color_data = Z;
		19'b0111001000101001010: color_data = Z;
		19'b0111001000101001011: color_data = Z;
		19'b0111001000101001100: color_data = Z;
		19'b0111001000101001101: color_data = Z;
		19'b0111001000101001110: color_data = Z;
		19'b0111001000101001111: color_data = Z;
		19'b0111001000101010000: color_data = Z;
		19'b0111001000101010001: color_data = Z;
		19'b0111001000101010010: color_data = Z;
		19'b0111001000101010011: color_data = Z;
		19'b0111001000101010100: color_data = Z;
		19'b0111001000101010101: color_data = Z;
		19'b0111001000101010110: color_data = Z;
		19'b0111001000101010111: color_data = Z;
		19'b0111001000101011000: color_data = Z;
		19'b0111001000101011001: color_data = Z;
		19'b0111001000101011010: color_data = Z;
		19'b0111001000101011011: color_data = Z;
		19'b0111001000101011100: color_data = Z;
		19'b0111001000101011101: color_data = Z;
		19'b0111001000101011110: color_data = Z;
		19'b0111001000101011111: color_data = Z;
		19'b0111001000101100000: color_data = Z;
		19'b0111001000101100001: color_data = Z;
		19'b0111001000101100010: color_data = Z;
		19'b0111001000101100011: color_data = Z;
		19'b0111001000101100100: color_data = Z;
		19'b0111001000101100101: color_data = Z;
		19'b0111001000101100110: color_data = Z;
		19'b0111001000101100111: color_data = Z;
		19'b0111001000101101000: color_data = Z;
		19'b0111001000101101001: color_data = Z;
		19'b0111001000101101010: color_data = Z;
		19'b0111001000101101011: color_data = Z;
		19'b0111001000101101111: color_data = Z;
		19'b0111001000101110000: color_data = Z;
		19'b0111001000101110001: color_data = Z;
		19'b0111001000101110010: color_data = Z;
		19'b0111001000101110011: color_data = Z;
		19'b0111001000101110100: color_data = Z;
		19'b0111001000101110101: color_data = Z;
		19'b0111001000101110110: color_data = Z;
		19'b0111001000101110111: color_data = Z;
		19'b0111001000101111000: color_data = Z;
		19'b0111001000101111001: color_data = Z;
		19'b0111001000101111010: color_data = Z;
		19'b0111001000101111011: color_data = Z;
		19'b0111001000101111100: color_data = Z;
		19'b0111001000101111101: color_data = Z;
		19'b0111001000101111110: color_data = Z;
		19'b0111001000101111111: color_data = Z;
		19'b0111001000110000000: color_data = Z;
		19'b0111001000110000001: color_data = Z;
		19'b0111001000110000010: color_data = Z;
		19'b0111001000110000011: color_data = Z;
		19'b0111001000110000100: color_data = Z;
		19'b0111001000110001001: color_data = Z;
		19'b0111001000110001010: color_data = Z;
		19'b0111001000110001011: color_data = Z;
		19'b0111001000110001100: color_data = Z;
		19'b0111001000110001101: color_data = Z;
		19'b0111001000110001110: color_data = Z;
		19'b0111001000110001111: color_data = Z;
		19'b0111001000110010000: color_data = Z;
		19'b0111001000110010001: color_data = Z;
		19'b0111001000110010010: color_data = Z;
		19'b0111001000110010011: color_data = Z;
		19'b0111001000110010100: color_data = Z;
		19'b0111001000110010101: color_data = Z;
		19'b0111001000110010110: color_data = Z;
		19'b0111001000110010111: color_data = Z;
		19'b0111001000110011000: color_data = Z;
		19'b0111001000110011001: color_data = Z;
		19'b0111001000110011010: color_data = Z;
		19'b0111001000110011011: color_data = Z;
		19'b0111001000110011100: color_data = Z;
		19'b0111001000110011101: color_data = Z;
		19'b0111001000110011110: color_data = Z;
		19'b0111001000110011111: color_data = Z;
		19'b0111001000110100000: color_data = Z;
		19'b0111001000110100001: color_data = Z;
		19'b0111001000110100010: color_data = Z;
		19'b0111001000110100011: color_data = Z;
		19'b0111001000110100100: color_data = Z;
		19'b0111001000110100101: color_data = Z;
		19'b0111001000110100110: color_data = Z;
		19'b0111001000110100111: color_data = Z;
		19'b0111001000110101000: color_data = Z;
		19'b0111001000110101001: color_data = Z;
		19'b0111001000110101010: color_data = Z;
		19'b0111001000110101011: color_data = Z;
		19'b0111001000110101100: color_data = Z;
		19'b0111001000110101101: color_data = Z;
		19'b0111001000110110100: color_data = Z;
		19'b0111001000110110101: color_data = Z;
		19'b0111001000110110110: color_data = Z;
		19'b0111001000110110111: color_data = Z;
		19'b0111001000110111000: color_data = Z;
		19'b0111001000110111001: color_data = Z;
		19'b0111001000110111010: color_data = Z;
		19'b0111001000110111011: color_data = Z;
		19'b0111001000110111100: color_data = Z;
		19'b0111001000110111101: color_data = Z;
		19'b0111001000110111110: color_data = Z;
		19'b0111001010010101010: color_data = Z;
		19'b0111001010010101011: color_data = Z;
		19'b0111001010010101100: color_data = Z;
		19'b0111001010010101101: color_data = Z;
		19'b0111001010010101110: color_data = Z;
		19'b0111001010010101111: color_data = Z;
		19'b0111001010010110000: color_data = Z;
		19'b0111001010010110001: color_data = Z;
		19'b0111001010010110010: color_data = Z;
		19'b0111001010010110011: color_data = Z;
		19'b0111001010010110100: color_data = Z;
		19'b0111001010010110101: color_data = Z;
		19'b0111001010010111010: color_data = Z;
		19'b0111001010010111011: color_data = Z;
		19'b0111001010010111100: color_data = Z;
		19'b0111001010010111101: color_data = Z;
		19'b0111001010010111110: color_data = Z;
		19'b0111001010010111111: color_data = Z;
		19'b0111001010011000000: color_data = Z;
		19'b0111001010100010110: color_data = Z;
		19'b0111001010100010111: color_data = Z;
		19'b0111001010100011000: color_data = Z;
		19'b0111001010100011001: color_data = Z;
		19'b0111001010100011010: color_data = Z;
		19'b0111001010100011011: color_data = Z;
		19'b0111001010100011100: color_data = Z;
		19'b0111001010100011101: color_data = Z;
		19'b0111001010100011110: color_data = Z;
		19'b0111001010100011111: color_data = Z;
		19'b0111001010100100000: color_data = Z;
		19'b0111001010100100001: color_data = Z;
		19'b0111001010100100010: color_data = Z;
		19'b0111001010100100011: color_data = Z;
		19'b0111001010100100100: color_data = Z;
		19'b0111001010100100101: color_data = Z;
		19'b0111001010100100110: color_data = Z;
		19'b0111001010100100111: color_data = Z;
		19'b0111001010100101011: color_data = Z;
		19'b0111001010100101100: color_data = Z;
		19'b0111001010100101101: color_data = Z;
		19'b0111001010100101110: color_data = Z;
		19'b0111001010100101111: color_data = Z;
		19'b0111001010100110000: color_data = Z;
		19'b0111001010100110001: color_data = Z;
		19'b0111001010100110010: color_data = Z;
		19'b0111001010100110011: color_data = Z;
		19'b0111001010100110100: color_data = Z;
		19'b0111001010100110101: color_data = Z;
		19'b0111001010100110110: color_data = Z;
		19'b0111001010100110111: color_data = Z;
		19'b0111001010100111000: color_data = Z;
		19'b0111001010100111001: color_data = Z;
		19'b0111001010100111010: color_data = Z;
		19'b0111001010100111100: color_data = Z;
		19'b0111001010100111101: color_data = Z;
		19'b0111001010100111110: color_data = Z;
		19'b0111001010100111111: color_data = Z;
		19'b0111001010101000000: color_data = Z;
		19'b0111001010101000001: color_data = Z;
		19'b0111001010101000010: color_data = Z;
		19'b0111001010101000011: color_data = Z;
		19'b0111001010101000100: color_data = Z;
		19'b0111001010101000101: color_data = Z;
		19'b0111001010101000110: color_data = Z;
		19'b0111001010101000111: color_data = Z;
		19'b0111001010101001000: color_data = Z;
		19'b0111001010101001001: color_data = Z;
		19'b0111001010101001010: color_data = Z;
		19'b0111001010101001011: color_data = Z;
		19'b0111001010101001100: color_data = Z;
		19'b0111001010101001101: color_data = Z;
		19'b0111001010101001110: color_data = Z;
		19'b0111001010101001111: color_data = Z;
		19'b0111001010101010000: color_data = Z;
		19'b0111001010101010001: color_data = Z;
		19'b0111001010101010010: color_data = Z;
		19'b0111001010101010011: color_data = Z;
		19'b0111001010101010100: color_data = Z;
		19'b0111001010101010101: color_data = Z;
		19'b0111001010101010110: color_data = Z;
		19'b0111001010101010111: color_data = Z;
		19'b0111001010101011000: color_data = Z;
		19'b0111001010101011001: color_data = Z;
		19'b0111001010101011010: color_data = Z;
		19'b0111001010101011011: color_data = Z;
		19'b0111001010101011100: color_data = Z;
		19'b0111001010101011101: color_data = Z;
		19'b0111001010101011110: color_data = Z;
		19'b0111001010101011111: color_data = Z;
		19'b0111001010101100000: color_data = Z;
		19'b0111001010101100001: color_data = Z;
		19'b0111001010101100010: color_data = Z;
		19'b0111001010101100011: color_data = Z;
		19'b0111001010101100100: color_data = Z;
		19'b0111001010101100101: color_data = Z;
		19'b0111001010101100110: color_data = Z;
		19'b0111001010101100111: color_data = Z;
		19'b0111001010101101000: color_data = Z;
		19'b0111001010101101001: color_data = Z;
		19'b0111001010101101010: color_data = Z;
		19'b0111001010101101011: color_data = Z;
		19'b0111001010101101111: color_data = Z;
		19'b0111001010101110000: color_data = Z;
		19'b0111001010101110001: color_data = Z;
		19'b0111001010101110010: color_data = Z;
		19'b0111001010101110011: color_data = Z;
		19'b0111001010101110100: color_data = Z;
		19'b0111001010101110101: color_data = Z;
		19'b0111001010101110110: color_data = Z;
		19'b0111001010101110111: color_data = Z;
		19'b0111001010101111000: color_data = Z;
		19'b0111001010101111001: color_data = Z;
		19'b0111001010101111010: color_data = Z;
		19'b0111001010101111011: color_data = Z;
		19'b0111001010101111100: color_data = Z;
		19'b0111001010101111101: color_data = Z;
		19'b0111001010101111110: color_data = Z;
		19'b0111001010101111111: color_data = Z;
		19'b0111001010110000000: color_data = Z;
		19'b0111001010110000001: color_data = Z;
		19'b0111001010110000010: color_data = Z;
		19'b0111001010110000011: color_data = Z;
		19'b0111001010110000100: color_data = Z;
		19'b0111001010110000101: color_data = Z;
		19'b0111001010110001010: color_data = Z;
		19'b0111001010110001011: color_data = Z;
		19'b0111001010110001100: color_data = Z;
		19'b0111001010110001101: color_data = Z;
		19'b0111001010110001110: color_data = Z;
		19'b0111001010110001111: color_data = Z;
		19'b0111001010110010000: color_data = Z;
		19'b0111001010110010001: color_data = Z;
		19'b0111001010110010010: color_data = Z;
		19'b0111001010110010011: color_data = Z;
		19'b0111001010110010100: color_data = Z;
		19'b0111001010110010101: color_data = Z;
		19'b0111001010110010110: color_data = Z;
		19'b0111001010110010111: color_data = Z;
		19'b0111001010110011000: color_data = Z;
		19'b0111001010110011001: color_data = Z;
		19'b0111001010110011010: color_data = Z;
		19'b0111001010110011011: color_data = Z;
		19'b0111001010110011100: color_data = Z;
		19'b0111001010110011101: color_data = Z;
		19'b0111001010110011110: color_data = Z;
		19'b0111001010110011111: color_data = Z;
		19'b0111001010110100000: color_data = Z;
		19'b0111001010110100001: color_data = Z;
		19'b0111001010110100010: color_data = Z;
		19'b0111001010110100011: color_data = Z;
		19'b0111001010110100100: color_data = Z;
		19'b0111001010110100101: color_data = Z;
		19'b0111001010110100110: color_data = Z;
		19'b0111001010110100111: color_data = Z;
		19'b0111001010110101000: color_data = Z;
		19'b0111001010110101001: color_data = Z;
		19'b0111001010110101010: color_data = Z;
		19'b0111001010110101011: color_data = Z;
		19'b0111001010110101100: color_data = Z;
		19'b0111001010110101101: color_data = Z;
		19'b0111001010110101110: color_data = Z;
		19'b0111001010110101111: color_data = Z;
		19'b0111001010110110100: color_data = Z;
		19'b0111001010110110101: color_data = Z;
		19'b0111001010110110110: color_data = Z;
		19'b0111001010110110111: color_data = Z;
		19'b0111001010110111000: color_data = Z;
		19'b0111001010110111001: color_data = Z;
		19'b0111001010110111010: color_data = Z;
		19'b0111001010110111011: color_data = Z;
		19'b0111001010110111100: color_data = Z;
		19'b0111001010110111101: color_data = Z;
		19'b0111001010110111110: color_data = Z;
		19'b0111001100010101010: color_data = Z;
		19'b0111001100010101011: color_data = Z;
		19'b0111001100010101100: color_data = Z;
		19'b0111001100010101101: color_data = Z;
		19'b0111001100010101110: color_data = Z;
		19'b0111001100010101111: color_data = Z;
		19'b0111001100010110000: color_data = Z;
		19'b0111001100010110001: color_data = Z;
		19'b0111001100010110010: color_data = Z;
		19'b0111001100010110011: color_data = Z;
		19'b0111001100010110100: color_data = Z;
		19'b0111001100010110101: color_data = Z;
		19'b0111001100010110110: color_data = Z;
		19'b0111001100010111011: color_data = Z;
		19'b0111001100010111100: color_data = Z;
		19'b0111001100010111101: color_data = Z;
		19'b0111001100010111110: color_data = Z;
		19'b0111001100010111111: color_data = Z;
		19'b0111001100011000000: color_data = Z;
		19'b0111001100011000001: color_data = Z;
		19'b0111001100100010110: color_data = Z;
		19'b0111001100100010111: color_data = Z;
		19'b0111001100100011000: color_data = Z;
		19'b0111001100100011001: color_data = Z;
		19'b0111001100100011010: color_data = Z;
		19'b0111001100100011011: color_data = Z;
		19'b0111001100100011100: color_data = Z;
		19'b0111001100100011101: color_data = Z;
		19'b0111001100100011110: color_data = Z;
		19'b0111001100100011111: color_data = Z;
		19'b0111001100100100000: color_data = Z;
		19'b0111001100100100001: color_data = Z;
		19'b0111001100100100010: color_data = Z;
		19'b0111001100100100011: color_data = Z;
		19'b0111001100100100100: color_data = Z;
		19'b0111001100100100101: color_data = Z;
		19'b0111001100100100110: color_data = Z;
		19'b0111001100100100111: color_data = Z;
		19'b0111001100100101000: color_data = Z;
		19'b0111001100100101010: color_data = Z;
		19'b0111001100100101011: color_data = Z;
		19'b0111001100100101100: color_data = Z;
		19'b0111001100100101101: color_data = Z;
		19'b0111001100100101110: color_data = Z;
		19'b0111001100100101111: color_data = Z;
		19'b0111001100100110000: color_data = Z;
		19'b0111001100100110001: color_data = Z;
		19'b0111001100100110010: color_data = Z;
		19'b0111001100100110011: color_data = Z;
		19'b0111001100100110100: color_data = Z;
		19'b0111001100100110101: color_data = Z;
		19'b0111001100100110110: color_data = Z;
		19'b0111001100100110111: color_data = Z;
		19'b0111001100100111000: color_data = Z;
		19'b0111001100100111001: color_data = Z;
		19'b0111001100100111100: color_data = Z;
		19'b0111001100100111101: color_data = Z;
		19'b0111001100100111110: color_data = Z;
		19'b0111001100100111111: color_data = Z;
		19'b0111001100101000000: color_data = Z;
		19'b0111001100101000001: color_data = Z;
		19'b0111001100101000010: color_data = Z;
		19'b0111001100101000011: color_data = Z;
		19'b0111001100101000100: color_data = Z;
		19'b0111001100101000101: color_data = Z;
		19'b0111001100101000110: color_data = Z;
		19'b0111001100101000111: color_data = Z;
		19'b0111001100101001000: color_data = Z;
		19'b0111001100101001001: color_data = Z;
		19'b0111001100101001010: color_data = Z;
		19'b0111001100101001011: color_data = Z;
		19'b0111001100101001100: color_data = Z;
		19'b0111001100101001101: color_data = Z;
		19'b0111001100101001110: color_data = Z;
		19'b0111001100101001111: color_data = Z;
		19'b0111001100101010000: color_data = Z;
		19'b0111001100101010001: color_data = Z;
		19'b0111001100101010010: color_data = Z;
		19'b0111001100101010011: color_data = Z;
		19'b0111001100101010100: color_data = Z;
		19'b0111001100101010101: color_data = Z;
		19'b0111001100101010110: color_data = Z;
		19'b0111001100101010111: color_data = Z;
		19'b0111001100101011000: color_data = Z;
		19'b0111001100101011001: color_data = Z;
		19'b0111001100101011010: color_data = Z;
		19'b0111001100101011011: color_data = Z;
		19'b0111001100101011100: color_data = Z;
		19'b0111001100101011101: color_data = Z;
		19'b0111001100101011110: color_data = Z;
		19'b0111001100101011111: color_data = Z;
		19'b0111001100101100000: color_data = Z;
		19'b0111001100101100001: color_data = Z;
		19'b0111001100101100010: color_data = Z;
		19'b0111001100101100011: color_data = Z;
		19'b0111001100101100100: color_data = Z;
		19'b0111001100101100101: color_data = Z;
		19'b0111001100101100110: color_data = Z;
		19'b0111001100101100111: color_data = Z;
		19'b0111001100101101000: color_data = Z;
		19'b0111001100101101001: color_data = Z;
		19'b0111001100101101010: color_data = Z;
		19'b0111001100101101011: color_data = Z;
		19'b0111001100101101100: color_data = Z;
		19'b0111001100101101101: color_data = Z;
		19'b0111001100101101111: color_data = Z;
		19'b0111001100101110000: color_data = Z;
		19'b0111001100101110001: color_data = Z;
		19'b0111001100101110010: color_data = Z;
		19'b0111001100101110011: color_data = Z;
		19'b0111001100101110100: color_data = Z;
		19'b0111001100101110101: color_data = Z;
		19'b0111001100101110110: color_data = Z;
		19'b0111001100101110111: color_data = Z;
		19'b0111001100101111000: color_data = Z;
		19'b0111001100101111001: color_data = Z;
		19'b0111001100101111010: color_data = Z;
		19'b0111001100101111011: color_data = Z;
		19'b0111001100101111100: color_data = Z;
		19'b0111001100101111101: color_data = Z;
		19'b0111001100101111110: color_data = Z;
		19'b0111001100101111111: color_data = Z;
		19'b0111001100110000000: color_data = Z;
		19'b0111001100110000001: color_data = Z;
		19'b0111001100110000010: color_data = Z;
		19'b0111001100110000011: color_data = Z;
		19'b0111001100110000100: color_data = Z;
		19'b0111001100110000101: color_data = Z;
		19'b0111001100110001010: color_data = Z;
		19'b0111001100110001011: color_data = Z;
		19'b0111001100110001100: color_data = Z;
		19'b0111001100110001101: color_data = Z;
		19'b0111001100110001110: color_data = Z;
		19'b0111001100110001111: color_data = Z;
		19'b0111001100110010000: color_data = Z;
		19'b0111001100110010001: color_data = Z;
		19'b0111001100110010010: color_data = Z;
		19'b0111001100110010011: color_data = Z;
		19'b0111001100110010100: color_data = Z;
		19'b0111001100110010111: color_data = Z;
		19'b0111001100110011000: color_data = Z;
		19'b0111001100110011001: color_data = Z;
		19'b0111001100110011010: color_data = Z;
		19'b0111001100110011011: color_data = Z;
		19'b0111001100110011100: color_data = Z;
		19'b0111001100110011101: color_data = Z;
		19'b0111001100110011110: color_data = Z;
		19'b0111001100110011111: color_data = Z;
		19'b0111001100110100000: color_data = Z;
		19'b0111001100110100001: color_data = Z;
		19'b0111001100110100010: color_data = Z;
		19'b0111001100110100011: color_data = Z;
		19'b0111001100110100100: color_data = Z;
		19'b0111001100110100101: color_data = Z;
		19'b0111001100110100110: color_data = Z;
		19'b0111001100110100111: color_data = Z;
		19'b0111001100110101000: color_data = Z;
		19'b0111001100110101001: color_data = Z;
		19'b0111001100110101010: color_data = Z;
		19'b0111001100110101011: color_data = Z;
		19'b0111001100110101100: color_data = Z;
		19'b0111001100110101101: color_data = Z;
		19'b0111001100110101110: color_data = Z;
		19'b0111001100110101111: color_data = Z;
		19'b0111001100110110011: color_data = Z;
		19'b0111001100110110100: color_data = Z;
		19'b0111001100110110101: color_data = Z;
		19'b0111001100110110110: color_data = Z;
		19'b0111001100110110111: color_data = Z;
		19'b0111001100110111000: color_data = Z;
		19'b0111001100110111001: color_data = Z;
		19'b0111001100110111010: color_data = Z;
		19'b0111001100110111011: color_data = Z;
		19'b0111001100110111100: color_data = Z;
		19'b0111001100110111101: color_data = Z;
		19'b0111001110010101010: color_data = Z;
		19'b0111001110010101011: color_data = Z;
		19'b0111001110010101100: color_data = Z;
		19'b0111001110010101101: color_data = Z;
		19'b0111001110010101110: color_data = Z;
		19'b0111001110010101111: color_data = Z;
		19'b0111001110010110000: color_data = Z;
		19'b0111001110010110001: color_data = Z;
		19'b0111001110010110010: color_data = Z;
		19'b0111001110010110011: color_data = Z;
		19'b0111001110010110100: color_data = Z;
		19'b0111001110010110101: color_data = Z;
		19'b0111001110010110110: color_data = Z;
		19'b0111001110010110111: color_data = Z;
		19'b0111001110010111100: color_data = Z;
		19'b0111001110010111101: color_data = Z;
		19'b0111001110010111110: color_data = Z;
		19'b0111001110010111111: color_data = Z;
		19'b0111001110011000000: color_data = Z;
		19'b0111001110011000001: color_data = Z;
		19'b0111001110011000010: color_data = Z;
		19'b0111001110100001101: color_data = Z;
		19'b0111001110100001110: color_data = Z;
		19'b0111001110100010101: color_data = Z;
		19'b0111001110100010110: color_data = Z;
		19'b0111001110100010111: color_data = Z;
		19'b0111001110100011011: color_data = Z;
		19'b0111001110100011100: color_data = Z;
		19'b0111001110100011101: color_data = Z;
		19'b0111001110100011110: color_data = Z;
		19'b0111001110100011111: color_data = Z;
		19'b0111001110100100000: color_data = Z;
		19'b0111001110100100001: color_data = Z;
		19'b0111001110100100010: color_data = Z;
		19'b0111001110100100011: color_data = Z;
		19'b0111001110100100100: color_data = Z;
		19'b0111001110100100101: color_data = Z;
		19'b0111001110100100110: color_data = Z;
		19'b0111001110100100111: color_data = Z;
		19'b0111001110100101000: color_data = Z;
		19'b0111001110100101010: color_data = Z;
		19'b0111001110100101011: color_data = Z;
		19'b0111001110100101100: color_data = Z;
		19'b0111001110100101101: color_data = Z;
		19'b0111001110100101110: color_data = Z;
		19'b0111001110100101111: color_data = Z;
		19'b0111001110100110000: color_data = Z;
		19'b0111001110100110001: color_data = Z;
		19'b0111001110100110010: color_data = Z;
		19'b0111001110100110011: color_data = Z;
		19'b0111001110100110100: color_data = Z;
		19'b0111001110100110101: color_data = Z;
		19'b0111001110100110110: color_data = Z;
		19'b0111001110100110111: color_data = Z;
		19'b0111001110100111000: color_data = Z;
		19'b0111001110100111001: color_data = Z;
		19'b0111001110100111100: color_data = Z;
		19'b0111001110100111101: color_data = Z;
		19'b0111001110100111110: color_data = Z;
		19'b0111001110100111111: color_data = Z;
		19'b0111001110101000000: color_data = Z;
		19'b0111001110101000001: color_data = Z;
		19'b0111001110101000010: color_data = Z;
		19'b0111001110101000011: color_data = Z;
		19'b0111001110101000100: color_data = Z;
		19'b0111001110101000101: color_data = Z;
		19'b0111001110101000110: color_data = Z;
		19'b0111001110101000111: color_data = Z;
		19'b0111001110101001000: color_data = Z;
		19'b0111001110101001001: color_data = Z;
		19'b0111001110101001010: color_data = Z;
		19'b0111001110101001011: color_data = Z;
		19'b0111001110101001100: color_data = Z;
		19'b0111001110101001101: color_data = Z;
		19'b0111001110101001110: color_data = Z;
		19'b0111001110101001111: color_data = Z;
		19'b0111001110101010000: color_data = Z;
		19'b0111001110101010001: color_data = Z;
		19'b0111001110101010010: color_data = Z;
		19'b0111001110101010011: color_data = Z;
		19'b0111001110101010100: color_data = Z;
		19'b0111001110101010101: color_data = Z;
		19'b0111001110101010110: color_data = Z;
		19'b0111001110101010111: color_data = Z;
		19'b0111001110101011000: color_data = Z;
		19'b0111001110101011001: color_data = Z;
		19'b0111001110101011010: color_data = Z;
		19'b0111001110101011011: color_data = Z;
		19'b0111001110101011100: color_data = Z;
		19'b0111001110101011101: color_data = Z;
		19'b0111001110101011110: color_data = Z;
		19'b0111001110101011111: color_data = Z;
		19'b0111001110101100000: color_data = Z;
		19'b0111001110101100001: color_data = Z;
		19'b0111001110101100010: color_data = Z;
		19'b0111001110101100011: color_data = Z;
		19'b0111001110101100100: color_data = Z;
		19'b0111001110101100101: color_data = Z;
		19'b0111001110101100110: color_data = Z;
		19'b0111001110101100111: color_data = Z;
		19'b0111001110101101000: color_data = Z;
		19'b0111001110101101001: color_data = Z;
		19'b0111001110101101010: color_data = Z;
		19'b0111001110101101011: color_data = Z;
		19'b0111001110101101100: color_data = Z;
		19'b0111001110101101101: color_data = Z;
		19'b0111001110101110000: color_data = Z;
		19'b0111001110101110001: color_data = Z;
		19'b0111001110101110010: color_data = Z;
		19'b0111001110101110011: color_data = Z;
		19'b0111001110101110100: color_data = Z;
		19'b0111001110101110101: color_data = Z;
		19'b0111001110101110110: color_data = Z;
		19'b0111001110101110111: color_data = Z;
		19'b0111001110101111000: color_data = Z;
		19'b0111001110101111001: color_data = Z;
		19'b0111001110101111010: color_data = Z;
		19'b0111001110101111011: color_data = Z;
		19'b0111001110101111100: color_data = Z;
		19'b0111001110101111101: color_data = Z;
		19'b0111001110101111110: color_data = Z;
		19'b0111001110101111111: color_data = Z;
		19'b0111001110110000000: color_data = Z;
		19'b0111001110110000001: color_data = Z;
		19'b0111001110110000010: color_data = Z;
		19'b0111001110110000011: color_data = Z;
		19'b0111001110110000100: color_data = Z;
		19'b0111001110110000101: color_data = Z;
		19'b0111001110110000110: color_data = Z;
		19'b0111001110110000111: color_data = Z;
		19'b0111001110110001011: color_data = Z;
		19'b0111001110110001100: color_data = Z;
		19'b0111001110110001101: color_data = Z;
		19'b0111001110110001110: color_data = Z;
		19'b0111001110110001111: color_data = Z;
		19'b0111001110110010000: color_data = Z;
		19'b0111001110110010010: color_data = Z;
		19'b0111001110110010011: color_data = Z;
		19'b0111001110110010100: color_data = Z;
		19'b0111001110110010101: color_data = Z;
		19'b0111001110110011000: color_data = Z;
		19'b0111001110110011001: color_data = Z;
		19'b0111001110110011010: color_data = Z;
		19'b0111001110110011011: color_data = Z;
		19'b0111001110110011100: color_data = Z;
		19'b0111001110110011101: color_data = Z;
		19'b0111001110110011110: color_data = Z;
		19'b0111001110110011111: color_data = Z;
		19'b0111001110110100000: color_data = Z;
		19'b0111001110110100001: color_data = Z;
		19'b0111001110110100010: color_data = Z;
		19'b0111001110110100011: color_data = Z;
		19'b0111001110110100100: color_data = Z;
		19'b0111001110110100101: color_data = Z;
		19'b0111001110110100110: color_data = Z;
		19'b0111001110110100111: color_data = Z;
		19'b0111001110110101000: color_data = Z;
		19'b0111001110110101001: color_data = Z;
		19'b0111001110110101010: color_data = Z;
		19'b0111001110110101011: color_data = Z;
		19'b0111001110110101100: color_data = Z;
		19'b0111001110110101101: color_data = Z;
		19'b0111001110110110011: color_data = Z;
		19'b0111001110110110100: color_data = Z;
		19'b0111001110110110101: color_data = Z;
		19'b0111001110110110110: color_data = Z;
		19'b0111001110110110111: color_data = Z;
		19'b0111001110110111000: color_data = Z;
		19'b0111001110110111001: color_data = Z;
		19'b0111001110110111010: color_data = Z;
		19'b0111001110110111011: color_data = Z;
		19'b0111001110110111111: color_data = Z;
		19'b0111001110111000000: color_data = Z;
		19'b0111010000010101010: color_data = Z;
		19'b0111010000010101011: color_data = Z;
		19'b0111010000010101100: color_data = Z;
		19'b0111010000010101101: color_data = Z;
		19'b0111010000010101110: color_data = Z;
		19'b0111010000010101111: color_data = Z;
		19'b0111010000010110000: color_data = Z;
		19'b0111010000010110001: color_data = Z;
		19'b0111010000010110010: color_data = Z;
		19'b0111010000010110011: color_data = Z;
		19'b0111010000010110100: color_data = Z;
		19'b0111010000010110101: color_data = Z;
		19'b0111010000010110110: color_data = Z;
		19'b0111010000010110111: color_data = Z;
		19'b0111010000010111100: color_data = Z;
		19'b0111010000010111101: color_data = Z;
		19'b0111010000010111110: color_data = Z;
		19'b0111010000010111111: color_data = Z;
		19'b0111010000011000000: color_data = Z;
		19'b0111010000011000001: color_data = Z;
		19'b0111010000011000010: color_data = Z;
		19'b0111010000011000011: color_data = Z;
		19'b0111010000100001011: color_data = Z;
		19'b0111010000100001100: color_data = Z;
		19'b0111010000100001101: color_data = Z;
		19'b0111010000100001110: color_data = Z;
		19'b0111010000100010100: color_data = Z;
		19'b0111010000100010101: color_data = Z;
		19'b0111010000100010110: color_data = Z;
		19'b0111010000100010111: color_data = Z;
		19'b0111010000100011011: color_data = Z;
		19'b0111010000100011100: color_data = Z;
		19'b0111010000100011101: color_data = Z;
		19'b0111010000100011110: color_data = Z;
		19'b0111010000100011111: color_data = Z;
		19'b0111010000100100000: color_data = Z;
		19'b0111010000100100001: color_data = Z;
		19'b0111010000100100010: color_data = Z;
		19'b0111010000100100011: color_data = Z;
		19'b0111010000100100100: color_data = Z;
		19'b0111010000100100101: color_data = Z;
		19'b0111010000100100110: color_data = Z;
		19'b0111010000100100111: color_data = Z;
		19'b0111010000100101000: color_data = Z;
		19'b0111010000100101001: color_data = Z;
		19'b0111010000100101010: color_data = Z;
		19'b0111010000100101011: color_data = Z;
		19'b0111010000100101100: color_data = Z;
		19'b0111010000100101101: color_data = Z;
		19'b0111010000100101110: color_data = Z;
		19'b0111010000100101111: color_data = Z;
		19'b0111010000100110000: color_data = Z;
		19'b0111010000100110001: color_data = Z;
		19'b0111010000100110010: color_data = Z;
		19'b0111010000100110011: color_data = Z;
		19'b0111010000100110100: color_data = Z;
		19'b0111010000100110101: color_data = Z;
		19'b0111010000100110110: color_data = Z;
		19'b0111010000100110111: color_data = Z;
		19'b0111010000100111000: color_data = Z;
		19'b0111010000100111011: color_data = Z;
		19'b0111010000100111100: color_data = Z;
		19'b0111010000100111101: color_data = Z;
		19'b0111010000100111110: color_data = Z;
		19'b0111010000100111111: color_data = Z;
		19'b0111010000101000000: color_data = Z;
		19'b0111010000101000001: color_data = Z;
		19'b0111010000101000010: color_data = Z;
		19'b0111010000101000011: color_data = Z;
		19'b0111010000101000100: color_data = Z;
		19'b0111010000101000101: color_data = Z;
		19'b0111010000101000110: color_data = Z;
		19'b0111010000101000111: color_data = Z;
		19'b0111010000101001000: color_data = Z;
		19'b0111010000101001001: color_data = Z;
		19'b0111010000101001010: color_data = Z;
		19'b0111010000101001011: color_data = Z;
		19'b0111010000101001100: color_data = Z;
		19'b0111010000101001101: color_data = Z;
		19'b0111010000101001110: color_data = Z;
		19'b0111010000101001111: color_data = Z;
		19'b0111010000101010000: color_data = Z;
		19'b0111010000101010001: color_data = Z;
		19'b0111010000101010010: color_data = Z;
		19'b0111010000101010011: color_data = Z;
		19'b0111010000101010100: color_data = Z;
		19'b0111010000101010101: color_data = Z;
		19'b0111010000101010110: color_data = Z;
		19'b0111010000101010111: color_data = Z;
		19'b0111010000101011000: color_data = Z;
		19'b0111010000101011001: color_data = Z;
		19'b0111010000101011010: color_data = Z;
		19'b0111010000101011011: color_data = Z;
		19'b0111010000101011100: color_data = Z;
		19'b0111010000101011101: color_data = Z;
		19'b0111010000101011110: color_data = Z;
		19'b0111010000101011111: color_data = Z;
		19'b0111010000101100000: color_data = Z;
		19'b0111010000101100001: color_data = Z;
		19'b0111010000101100010: color_data = Z;
		19'b0111010000101100011: color_data = Z;
		19'b0111010000101100100: color_data = Z;
		19'b0111010000101100101: color_data = Z;
		19'b0111010000101100110: color_data = Z;
		19'b0111010000101100111: color_data = Z;
		19'b0111010000101101000: color_data = Z;
		19'b0111010000101101001: color_data = Z;
		19'b0111010000101101010: color_data = Z;
		19'b0111010000101101011: color_data = Z;
		19'b0111010000101101100: color_data = Z;
		19'b0111010000101101101: color_data = Z;
		19'b0111010000101101110: color_data = Z;
		19'b0111010000101110000: color_data = Z;
		19'b0111010000101110001: color_data = Z;
		19'b0111010000101110010: color_data = Z;
		19'b0111010000101110011: color_data = Z;
		19'b0111010000101110100: color_data = Z;
		19'b0111010000101110101: color_data = Z;
		19'b0111010000101110110: color_data = Z;
		19'b0111010000101110111: color_data = Z;
		19'b0111010000101111000: color_data = Z;
		19'b0111010000101111001: color_data = Z;
		19'b0111010000101111010: color_data = Z;
		19'b0111010000101111011: color_data = Z;
		19'b0111010000101111100: color_data = Z;
		19'b0111010000101111101: color_data = Z;
		19'b0111010000101111110: color_data = Z;
		19'b0111010000101111111: color_data = Z;
		19'b0111010000110000000: color_data = Z;
		19'b0111010000110000001: color_data = Z;
		19'b0111010000110000010: color_data = Z;
		19'b0111010000110000011: color_data = Z;
		19'b0111010000110000100: color_data = Z;
		19'b0111010000110000101: color_data = Z;
		19'b0111010000110000110: color_data = Z;
		19'b0111010000110000111: color_data = Z;
		19'b0111010000110001011: color_data = Z;
		19'b0111010000110001100: color_data = Z;
		19'b0111010000110001101: color_data = Z;
		19'b0111010000110001110: color_data = Z;
		19'b0111010000110001111: color_data = Z;
		19'b0111010000110010000: color_data = Z;
		19'b0111010000110010001: color_data = Z;
		19'b0111010000110010010: color_data = Z;
		19'b0111010000110010011: color_data = Z;
		19'b0111010000110010100: color_data = Z;
		19'b0111010000110010101: color_data = Z;
		19'b0111010000110010110: color_data = Z;
		19'b0111010000110011001: color_data = Z;
		19'b0111010000110011010: color_data = Z;
		19'b0111010000110011011: color_data = Z;
		19'b0111010000110011100: color_data = Z;
		19'b0111010000110011101: color_data = Z;
		19'b0111010000110011110: color_data = Z;
		19'b0111010000110011111: color_data = Z;
		19'b0111010000110100000: color_data = Z;
		19'b0111010000110100001: color_data = Z;
		19'b0111010000110100010: color_data = Z;
		19'b0111010000110100011: color_data = Z;
		19'b0111010000110100100: color_data = Z;
		19'b0111010000110100101: color_data = Z;
		19'b0111010000110100110: color_data = Z;
		19'b0111010000110100111: color_data = Z;
		19'b0111010000110101000: color_data = Z;
		19'b0111010000110101001: color_data = Z;
		19'b0111010000110101010: color_data = Z;
		19'b0111010000110101011: color_data = Z;
		19'b0111010000110101100: color_data = Z;
		19'b0111010000110110011: color_data = Z;
		19'b0111010000110110100: color_data = Z;
		19'b0111010000110110101: color_data = Z;
		19'b0111010000110110110: color_data = Z;
		19'b0111010000110110111: color_data = Z;
		19'b0111010000110111000: color_data = Z;
		19'b0111010000110111001: color_data = Z;
		19'b0111010000110111010: color_data = Z;
		19'b0111010000110111011: color_data = Z;
		19'b0111010000110111101: color_data = Z;
		19'b0111010000110111110: color_data = Z;
		19'b0111010000110111111: color_data = Z;
		19'b0111010000111000000: color_data = Z;
		19'b0111010000111000001: color_data = Z;
		19'b0111010010010101011: color_data = Z;
		19'b0111010010010101100: color_data = Z;
		19'b0111010010010101101: color_data = Z;
		19'b0111010010010101110: color_data = Z;
		19'b0111010010010101111: color_data = Z;
		19'b0111010010010110000: color_data = Z;
		19'b0111010010010110001: color_data = Z;
		19'b0111010010010110010: color_data = Z;
		19'b0111010010010110011: color_data = Z;
		19'b0111010010010110100: color_data = Z;
		19'b0111010010010110101: color_data = Z;
		19'b0111010010010110110: color_data = Z;
		19'b0111010010010110111: color_data = Z;
		19'b0111010010010111100: color_data = Z;
		19'b0111010010010111101: color_data = Z;
		19'b0111010010010111110: color_data = Z;
		19'b0111010010010111111: color_data = Z;
		19'b0111010010011000000: color_data = Z;
		19'b0111010010011000001: color_data = Z;
		19'b0111010010011000010: color_data = Z;
		19'b0111010010011000011: color_data = Z;
		19'b0111010010011000100: color_data = Z;
		19'b0111010010011001000: color_data = Z;
		19'b0111010010011001001: color_data = Z;
		19'b0111010010011001010: color_data = Z;
		19'b0111010010100001010: color_data = Z;
		19'b0111010010100001011: color_data = Z;
		19'b0111010010100001100: color_data = Z;
		19'b0111010010100001101: color_data = Z;
		19'b0111010010100010100: color_data = Z;
		19'b0111010010100010101: color_data = Z;
		19'b0111010010100010110: color_data = Z;
		19'b0111010010100011011: color_data = Z;
		19'b0111010010100011100: color_data = Z;
		19'b0111010010100011101: color_data = Z;
		19'b0111010010100011110: color_data = Z;
		19'b0111010010100011111: color_data = Z;
		19'b0111010010100100000: color_data = Z;
		19'b0111010010100100001: color_data = Z;
		19'b0111010010100100010: color_data = Z;
		19'b0111010010100100011: color_data = Z;
		19'b0111010010100100100: color_data = Z;
		19'b0111010010100100101: color_data = Z;
		19'b0111010010100100110: color_data = Z;
		19'b0111010010100100111: color_data = Z;
		19'b0111010010100101000: color_data = Z;
		19'b0111010010100101001: color_data = Z;
		19'b0111010010100101010: color_data = Z;
		19'b0111010010100101011: color_data = Z;
		19'b0111010010100101100: color_data = Z;
		19'b0111010010100101101: color_data = Z;
		19'b0111010010100101110: color_data = Z;
		19'b0111010010100101111: color_data = Z;
		19'b0111010010100110000: color_data = Z;
		19'b0111010010100110001: color_data = Z;
		19'b0111010010100110010: color_data = Z;
		19'b0111010010100110011: color_data = Z;
		19'b0111010010100110100: color_data = Z;
		19'b0111010010100110101: color_data = Z;
		19'b0111010010100110110: color_data = Z;
		19'b0111010010100110111: color_data = Z;
		19'b0111010010100111000: color_data = Z;
		19'b0111010010100111010: color_data = Z;
		19'b0111010010100111011: color_data = Z;
		19'b0111010010100111100: color_data = Z;
		19'b0111010010100111101: color_data = Z;
		19'b0111010010100111110: color_data = Z;
		19'b0111010010100111111: color_data = Z;
		19'b0111010010101000000: color_data = Z;
		19'b0111010010101000001: color_data = Z;
		19'b0111010010101000010: color_data = Z;
		19'b0111010010101000011: color_data = Z;
		19'b0111010010101000100: color_data = Z;
		19'b0111010010101000101: color_data = Z;
		19'b0111010010101000110: color_data = Z;
		19'b0111010010101000111: color_data = Z;
		19'b0111010010101001000: color_data = Z;
		19'b0111010010101001001: color_data = Z;
		19'b0111010010101001010: color_data = Z;
		19'b0111010010101001011: color_data = Z;
		19'b0111010010101001100: color_data = Z;
		19'b0111010010101001101: color_data = Z;
		19'b0111010010101001110: color_data = Z;
		19'b0111010010101001111: color_data = Z;
		19'b0111010010101010000: color_data = Z;
		19'b0111010010101010001: color_data = Z;
		19'b0111010010101010010: color_data = Z;
		19'b0111010010101010011: color_data = Z;
		19'b0111010010101010100: color_data = Z;
		19'b0111010010101010101: color_data = Z;
		19'b0111010010101010110: color_data = Z;
		19'b0111010010101010111: color_data = Z;
		19'b0111010010101011000: color_data = Z;
		19'b0111010010101011001: color_data = Z;
		19'b0111010010101011010: color_data = Z;
		19'b0111010010101011011: color_data = Z;
		19'b0111010010101011100: color_data = Z;
		19'b0111010010101011101: color_data = Z;
		19'b0111010010101011110: color_data = Z;
		19'b0111010010101011111: color_data = Z;
		19'b0111010010101100000: color_data = Z;
		19'b0111010010101100001: color_data = Z;
		19'b0111010010101100010: color_data = Z;
		19'b0111010010101100011: color_data = Z;
		19'b0111010010101100100: color_data = Z;
		19'b0111010010101100101: color_data = Z;
		19'b0111010010101100110: color_data = Z;
		19'b0111010010101100111: color_data = Z;
		19'b0111010010101101000: color_data = Z;
		19'b0111010010101101001: color_data = Z;
		19'b0111010010101101010: color_data = Z;
		19'b0111010010101101011: color_data = Z;
		19'b0111010010101101100: color_data = Z;
		19'b0111010010101101101: color_data = Z;
		19'b0111010010101101110: color_data = Z;
		19'b0111010010101101111: color_data = Z;
		19'b0111010010101110000: color_data = Z;
		19'b0111010010101110001: color_data = Z;
		19'b0111010010101110010: color_data = Z;
		19'b0111010010101110011: color_data = Z;
		19'b0111010010101110100: color_data = Z;
		19'b0111010010101110101: color_data = Z;
		19'b0111010010101110110: color_data = Z;
		19'b0111010010101110111: color_data = Z;
		19'b0111010010101111000: color_data = Z;
		19'b0111010010101111001: color_data = Z;
		19'b0111010010101111010: color_data = Z;
		19'b0111010010101111011: color_data = Z;
		19'b0111010010101111100: color_data = Z;
		19'b0111010010101111101: color_data = Z;
		19'b0111010010101111110: color_data = Z;
		19'b0111010010101111111: color_data = Z;
		19'b0111010010110000000: color_data = Z;
		19'b0111010010110000001: color_data = Z;
		19'b0111010010110000010: color_data = Z;
		19'b0111010010110000011: color_data = Z;
		19'b0111010010110000100: color_data = Z;
		19'b0111010010110000101: color_data = Z;
		19'b0111010010110000110: color_data = Z;
		19'b0111010010110000111: color_data = Z;
		19'b0111010010110001100: color_data = Z;
		19'b0111010010110001101: color_data = Z;
		19'b0111010010110001110: color_data = Z;
		19'b0111010010110001111: color_data = Z;
		19'b0111010010110010000: color_data = Z;
		19'b0111010010110010001: color_data = Z;
		19'b0111010010110010010: color_data = Z;
		19'b0111010010110010011: color_data = Z;
		19'b0111010010110010100: color_data = Z;
		19'b0111010010110010101: color_data = Z;
		19'b0111010010110010110: color_data = Z;
		19'b0111010010110010111: color_data = Z;
		19'b0111010010110011000: color_data = Z;
		19'b0111010010110011001: color_data = Z;
		19'b0111010010110011010: color_data = Z;
		19'b0111010010110011011: color_data = Z;
		19'b0111010010110011100: color_data = Z;
		19'b0111010010110011101: color_data = Z;
		19'b0111010010110011110: color_data = Z;
		19'b0111010010110011111: color_data = Z;
		19'b0111010010110100000: color_data = Z;
		19'b0111010010110100001: color_data = Z;
		19'b0111010010110100010: color_data = Z;
		19'b0111010010110100011: color_data = Z;
		19'b0111010010110100100: color_data = Z;
		19'b0111010010110100101: color_data = Z;
		19'b0111010010110100110: color_data = Z;
		19'b0111010010110100111: color_data = Z;
		19'b0111010010110101000: color_data = Z;
		19'b0111010010110101001: color_data = Z;
		19'b0111010010110101010: color_data = Z;
		19'b0111010010110101011: color_data = Z;
		19'b0111010010110110010: color_data = Z;
		19'b0111010010110110011: color_data = Z;
		19'b0111010010110110100: color_data = Z;
		19'b0111010010110110101: color_data = Z;
		19'b0111010010110110110: color_data = Z;
		19'b0111010010110110111: color_data = Z;
		19'b0111010010110111000: color_data = Z;
		19'b0111010010110111001: color_data = Z;
		19'b0111010010110111010: color_data = Z;
		19'b0111010010110111011: color_data = Z;
		19'b0111010010110111100: color_data = Z;
		19'b0111010010110111101: color_data = Z;
		19'b0111010010110111110: color_data = Z;
		19'b0111010010110111111: color_data = Z;
		19'b0111010010111000000: color_data = Z;
		19'b0111010010111000001: color_data = Z;
		19'b0111010100010101011: color_data = Z;
		19'b0111010100010101100: color_data = Z;
		19'b0111010100010101101: color_data = Z;
		19'b0111010100010101110: color_data = Z;
		19'b0111010100010101111: color_data = Z;
		19'b0111010100010110000: color_data = Z;
		19'b0111010100010110001: color_data = Z;
		19'b0111010100010110010: color_data = Z;
		19'b0111010100010110011: color_data = Z;
		19'b0111010100010110100: color_data = Z;
		19'b0111010100010110101: color_data = Z;
		19'b0111010100010110110: color_data = Z;
		19'b0111010100010110111: color_data = Z;
		19'b0111010100010111000: color_data = Z;
		19'b0111010100010111101: color_data = Z;
		19'b0111010100010111110: color_data = Z;
		19'b0111010100010111111: color_data = Z;
		19'b0111010100011000000: color_data = Z;
		19'b0111010100011000001: color_data = Z;
		19'b0111010100011000010: color_data = Z;
		19'b0111010100011000011: color_data = Z;
		19'b0111010100011000100: color_data = Z;
		19'b0111010100011000101: color_data = Z;
		19'b0111010100011000110: color_data = Z;
		19'b0111010100011000111: color_data = Z;
		19'b0111010100011001000: color_data = Z;
		19'b0111010100011001001: color_data = Z;
		19'b0111010100011001010: color_data = Z;
		19'b0111010100011001011: color_data = Z;
		19'b0111010100011001100: color_data = Z;
		19'b0111010100100001001: color_data = Z;
		19'b0111010100100001010: color_data = Z;
		19'b0111010100100001011: color_data = Z;
		19'b0111010100100001100: color_data = Z;
		19'b0111010100100001101: color_data = Z;
		19'b0111010100100010011: color_data = Z;
		19'b0111010100100010100: color_data = Z;
		19'b0111010100100010101: color_data = Z;
		19'b0111010100100010110: color_data = Z;
		19'b0111010100100011011: color_data = Z;
		19'b0111010100100011100: color_data = Z;
		19'b0111010100100011101: color_data = Z;
		19'b0111010100100011110: color_data = Z;
		19'b0111010100100011111: color_data = Z;
		19'b0111010100100100000: color_data = Z;
		19'b0111010100100100001: color_data = Z;
		19'b0111010100100100010: color_data = Z;
		19'b0111010100100100011: color_data = Z;
		19'b0111010100100100100: color_data = Z;
		19'b0111010100100100101: color_data = Z;
		19'b0111010100100100110: color_data = Z;
		19'b0111010100100100111: color_data = Z;
		19'b0111010100100101000: color_data = Z;
		19'b0111010100100101001: color_data = Z;
		19'b0111010100100101010: color_data = Z;
		19'b0111010100100101011: color_data = Z;
		19'b0111010100100101100: color_data = Z;
		19'b0111010100100101101: color_data = Z;
		19'b0111010100100101110: color_data = Z;
		19'b0111010100100101111: color_data = Z;
		19'b0111010100100110000: color_data = Z;
		19'b0111010100100110001: color_data = Z;
		19'b0111010100100110010: color_data = Z;
		19'b0111010100100110011: color_data = Z;
		19'b0111010100100110100: color_data = Z;
		19'b0111010100100110101: color_data = Z;
		19'b0111010100100110110: color_data = Z;
		19'b0111010100100110111: color_data = Z;
		19'b0111010100100111010: color_data = Z;
		19'b0111010100100111011: color_data = Z;
		19'b0111010100100111100: color_data = Z;
		19'b0111010100100111101: color_data = Z;
		19'b0111010100100111110: color_data = Z;
		19'b0111010100100111111: color_data = Z;
		19'b0111010100101000000: color_data = Z;
		19'b0111010100101000001: color_data = Z;
		19'b0111010100101000010: color_data = Z;
		19'b0111010100101000011: color_data = Z;
		19'b0111010100101000100: color_data = Z;
		19'b0111010100101000101: color_data = Z;
		19'b0111010100101000110: color_data = Z;
		19'b0111010100101000111: color_data = Z;
		19'b0111010100101001000: color_data = Z;
		19'b0111010100101001001: color_data = Z;
		19'b0111010100101001010: color_data = Z;
		19'b0111010100101001011: color_data = Z;
		19'b0111010100101001100: color_data = Z;
		19'b0111010100101001101: color_data = Z;
		19'b0111010100101001110: color_data = Z;
		19'b0111010100101001111: color_data = Z;
		19'b0111010100101010000: color_data = Z;
		19'b0111010100101010001: color_data = Z;
		19'b0111010100101010010: color_data = Z;
		19'b0111010100101010011: color_data = Z;
		19'b0111010100101010100: color_data = Z;
		19'b0111010100101010101: color_data = Z;
		19'b0111010100101010110: color_data = Z;
		19'b0111010100101010111: color_data = Z;
		19'b0111010100101011000: color_data = Z;
		19'b0111010100101011001: color_data = Z;
		19'b0111010100101011010: color_data = Z;
		19'b0111010100101011011: color_data = Z;
		19'b0111010100101011100: color_data = Z;
		19'b0111010100101011101: color_data = Z;
		19'b0111010100101011110: color_data = Z;
		19'b0111010100101011111: color_data = Z;
		19'b0111010100101100000: color_data = Z;
		19'b0111010100101100001: color_data = Z;
		19'b0111010100101100010: color_data = Z;
		19'b0111010100101100011: color_data = Z;
		19'b0111010100101100100: color_data = Z;
		19'b0111010100101100101: color_data = Z;
		19'b0111010100101100110: color_data = Z;
		19'b0111010100101100111: color_data = Z;
		19'b0111010100101101000: color_data = Z;
		19'b0111010100101101001: color_data = Z;
		19'b0111010100101101010: color_data = Z;
		19'b0111010100101101011: color_data = Z;
		19'b0111010100101101101: color_data = Z;
		19'b0111010100101101110: color_data = Z;
		19'b0111010100101101111: color_data = Z;
		19'b0111010100101110000: color_data = Z;
		19'b0111010100101110001: color_data = Z;
		19'b0111010100101110010: color_data = Z;
		19'b0111010100101110011: color_data = Z;
		19'b0111010100101110100: color_data = Z;
		19'b0111010100101110101: color_data = Z;
		19'b0111010100101110110: color_data = Z;
		19'b0111010100101110111: color_data = Z;
		19'b0111010100101111000: color_data = Z;
		19'b0111010100101111001: color_data = Z;
		19'b0111010100101111010: color_data = Z;
		19'b0111010100101111011: color_data = Z;
		19'b0111010100101111100: color_data = Z;
		19'b0111010100101111101: color_data = Z;
		19'b0111010100101111110: color_data = Z;
		19'b0111010100101111111: color_data = Z;
		19'b0111010100110000000: color_data = Z;
		19'b0111010100110000001: color_data = Z;
		19'b0111010100110000010: color_data = Z;
		19'b0111010100110000011: color_data = Z;
		19'b0111010100110000100: color_data = Z;
		19'b0111010100110000101: color_data = Z;
		19'b0111010100110000110: color_data = Z;
		19'b0111010100110001100: color_data = Z;
		19'b0111010100110001101: color_data = Z;
		19'b0111010100110001111: color_data = Z;
		19'b0111010100110010000: color_data = Z;
		19'b0111010100110010001: color_data = Z;
		19'b0111010100110010010: color_data = Z;
		19'b0111010100110010011: color_data = Z;
		19'b0111010100110010100: color_data = Z;
		19'b0111010100110010101: color_data = Z;
		19'b0111010100110010110: color_data = Z;
		19'b0111010100110010111: color_data = Z;
		19'b0111010100110011000: color_data = Z;
		19'b0111010100110011001: color_data = Z;
		19'b0111010100110011010: color_data = Z;
		19'b0111010100110011011: color_data = Z;
		19'b0111010100110011100: color_data = Z;
		19'b0111010100110011101: color_data = Z;
		19'b0111010100110011110: color_data = Z;
		19'b0111010100110011111: color_data = Z;
		19'b0111010100110100000: color_data = Z;
		19'b0111010100110100001: color_data = Z;
		19'b0111010100110100010: color_data = Z;
		19'b0111010100110100011: color_data = Z;
		19'b0111010100110100100: color_data = Z;
		19'b0111010100110100101: color_data = Z;
		19'b0111010100110100110: color_data = Z;
		19'b0111010100110100111: color_data = Z;
		19'b0111010100110101000: color_data = Z;
		19'b0111010100110101001: color_data = Z;
		19'b0111010100110101010: color_data = Z;
		19'b0111010100110110001: color_data = Z;
		19'b0111010100110110010: color_data = Z;
		19'b0111010100110110011: color_data = Z;
		19'b0111010100110110100: color_data = Z;
		19'b0111010100110110101: color_data = Z;
		19'b0111010100110110110: color_data = Z;
		19'b0111010100110110111: color_data = Z;
		19'b0111010100110111000: color_data = Z;
		19'b0111010100110111001: color_data = Z;
		19'b0111010100110111011: color_data = Z;
		19'b0111010100110111100: color_data = Z;
		19'b0111010100110111101: color_data = Z;
		19'b0111010100110111110: color_data = Z;
		19'b0111010100110111111: color_data = Z;
		19'b0111010100111000000: color_data = Z;
		19'b0111010100111000001: color_data = Z;
		19'b0111010110010101011: color_data = Z;
		19'b0111010110010101100: color_data = Z;
		19'b0111010110010101101: color_data = Z;
		19'b0111010110010101110: color_data = Z;
		19'b0111010110010101111: color_data = Z;
		19'b0111010110010110000: color_data = Z;
		19'b0111010110010110001: color_data = Z;
		19'b0111010110010110010: color_data = Z;
		19'b0111010110010110011: color_data = Z;
		19'b0111010110010110100: color_data = Z;
		19'b0111010110010110101: color_data = Z;
		19'b0111010110010110110: color_data = Z;
		19'b0111010110010110111: color_data = Z;
		19'b0111010110010111000: color_data = Z;
		19'b0111010110010111101: color_data = Z;
		19'b0111010110010111110: color_data = Z;
		19'b0111010110010111111: color_data = Z;
		19'b0111010110011000000: color_data = Z;
		19'b0111010110011000001: color_data = Z;
		19'b0111010110011000010: color_data = Z;
		19'b0111010110011000011: color_data = Z;
		19'b0111010110011000100: color_data = Z;
		19'b0111010110011000101: color_data = Z;
		19'b0111010110011000110: color_data = Z;
		19'b0111010110011000111: color_data = Z;
		19'b0111010110011001000: color_data = Z;
		19'b0111010110011001001: color_data = Z;
		19'b0111010110011001010: color_data = Z;
		19'b0111010110011001011: color_data = Z;
		19'b0111010110011001100: color_data = Z;
		19'b0111010110011001101: color_data = Z;
		19'b0111010110011001110: color_data = Z;
		19'b0111010110011001111: color_data = Z;
		19'b0111010110011010000: color_data = Z;
		19'b0111010110011010001: color_data = Z;
		19'b0111010110011010010: color_data = Z;
		19'b0111010110011010011: color_data = Z;
		19'b0111010110100001001: color_data = Z;
		19'b0111010110100001010: color_data = Z;
		19'b0111010110100001011: color_data = Z;
		19'b0111010110100001100: color_data = Z;
		19'b0111010110100010011: color_data = Z;
		19'b0111010110100010100: color_data = Z;
		19'b0111010110100010101: color_data = Z;
		19'b0111010110100010110: color_data = Z;
		19'b0111010110100011011: color_data = Z;
		19'b0111010110100011100: color_data = Z;
		19'b0111010110100011101: color_data = Z;
		19'b0111010110100011110: color_data = Z;
		19'b0111010110100011111: color_data = Z;
		19'b0111010110100100000: color_data = Z;
		19'b0111010110100100001: color_data = Z;
		19'b0111010110100100010: color_data = Z;
		19'b0111010110100100011: color_data = Z;
		19'b0111010110100100100: color_data = Z;
		19'b0111010110100100101: color_data = Z;
		19'b0111010110100100110: color_data = Z;
		19'b0111010110100100111: color_data = Z;
		19'b0111010110100101000: color_data = Z;
		19'b0111010110100101001: color_data = Z;
		19'b0111010110100101010: color_data = Z;
		19'b0111010110100101011: color_data = Z;
		19'b0111010110100101100: color_data = Z;
		19'b0111010110100101101: color_data = Z;
		19'b0111010110100101110: color_data = Z;
		19'b0111010110100101111: color_data = Z;
		19'b0111010110100110000: color_data = Z;
		19'b0111010110100110001: color_data = Z;
		19'b0111010110100110010: color_data = Z;
		19'b0111010110100110011: color_data = Z;
		19'b0111010110100110100: color_data = Z;
		19'b0111010110100110101: color_data = Z;
		19'b0111010110100110110: color_data = Z;
		19'b0111010110100111001: color_data = Z;
		19'b0111010110100111010: color_data = Z;
		19'b0111010110100111011: color_data = Z;
		19'b0111010110100111100: color_data = Z;
		19'b0111010110100111101: color_data = Z;
		19'b0111010110100111110: color_data = Z;
		19'b0111010110100111111: color_data = Z;
		19'b0111010110101000000: color_data = Z;
		19'b0111010110101000001: color_data = Z;
		19'b0111010110101000010: color_data = Z;
		19'b0111010110101000011: color_data = Z;
		19'b0111010110101000100: color_data = Z;
		19'b0111010110101000101: color_data = Z;
		19'b0111010110101000110: color_data = Z;
		19'b0111010110101000111: color_data = Z;
		19'b0111010110101001000: color_data = Z;
		19'b0111010110101001001: color_data = Z;
		19'b0111010110101001010: color_data = Z;
		19'b0111010110101001011: color_data = Z;
		19'b0111010110101001100: color_data = Z;
		19'b0111010110101001101: color_data = Z;
		19'b0111010110101001110: color_data = Z;
		19'b0111010110101001111: color_data = Z;
		19'b0111010110101010000: color_data = Z;
		19'b0111010110101010001: color_data = Z;
		19'b0111010110101010010: color_data = Z;
		19'b0111010110101010011: color_data = Z;
		19'b0111010110101010100: color_data = Z;
		19'b0111010110101010101: color_data = Z;
		19'b0111010110101010110: color_data = Z;
		19'b0111010110101010111: color_data = Z;
		19'b0111010110101011000: color_data = Z;
		19'b0111010110101011001: color_data = Z;
		19'b0111010110101011010: color_data = Z;
		19'b0111010110101011011: color_data = Z;
		19'b0111010110101011100: color_data = Z;
		19'b0111010110101011101: color_data = Z;
		19'b0111010110101011110: color_data = Z;
		19'b0111010110101011111: color_data = Z;
		19'b0111010110101100000: color_data = Z;
		19'b0111010110101100001: color_data = Z;
		19'b0111010110101100010: color_data = Z;
		19'b0111010110101100011: color_data = Z;
		19'b0111010110101100100: color_data = Z;
		19'b0111010110101100101: color_data = Z;
		19'b0111010110101100110: color_data = Z;
		19'b0111010110101100111: color_data = Z;
		19'b0111010110101101000: color_data = Z;
		19'b0111010110101101001: color_data = Z;
		19'b0111010110101101010: color_data = Z;
		19'b0111010110101101011: color_data = Z;
		19'b0111010110101101100: color_data = Z;
		19'b0111010110101101101: color_data = Z;
		19'b0111010110101101110: color_data = Z;
		19'b0111010110101101111: color_data = Z;
		19'b0111010110101110000: color_data = Z;
		19'b0111010110101110001: color_data = Z;
		19'b0111010110101110010: color_data = Z;
		19'b0111010110101110011: color_data = Z;
		19'b0111010110101110100: color_data = Z;
		19'b0111010110101110101: color_data = Z;
		19'b0111010110101110110: color_data = Z;
		19'b0111010110101110111: color_data = Z;
		19'b0111010110101111000: color_data = Z;
		19'b0111010110101111001: color_data = Z;
		19'b0111010110101111010: color_data = Z;
		19'b0111010110101111011: color_data = Z;
		19'b0111010110101111100: color_data = Z;
		19'b0111010110101111101: color_data = Z;
		19'b0111010110101111110: color_data = Z;
		19'b0111010110101111111: color_data = Z;
		19'b0111010110110000000: color_data = Z;
		19'b0111010110110000001: color_data = Z;
		19'b0111010110110000010: color_data = Z;
		19'b0111010110110000011: color_data = Z;
		19'b0111010110110000100: color_data = Z;
		19'b0111010110110000101: color_data = Z;
		19'b0111010110110000110: color_data = Z;
		19'b0111010110110000111: color_data = Z;
		19'b0111010110110001000: color_data = Z;
		19'b0111010110110001101: color_data = Z;
		19'b0111010110110001111: color_data = Z;
		19'b0111010110110010000: color_data = Z;
		19'b0111010110110010001: color_data = Z;
		19'b0111010110110010010: color_data = Z;
		19'b0111010110110010011: color_data = Z;
		19'b0111010110110010100: color_data = Z;
		19'b0111010110110010101: color_data = Z;
		19'b0111010110110010110: color_data = Z;
		19'b0111010110110010111: color_data = Z;
		19'b0111010110110011000: color_data = Z;
		19'b0111010110110011001: color_data = Z;
		19'b0111010110110011010: color_data = Z;
		19'b0111010110110011011: color_data = Z;
		19'b0111010110110011100: color_data = Z;
		19'b0111010110110011101: color_data = Z;
		19'b0111010110110011110: color_data = Z;
		19'b0111010110110011111: color_data = Z;
		19'b0111010110110100000: color_data = Z;
		19'b0111010110110100001: color_data = Z;
		19'b0111010110110100010: color_data = Z;
		19'b0111010110110100011: color_data = Z;
		19'b0111010110110100100: color_data = Z;
		19'b0111010110110100101: color_data = Z;
		19'b0111010110110100110: color_data = Z;
		19'b0111010110110100111: color_data = Z;
		19'b0111010110110101000: color_data = Z;
		19'b0111010110110101001: color_data = Z;
		19'b0111010110110101010: color_data = Z;
		19'b0111010110110101011: color_data = Z;
		19'b0111010110110101100: color_data = Z;
		19'b0111010110110101101: color_data = Z;
		19'b0111010110110101110: color_data = Z;
		19'b0111010110110101111: color_data = Z;
		19'b0111010110110110000: color_data = Z;
		19'b0111010110110110001: color_data = Z;
		19'b0111010110110110010: color_data = Z;
		19'b0111010110110110011: color_data = Z;
		19'b0111010110110110100: color_data = Z;
		19'b0111010110110110101: color_data = Z;
		19'b0111010110110110110: color_data = Z;
		19'b0111010110110110111: color_data = Z;
		19'b0111010110110111000: color_data = Z;
		19'b0111010110110111001: color_data = Z;
		19'b0111010110110111010: color_data = Z;
		19'b0111010110110111011: color_data = Z;
		19'b0111010110110111100: color_data = Z;
		19'b0111010110110111101: color_data = Z;
		19'b0111010110110111110: color_data = Z;
		19'b0111010110110111111: color_data = Z;
		19'b0111010110111000000: color_data = Z;
		19'b0111010110111000001: color_data = Z;
		19'b0111011000010101100: color_data = Z;
		19'b0111011000010101101: color_data = Z;
		19'b0111011000010101110: color_data = Z;
		19'b0111011000010101111: color_data = Z;
		19'b0111011000010110000: color_data = Z;
		19'b0111011000010110001: color_data = Z;
		19'b0111011000010110010: color_data = Z;
		19'b0111011000010110011: color_data = Z;
		19'b0111011000010110100: color_data = Z;
		19'b0111011000010110101: color_data = Z;
		19'b0111011000010110110: color_data = Z;
		19'b0111011000010110111: color_data = Z;
		19'b0111011000010111000: color_data = Z;
		19'b0111011000010111001: color_data = Z;
		19'b0111011000010111111: color_data = Z;
		19'b0111011000011000000: color_data = Z;
		19'b0111011000011000001: color_data = Z;
		19'b0111011000011000010: color_data = Z;
		19'b0111011000011000011: color_data = Z;
		19'b0111011000011000100: color_data = Z;
		19'b0111011000011000101: color_data = Z;
		19'b0111011000011000110: color_data = Z;
		19'b0111011000011000111: color_data = Z;
		19'b0111011000011001000: color_data = Z;
		19'b0111011000011001001: color_data = Z;
		19'b0111011000011001010: color_data = Z;
		19'b0111011000011001011: color_data = Z;
		19'b0111011000011001100: color_data = Z;
		19'b0111011000011001101: color_data = Z;
		19'b0111011000011001110: color_data = Z;
		19'b0111011000011001111: color_data = Z;
		19'b0111011000011010000: color_data = Z;
		19'b0111011000011010001: color_data = Z;
		19'b0111011000011010010: color_data = Z;
		19'b0111011000011010011: color_data = Z;
		19'b0111011000011010100: color_data = Z;
		19'b0111011000011010101: color_data = Z;
		19'b0111011000100001000: color_data = Z;
		19'b0111011000100001001: color_data = Z;
		19'b0111011000100001010: color_data = Z;
		19'b0111011000100001011: color_data = Z;
		19'b0111011000100001100: color_data = Z;
		19'b0111011000100010010: color_data = Z;
		19'b0111011000100010011: color_data = Z;
		19'b0111011000100010100: color_data = Z;
		19'b0111011000100010101: color_data = Z;
		19'b0111011000100011010: color_data = Z;
		19'b0111011000100011011: color_data = Z;
		19'b0111011000100011100: color_data = Z;
		19'b0111011000100011101: color_data = Z;
		19'b0111011000100011110: color_data = Z;
		19'b0111011000100011111: color_data = Z;
		19'b0111011000100100000: color_data = Z;
		19'b0111011000100100001: color_data = Z;
		19'b0111011000100100010: color_data = Z;
		19'b0111011000100100011: color_data = Z;
		19'b0111011000100100100: color_data = Z;
		19'b0111011000100100101: color_data = Z;
		19'b0111011000100100110: color_data = Z;
		19'b0111011000100100111: color_data = Z;
		19'b0111011000100101000: color_data = Z;
		19'b0111011000100101001: color_data = Z;
		19'b0111011000100101010: color_data = Z;
		19'b0111011000100101011: color_data = Z;
		19'b0111011000100101100: color_data = Z;
		19'b0111011000100101101: color_data = Z;
		19'b0111011000100101110: color_data = Z;
		19'b0111011000100101111: color_data = Z;
		19'b0111011000100110000: color_data = Z;
		19'b0111011000100110001: color_data = Z;
		19'b0111011000100110010: color_data = Z;
		19'b0111011000100110011: color_data = Z;
		19'b0111011000100110100: color_data = Z;
		19'b0111011000100110101: color_data = Z;
		19'b0111011000100110110: color_data = Z;
		19'b0111011000100111000: color_data = Z;
		19'b0111011000100111001: color_data = Z;
		19'b0111011000100111010: color_data = Z;
		19'b0111011000100111011: color_data = Z;
		19'b0111011000100111100: color_data = Z;
		19'b0111011000100111101: color_data = Z;
		19'b0111011000100111110: color_data = Z;
		19'b0111011000100111111: color_data = Z;
		19'b0111011000101000000: color_data = Z;
		19'b0111011000101000001: color_data = Z;
		19'b0111011000101000010: color_data = Z;
		19'b0111011000101000011: color_data = Z;
		19'b0111011000101000100: color_data = Z;
		19'b0111011000101000101: color_data = Z;
		19'b0111011000101000110: color_data = Z;
		19'b0111011000101000111: color_data = Z;
		19'b0111011000101001000: color_data = Z;
		19'b0111011000101001001: color_data = Z;
		19'b0111011000101001010: color_data = Z;
		19'b0111011000101001011: color_data = Z;
		19'b0111011000101001100: color_data = Z;
		19'b0111011000101001101: color_data = Z;
		19'b0111011000101001110: color_data = Z;
		19'b0111011000101001111: color_data = Z;
		19'b0111011000101010000: color_data = Z;
		19'b0111011000101010001: color_data = Z;
		19'b0111011000101010010: color_data = Z;
		19'b0111011000101010011: color_data = Z;
		19'b0111011000101010100: color_data = Z;
		19'b0111011000101010101: color_data = Z;
		19'b0111011000101010110: color_data = Z;
		19'b0111011000101010111: color_data = Z;
		19'b0111011000101011000: color_data = Z;
		19'b0111011000101011001: color_data = Z;
		19'b0111011000101011010: color_data = Z;
		19'b0111011000101011011: color_data = Z;
		19'b0111011000101011100: color_data = Z;
		19'b0111011000101011101: color_data = Z;
		19'b0111011000101011110: color_data = Z;
		19'b0111011000101011111: color_data = Z;
		19'b0111011000101100000: color_data = Z;
		19'b0111011000101100001: color_data = Z;
		19'b0111011000101100010: color_data = Z;
		19'b0111011000101100011: color_data = Z;
		19'b0111011000101100100: color_data = Z;
		19'b0111011000101100101: color_data = Z;
		19'b0111011000101100110: color_data = Z;
		19'b0111011000101100111: color_data = Z;
		19'b0111011000101101000: color_data = Z;
		19'b0111011000101101001: color_data = Z;
		19'b0111011000101101010: color_data = Z;
		19'b0111011000101101011: color_data = Z;
		19'b0111011000101101100: color_data = Z;
		19'b0111011000101101101: color_data = Z;
		19'b0111011000101101110: color_data = Z;
		19'b0111011000101101111: color_data = Z;
		19'b0111011000101110000: color_data = Z;
		19'b0111011000101110001: color_data = Z;
		19'b0111011000101110010: color_data = Z;
		19'b0111011000101110011: color_data = Z;
		19'b0111011000101110100: color_data = Z;
		19'b0111011000101110101: color_data = Z;
		19'b0111011000101110110: color_data = Z;
		19'b0111011000101110111: color_data = Z;
		19'b0111011000101111000: color_data = Z;
		19'b0111011000101111001: color_data = Z;
		19'b0111011000101111010: color_data = Z;
		19'b0111011000101111011: color_data = Z;
		19'b0111011000101111100: color_data = Z;
		19'b0111011000101111101: color_data = Z;
		19'b0111011000101111110: color_data = Z;
		19'b0111011000101111111: color_data = Z;
		19'b0111011000110000000: color_data = Z;
		19'b0111011000110000001: color_data = Z;
		19'b0111011000110000010: color_data = Z;
		19'b0111011000110000011: color_data = Z;
		19'b0111011000110000100: color_data = Z;
		19'b0111011000110000101: color_data = Z;
		19'b0111011000110000110: color_data = Z;
		19'b0111011000110000111: color_data = Z;
		19'b0111011000110001000: color_data = Z;
		19'b0111011000110001001: color_data = Z;
		19'b0111011000110010000: color_data = Z;
		19'b0111011000110010001: color_data = Z;
		19'b0111011000110010010: color_data = Z;
		19'b0111011000110010011: color_data = Z;
		19'b0111011000110010100: color_data = Z;
		19'b0111011000110010101: color_data = Z;
		19'b0111011000110010110: color_data = Z;
		19'b0111011000110010111: color_data = Z;
		19'b0111011000110011000: color_data = Z;
		19'b0111011000110011001: color_data = Z;
		19'b0111011000110011010: color_data = Z;
		19'b0111011000110011011: color_data = Z;
		19'b0111011000110011100: color_data = Z;
		19'b0111011000110011101: color_data = Z;
		19'b0111011000110011110: color_data = Z;
		19'b0111011000110011111: color_data = Z;
		19'b0111011000110100000: color_data = Z;
		19'b0111011000110100001: color_data = Z;
		19'b0111011000110100010: color_data = Z;
		19'b0111011000110100011: color_data = Z;
		19'b0111011000110100100: color_data = Z;
		19'b0111011000110100101: color_data = Z;
		19'b0111011000110100110: color_data = Z;
		19'b0111011000110100111: color_data = Z;
		19'b0111011000110101000: color_data = Z;
		19'b0111011000110101001: color_data = Z;
		19'b0111011000110101010: color_data = Z;
		19'b0111011000110101011: color_data = Z;
		19'b0111011000110101100: color_data = Z;
		19'b0111011000110101101: color_data = Z;
		19'b0111011000110101110: color_data = Z;
		19'b0111011000110101111: color_data = Z;
		19'b0111011000110110000: color_data = Z;
		19'b0111011000110110001: color_data = Z;
		19'b0111011000110110010: color_data = Z;
		19'b0111011000110110011: color_data = Z;
		19'b0111011000110110100: color_data = Z;
		19'b0111011000110110101: color_data = Z;
		19'b0111011000110110110: color_data = Z;
		19'b0111011000110110111: color_data = Z;
		19'b0111011000110111000: color_data = Z;
		19'b0111011000110111001: color_data = Z;
		19'b0111011000110111010: color_data = Z;
		19'b0111011000110111011: color_data = Z;
		19'b0111011000110111100: color_data = Z;
		19'b0111011000110111101: color_data = Z;
		19'b0111011000110111110: color_data = Z;
		19'b0111011000110111111: color_data = Z;
		19'b0111011000111000000: color_data = Z;
		19'b0111011000111000001: color_data = Z;
		19'b0111011000111000010: color_data = Z;
		19'b0111011010010101100: color_data = Z;
		19'b0111011010010101101: color_data = Z;
		19'b0111011010010101110: color_data = Z;
		19'b0111011010010101111: color_data = Z;
		19'b0111011010010110000: color_data = Z;
		19'b0111011010010110001: color_data = Z;
		19'b0111011010010110010: color_data = Z;
		19'b0111011010010110011: color_data = Z;
		19'b0111011010010110100: color_data = Z;
		19'b0111011010010110101: color_data = Z;
		19'b0111011010010110110: color_data = Z;
		19'b0111011010010110111: color_data = Z;
		19'b0111011010010111000: color_data = Z;
		19'b0111011010010111001: color_data = Z;
		19'b0111011010010111010: color_data = Z;
		19'b0111011010010111111: color_data = Z;
		19'b0111011010011000000: color_data = Z;
		19'b0111011010011000001: color_data = Z;
		19'b0111011010011000010: color_data = Z;
		19'b0111011010011000011: color_data = Z;
		19'b0111011010011000100: color_data = Z;
		19'b0111011010011000101: color_data = Z;
		19'b0111011010011000110: color_data = Z;
		19'b0111011010011000111: color_data = Z;
		19'b0111011010011001000: color_data = Z;
		19'b0111011010011001001: color_data = Z;
		19'b0111011010011001010: color_data = Z;
		19'b0111011010011001011: color_data = Z;
		19'b0111011010011001100: color_data = Z;
		19'b0111011010011001101: color_data = Z;
		19'b0111011010011001110: color_data = Z;
		19'b0111011010011001111: color_data = Z;
		19'b0111011010011010000: color_data = Z;
		19'b0111011010011010001: color_data = Z;
		19'b0111011010011010010: color_data = Z;
		19'b0111011010011010011: color_data = Z;
		19'b0111011010011010100: color_data = Z;
		19'b0111011010011010101: color_data = Z;
		19'b0111011010011010110: color_data = Z;
		19'b0111011010011010111: color_data = Z;
		19'b0111011010100001000: color_data = Z;
		19'b0111011010100001001: color_data = Z;
		19'b0111011010100001010: color_data = Z;
		19'b0111011010100001011: color_data = Z;
		19'b0111011010100001100: color_data = Z;
		19'b0111011010100010001: color_data = Z;
		19'b0111011010100010010: color_data = Z;
		19'b0111011010100010011: color_data = Z;
		19'b0111011010100010100: color_data = Z;
		19'b0111011010100010101: color_data = Z;
		19'b0111011010100011001: color_data = Z;
		19'b0111011010100011010: color_data = Z;
		19'b0111011010100011011: color_data = Z;
		19'b0111011010100011100: color_data = Z;
		19'b0111011010100011101: color_data = Z;
		19'b0111011010100011110: color_data = Z;
		19'b0111011010100011111: color_data = Z;
		19'b0111011010100100000: color_data = Z;
		19'b0111011010100100001: color_data = Z;
		19'b0111011010100100010: color_data = Z;
		19'b0111011010100100011: color_data = Z;
		19'b0111011010100100100: color_data = Z;
		19'b0111011010100100101: color_data = Z;
		19'b0111011010100100110: color_data = Z;
		19'b0111011010100100111: color_data = Z;
		19'b0111011010100101000: color_data = Z;
		19'b0111011010100101001: color_data = Z;
		19'b0111011010100101010: color_data = Z;
		19'b0111011010100101011: color_data = Z;
		19'b0111011010100101100: color_data = Z;
		19'b0111011010100101101: color_data = Z;
		19'b0111011010100101110: color_data = Z;
		19'b0111011010100101111: color_data = Z;
		19'b0111011010100110000: color_data = Z;
		19'b0111011010100110001: color_data = Z;
		19'b0111011010100110010: color_data = Z;
		19'b0111011010100110011: color_data = Z;
		19'b0111011010100110100: color_data = Z;
		19'b0111011010100110101: color_data = Z;
		19'b0111011010100110110: color_data = Z;
		19'b0111011010100111000: color_data = Z;
		19'b0111011010100111001: color_data = Z;
		19'b0111011010100111010: color_data = Z;
		19'b0111011010100111011: color_data = Z;
		19'b0111011010100111100: color_data = Z;
		19'b0111011010100111101: color_data = Z;
		19'b0111011010100111110: color_data = Z;
		19'b0111011010100111111: color_data = Z;
		19'b0111011010101000000: color_data = Z;
		19'b0111011010101000001: color_data = Z;
		19'b0111011010101000010: color_data = Z;
		19'b0111011010101000011: color_data = Z;
		19'b0111011010101000100: color_data = Z;
		19'b0111011010101000101: color_data = Z;
		19'b0111011010101000110: color_data = Z;
		19'b0111011010101000111: color_data = Z;
		19'b0111011010101001000: color_data = Z;
		19'b0111011010101001001: color_data = Z;
		19'b0111011010101001010: color_data = Z;
		19'b0111011010101001011: color_data = Z;
		19'b0111011010101001100: color_data = Z;
		19'b0111011010101001101: color_data = Z;
		19'b0111011010101001110: color_data = Z;
		19'b0111011010101001111: color_data = Z;
		19'b0111011010101010000: color_data = Z;
		19'b0111011010101010001: color_data = Z;
		19'b0111011010101010010: color_data = Z;
		19'b0111011010101010011: color_data = Z;
		19'b0111011010101010100: color_data = Z;
		19'b0111011010101010101: color_data = Z;
		19'b0111011010101010110: color_data = Z;
		19'b0111011010101010111: color_data = Z;
		19'b0111011010101011000: color_data = Z;
		19'b0111011010101011001: color_data = Z;
		19'b0111011010101011010: color_data = Z;
		19'b0111011010101011011: color_data = Z;
		19'b0111011010101011100: color_data = Z;
		19'b0111011010101011101: color_data = Z;
		19'b0111011010101011110: color_data = Z;
		19'b0111011010101011111: color_data = Z;
		19'b0111011010101100000: color_data = Z;
		19'b0111011010101100001: color_data = Z;
		19'b0111011010101100010: color_data = Z;
		19'b0111011010101100011: color_data = Z;
		19'b0111011010101100100: color_data = Z;
		19'b0111011010101100101: color_data = Z;
		19'b0111011010101100110: color_data = Z;
		19'b0111011010101100111: color_data = Z;
		19'b0111011010101101000: color_data = Z;
		19'b0111011010101101001: color_data = Z;
		19'b0111011010101101010: color_data = Z;
		19'b0111011010101101011: color_data = Z;
		19'b0111011010101101100: color_data = Z;
		19'b0111011010101101101: color_data = Z;
		19'b0111011010101101110: color_data = Z;
		19'b0111011010101101111: color_data = Z;
		19'b0111011010101110000: color_data = Z;
		19'b0111011010101110001: color_data = Z;
		19'b0111011010101110010: color_data = Z;
		19'b0111011010101110011: color_data = Z;
		19'b0111011010101110100: color_data = Z;
		19'b0111011010101110101: color_data = Z;
		19'b0111011010101110110: color_data = Z;
		19'b0111011010101110111: color_data = Z;
		19'b0111011010101111000: color_data = Z;
		19'b0111011010101111001: color_data = Z;
		19'b0111011010101111010: color_data = Z;
		19'b0111011010101111011: color_data = Z;
		19'b0111011010101111100: color_data = Z;
		19'b0111011010101111101: color_data = Z;
		19'b0111011010101111110: color_data = Z;
		19'b0111011010101111111: color_data = Z;
		19'b0111011010110000000: color_data = Z;
		19'b0111011010110000001: color_data = Z;
		19'b0111011010110000010: color_data = Z;
		19'b0111011010110000011: color_data = Z;
		19'b0111011010110000100: color_data = Z;
		19'b0111011010110000101: color_data = Z;
		19'b0111011010110000110: color_data = Z;
		19'b0111011010110000111: color_data = Z;
		19'b0111011010110001000: color_data = Z;
		19'b0111011010110001001: color_data = Z;
		19'b0111011010110001010: color_data = Z;
		19'b0111011010110001011: color_data = Z;
		19'b0111011010110001100: color_data = Z;
		19'b0111011010110010001: color_data = Z;
		19'b0111011010110010010: color_data = Z;
		19'b0111011010110010011: color_data = Z;
		19'b0111011010110010100: color_data = Z;
		19'b0111011010110010101: color_data = Z;
		19'b0111011010110010110: color_data = Z;
		19'b0111011010110010111: color_data = Z;
		19'b0111011010110011000: color_data = Z;
		19'b0111011010110011001: color_data = Z;
		19'b0111011010110011010: color_data = Z;
		19'b0111011010110011011: color_data = Z;
		19'b0111011010110011100: color_data = Z;
		19'b0111011010110011101: color_data = Z;
		19'b0111011010110011110: color_data = Z;
		19'b0111011010110011111: color_data = Z;
		19'b0111011010110100000: color_data = Z;
		19'b0111011010110100001: color_data = Z;
		19'b0111011010110100010: color_data = Z;
		19'b0111011010110100011: color_data = Z;
		19'b0111011010110100100: color_data = Z;
		19'b0111011010110100101: color_data = Z;
		19'b0111011010110100110: color_data = Z;
		19'b0111011010110100111: color_data = Z;
		19'b0111011010110101000: color_data = Z;
		19'b0111011010110101001: color_data = Z;
		19'b0111011010110101010: color_data = Z;
		19'b0111011010110101011: color_data = Z;
		19'b0111011010110101100: color_data = Z;
		19'b0111011010110101101: color_data = Z;
		19'b0111011010110101110: color_data = Z;
		19'b0111011010110101111: color_data = Z;
		19'b0111011010110110000: color_data = Z;
		19'b0111011010110110001: color_data = Z;
		19'b0111011010110110010: color_data = Z;
		19'b0111011010110110011: color_data = Z;
		19'b0111011010110110100: color_data = Z;
		19'b0111011010110110101: color_data = Z;
		19'b0111011010110110110: color_data = Z;
		19'b0111011010110110111: color_data = Z;
		19'b0111011010110111000: color_data = Z;
		19'b0111011010110111001: color_data = Z;
		19'b0111011010110111010: color_data = Z;
		19'b0111011010110111011: color_data = Z;
		19'b0111011010110111100: color_data = Z;
		19'b0111011010110111101: color_data = Z;
		19'b0111011010110111110: color_data = Z;
		19'b0111011010110111111: color_data = Z;
		19'b0111011010111000000: color_data = Z;
		19'b0111011010111000001: color_data = Z;
		19'b0111011010111000010: color_data = Z;
		19'b0111011100010101100: color_data = Z;
		19'b0111011100010101101: color_data = Z;
		19'b0111011100010101110: color_data = Z;
		19'b0111011100010101111: color_data = Z;
		19'b0111011100010110000: color_data = Z;
		19'b0111011100010110001: color_data = Z;
		19'b0111011100010110010: color_data = Z;
		19'b0111011100010110011: color_data = Z;
		19'b0111011100010110100: color_data = Z;
		19'b0111011100010110101: color_data = Z;
		19'b0111011100010110110: color_data = Z;
		19'b0111011100010110111: color_data = Z;
		19'b0111011100010111000: color_data = Z;
		19'b0111011100010111001: color_data = Z;
		19'b0111011100010111010: color_data = Z;
		19'b0111011100011000010: color_data = Z;
		19'b0111011100011000011: color_data = Z;
		19'b0111011100011000100: color_data = Z;
		19'b0111011100011000101: color_data = Z;
		19'b0111011100011000110: color_data = Z;
		19'b0111011100011000111: color_data = Z;
		19'b0111011100011001000: color_data = Z;
		19'b0111011100011001001: color_data = Z;
		19'b0111011100011001010: color_data = Z;
		19'b0111011100011001011: color_data = Z;
		19'b0111011100011001100: color_data = Z;
		19'b0111011100011001101: color_data = Z;
		19'b0111011100011001110: color_data = Z;
		19'b0111011100011001111: color_data = Z;
		19'b0111011100011010000: color_data = Z;
		19'b0111011100011010001: color_data = Z;
		19'b0111011100011010010: color_data = Z;
		19'b0111011100011010011: color_data = Z;
		19'b0111011100011010100: color_data = Z;
		19'b0111011100011010101: color_data = Z;
		19'b0111011100011010110: color_data = Z;
		19'b0111011100011010111: color_data = Z;
		19'b0111011100011011000: color_data = Z;
		19'b0111011100100001000: color_data = Z;
		19'b0111011100100001001: color_data = Z;
		19'b0111011100100001010: color_data = Z;
		19'b0111011100100001011: color_data = Z;
		19'b0111011100100010001: color_data = Z;
		19'b0111011100100010010: color_data = Z;
		19'b0111011100100010011: color_data = Z;
		19'b0111011100100010100: color_data = Z;
		19'b0111011100100011001: color_data = Z;
		19'b0111011100100011010: color_data = Z;
		19'b0111011100100011011: color_data = Z;
		19'b0111011100100011100: color_data = Z;
		19'b0111011100100011101: color_data = Z;
		19'b0111011100100011110: color_data = Z;
		19'b0111011100100011111: color_data = Z;
		19'b0111011100100100000: color_data = Z;
		19'b0111011100100100001: color_data = Z;
		19'b0111011100100100010: color_data = Z;
		19'b0111011100100100011: color_data = Z;
		19'b0111011100100100100: color_data = Z;
		19'b0111011100100100101: color_data = Z;
		19'b0111011100100100110: color_data = Z;
		19'b0111011100100101000: color_data = Z;
		19'b0111011100100101001: color_data = Z;
		19'b0111011100100101010: color_data = Z;
		19'b0111011100100101011: color_data = Z;
		19'b0111011100100101100: color_data = Z;
		19'b0111011100100101101: color_data = Z;
		19'b0111011100100101110: color_data = Z;
		19'b0111011100100101111: color_data = Z;
		19'b0111011100100110000: color_data = Z;
		19'b0111011100100110001: color_data = Z;
		19'b0111011100100110010: color_data = Z;
		19'b0111011100100110011: color_data = Z;
		19'b0111011100100110100: color_data = Z;
		19'b0111011100100110101: color_data = Z;
		19'b0111011100100110110: color_data = Z;
		19'b0111011100100110111: color_data = Z;
		19'b0111011100100111000: color_data = Z;
		19'b0111011100100111001: color_data = Z;
		19'b0111011100100111010: color_data = Z;
		19'b0111011100100111011: color_data = Z;
		19'b0111011100100111100: color_data = Z;
		19'b0111011100100111101: color_data = Z;
		19'b0111011100100111110: color_data = Z;
		19'b0111011100100111111: color_data = Z;
		19'b0111011100101000000: color_data = Z;
		19'b0111011100101000001: color_data = Z;
		19'b0111011100101000010: color_data = Z;
		19'b0111011100101000011: color_data = Z;
		19'b0111011100101000100: color_data = Z;
		19'b0111011100101000101: color_data = Z;
		19'b0111011100101000110: color_data = Z;
		19'b0111011100101000111: color_data = Z;
		19'b0111011100101001000: color_data = Z;
		19'b0111011100101001001: color_data = Z;
		19'b0111011100101001010: color_data = Z;
		19'b0111011100101001011: color_data = Z;
		19'b0111011100101001100: color_data = Z;
		19'b0111011100101001101: color_data = Z;
		19'b0111011100101001110: color_data = Z;
		19'b0111011100101001111: color_data = Z;
		19'b0111011100101010000: color_data = Z;
		19'b0111011100101010001: color_data = Z;
		19'b0111011100101010010: color_data = Z;
		19'b0111011100101010011: color_data = Z;
		19'b0111011100101010100: color_data = Z;
		19'b0111011100101010101: color_data = Z;
		19'b0111011100101010110: color_data = Z;
		19'b0111011100101010111: color_data = Z;
		19'b0111011100101011000: color_data = Z;
		19'b0111011100101011001: color_data = Z;
		19'b0111011100101011010: color_data = Z;
		19'b0111011100101011011: color_data = Z;
		19'b0111011100101011100: color_data = Z;
		19'b0111011100101011101: color_data = Z;
		19'b0111011100101011110: color_data = Z;
		19'b0111011100101011111: color_data = Z;
		19'b0111011100101100000: color_data = Z;
		19'b0111011100101100001: color_data = Z;
		19'b0111011100101100010: color_data = Z;
		19'b0111011100101100011: color_data = Z;
		19'b0111011100101100100: color_data = Z;
		19'b0111011100101100101: color_data = Z;
		19'b0111011100101100110: color_data = Z;
		19'b0111011100101100111: color_data = Z;
		19'b0111011100101101000: color_data = Z;
		19'b0111011100101101001: color_data = Z;
		19'b0111011100101101010: color_data = Z;
		19'b0111011100101101011: color_data = Z;
		19'b0111011100101101100: color_data = Z;
		19'b0111011100101101101: color_data = Z;
		19'b0111011100101101110: color_data = Z;
		19'b0111011100101101111: color_data = Z;
		19'b0111011100101110000: color_data = Z;
		19'b0111011100101110001: color_data = Z;
		19'b0111011100101110010: color_data = Z;
		19'b0111011100101110011: color_data = Z;
		19'b0111011100101110100: color_data = Z;
		19'b0111011100101110101: color_data = Z;
		19'b0111011100101110110: color_data = Z;
		19'b0111011100101110111: color_data = Z;
		19'b0111011100101111000: color_data = Z;
		19'b0111011100101111001: color_data = Z;
		19'b0111011100101111010: color_data = Z;
		19'b0111011100101111011: color_data = Z;
		19'b0111011100101111100: color_data = Z;
		19'b0111011100101111101: color_data = Z;
		19'b0111011100101111110: color_data = Z;
		19'b0111011100101111111: color_data = Z;
		19'b0111011100110000000: color_data = Z;
		19'b0111011100110000001: color_data = Z;
		19'b0111011100110000010: color_data = Z;
		19'b0111011100110000011: color_data = Z;
		19'b0111011100110000100: color_data = Z;
		19'b0111011100110000101: color_data = Z;
		19'b0111011100110000110: color_data = Z;
		19'b0111011100110000111: color_data = Z;
		19'b0111011100110001000: color_data = Z;
		19'b0111011100110001001: color_data = Z;
		19'b0111011100110001010: color_data = Z;
		19'b0111011100110001011: color_data = Z;
		19'b0111011100110001100: color_data = Z;
		19'b0111011100110010100: color_data = Z;
		19'b0111011100110010101: color_data = Z;
		19'b0111011100110010110: color_data = Z;
		19'b0111011100110010111: color_data = Z;
		19'b0111011100110011000: color_data = Z;
		19'b0111011100110011001: color_data = Z;
		19'b0111011100110011010: color_data = Z;
		19'b0111011100110011011: color_data = Z;
		19'b0111011100110011100: color_data = Z;
		19'b0111011100110011101: color_data = Z;
		19'b0111011100110011110: color_data = Z;
		19'b0111011100110011111: color_data = Z;
		19'b0111011100110100000: color_data = Z;
		19'b0111011100110100001: color_data = Z;
		19'b0111011100110100010: color_data = Z;
		19'b0111011100110100011: color_data = Z;
		19'b0111011100110100100: color_data = Z;
		19'b0111011100110100101: color_data = Z;
		19'b0111011100110100110: color_data = Z;
		19'b0111011100110100111: color_data = Z;
		19'b0111011100110101000: color_data = Z;
		19'b0111011100110101001: color_data = Z;
		19'b0111011100110101010: color_data = Z;
		19'b0111011100110101011: color_data = Z;
		19'b0111011100110101100: color_data = Z;
		19'b0111011100110101101: color_data = Z;
		19'b0111011100110101110: color_data = Z;
		19'b0111011100110101111: color_data = Z;
		19'b0111011100110110000: color_data = Z;
		19'b0111011100110110001: color_data = Z;
		19'b0111011100110110010: color_data = Z;
		19'b0111011100110110011: color_data = Z;
		19'b0111011100110110100: color_data = Z;
		19'b0111011100110110101: color_data = Z;
		19'b0111011100110110110: color_data = Z;
		19'b0111011100110110111: color_data = Z;
		19'b0111011100110111000: color_data = Z;
		19'b0111011100110111001: color_data = Z;
		19'b0111011100110111010: color_data = Z;
		19'b0111011100110111011: color_data = Z;
		19'b0111011100110111100: color_data = Z;
		19'b0111011100110111101: color_data = Z;
		19'b0111011100110111110: color_data = Z;
		19'b0111011100110111111: color_data = Z;
		19'b0111011100111000000: color_data = Z;
		19'b0111011100111000001: color_data = Z;
		19'b0111011100111000010: color_data = Z;
		19'b0111011100111000011: color_data = Z;
		19'b0111011100111000100: color_data = Z;
		19'b0111011100111000101: color_data = Z;
		19'b0111011110010101101: color_data = Z;
		19'b0111011110010101110: color_data = Z;
		19'b0111011110010101111: color_data = Z;
		19'b0111011110010110000: color_data = Z;
		19'b0111011110010110001: color_data = Z;
		19'b0111011110010110010: color_data = Z;
		19'b0111011110010110011: color_data = Z;
		19'b0111011110010110100: color_data = Z;
		19'b0111011110010110101: color_data = Z;
		19'b0111011110010110110: color_data = Z;
		19'b0111011110010110111: color_data = Z;
		19'b0111011110010111000: color_data = Z;
		19'b0111011110010111001: color_data = Z;
		19'b0111011110010111010: color_data = Z;
		19'b0111011110010111011: color_data = Z;
		19'b0111011110011000011: color_data = Z;
		19'b0111011110011000100: color_data = Z;
		19'b0111011110011000101: color_data = Z;
		19'b0111011110011000110: color_data = Z;
		19'b0111011110011000111: color_data = Z;
		19'b0111011110011001000: color_data = Z;
		19'b0111011110011001001: color_data = Z;
		19'b0111011110011001010: color_data = Z;
		19'b0111011110011001011: color_data = Z;
		19'b0111011110011001100: color_data = Z;
		19'b0111011110011001101: color_data = Z;
		19'b0111011110011001110: color_data = Z;
		19'b0111011110011001111: color_data = Z;
		19'b0111011110011010000: color_data = Z;
		19'b0111011110011010001: color_data = Z;
		19'b0111011110011010010: color_data = Z;
		19'b0111011110011010011: color_data = Z;
		19'b0111011110011010100: color_data = Z;
		19'b0111011110011010101: color_data = Z;
		19'b0111011110011010110: color_data = Z;
		19'b0111011110011010111: color_data = Z;
		19'b0111011110011011000: color_data = Z;
		19'b0111011110100001001: color_data = Z;
		19'b0111011110100001010: color_data = Z;
		19'b0111011110100001011: color_data = Z;
		19'b0111011110100010001: color_data = Z;
		19'b0111011110100010010: color_data = Z;
		19'b0111011110100010011: color_data = Z;
		19'b0111011110100010100: color_data = Z;
		19'b0111011110100011000: color_data = Z;
		19'b0111011110100011001: color_data = Z;
		19'b0111011110100011010: color_data = Z;
		19'b0111011110100011011: color_data = Z;
		19'b0111011110100011100: color_data = Z;
		19'b0111011110100011101: color_data = Z;
		19'b0111011110100011110: color_data = Z;
		19'b0111011110100011111: color_data = Z;
		19'b0111011110100100000: color_data = Z;
		19'b0111011110100100001: color_data = Z;
		19'b0111011110100100010: color_data = Z;
		19'b0111011110100100011: color_data = Z;
		19'b0111011110100100100: color_data = Z;
		19'b0111011110100100101: color_data = Z;
		19'b0111011110100101000: color_data = Z;
		19'b0111011110100101001: color_data = Z;
		19'b0111011110100101010: color_data = Z;
		19'b0111011110100101011: color_data = Z;
		19'b0111011110100101100: color_data = Z;
		19'b0111011110100101101: color_data = Z;
		19'b0111011110100101110: color_data = Z;
		19'b0111011110100101111: color_data = Z;
		19'b0111011110100110000: color_data = Z;
		19'b0111011110100110001: color_data = Z;
		19'b0111011110100110010: color_data = Z;
		19'b0111011110100110011: color_data = Z;
		19'b0111011110100110100: color_data = Z;
		19'b0111011110100110101: color_data = Z;
		19'b0111011110100110110: color_data = Z;
		19'b0111011110100110111: color_data = Z;
		19'b0111011110100111000: color_data = Z;
		19'b0111011110100111001: color_data = Z;
		19'b0111011110100111010: color_data = Z;
		19'b0111011110100111011: color_data = Z;
		19'b0111011110100111100: color_data = Z;
		19'b0111011110100111101: color_data = Z;
		19'b0111011110100111110: color_data = Z;
		19'b0111011110100111111: color_data = Z;
		19'b0111011110101000000: color_data = Z;
		19'b0111011110101000001: color_data = Z;
		19'b0111011110101000010: color_data = Z;
		19'b0111011110101000011: color_data = Z;
		19'b0111011110101000100: color_data = Z;
		19'b0111011110101000101: color_data = Z;
		19'b0111011110101000110: color_data = Z;
		19'b0111011110101000111: color_data = Z;
		19'b0111011110101001000: color_data = Z;
		19'b0111011110101001001: color_data = Z;
		19'b0111011110101001010: color_data = Z;
		19'b0111011110101001011: color_data = Z;
		19'b0111011110101001100: color_data = Z;
		19'b0111011110101001101: color_data = Z;
		19'b0111011110101001110: color_data = Z;
		19'b0111011110101001111: color_data = Z;
		19'b0111011110101010000: color_data = Z;
		19'b0111011110101010001: color_data = Z;
		19'b0111011110101010010: color_data = Z;
		19'b0111011110101010011: color_data = Z;
		19'b0111011110101010100: color_data = Z;
		19'b0111011110101010101: color_data = Z;
		19'b0111011110101010110: color_data = Z;
		19'b0111011110101010111: color_data = Z;
		19'b0111011110101011000: color_data = Z;
		19'b0111011110101011001: color_data = Z;
		19'b0111011110101011010: color_data = Z;
		19'b0111011110101011011: color_data = Z;
		19'b0111011110101011100: color_data = Z;
		19'b0111011110101011101: color_data = Z;
		19'b0111011110101011110: color_data = Z;
		19'b0111011110101011111: color_data = Z;
		19'b0111011110101100000: color_data = Z;
		19'b0111011110101100001: color_data = Z;
		19'b0111011110101100010: color_data = Z;
		19'b0111011110101100011: color_data = Z;
		19'b0111011110101100100: color_data = Z;
		19'b0111011110101100101: color_data = Z;
		19'b0111011110101100110: color_data = Z;
		19'b0111011110101100111: color_data = Z;
		19'b0111011110101101000: color_data = Z;
		19'b0111011110101101001: color_data = Z;
		19'b0111011110101101010: color_data = Z;
		19'b0111011110101101011: color_data = Z;
		19'b0111011110101101100: color_data = Z;
		19'b0111011110101101101: color_data = Z;
		19'b0111011110101101110: color_data = Z;
		19'b0111011110101101111: color_data = Z;
		19'b0111011110101110000: color_data = Z;
		19'b0111011110101110001: color_data = Z;
		19'b0111011110101110010: color_data = Z;
		19'b0111011110101110011: color_data = Z;
		19'b0111011110101110100: color_data = Z;
		19'b0111011110101110101: color_data = Z;
		19'b0111011110101110110: color_data = Z;
		19'b0111011110101110111: color_data = Z;
		19'b0111011110101111000: color_data = Z;
		19'b0111011110101111001: color_data = Z;
		19'b0111011110101111010: color_data = Z;
		19'b0111011110101111011: color_data = Z;
		19'b0111011110101111100: color_data = Z;
		19'b0111011110101111101: color_data = Z;
		19'b0111011110101111110: color_data = Z;
		19'b0111011110101111111: color_data = Z;
		19'b0111011110110000000: color_data = Z;
		19'b0111011110110000001: color_data = Z;
		19'b0111011110110000010: color_data = Z;
		19'b0111011110110000011: color_data = Z;
		19'b0111011110110000100: color_data = Z;
		19'b0111011110110000101: color_data = Z;
		19'b0111011110110000110: color_data = Z;
		19'b0111011110110000111: color_data = Z;
		19'b0111011110110001000: color_data = Z;
		19'b0111011110110001001: color_data = Z;
		19'b0111011110110001010: color_data = Z;
		19'b0111011110110001011: color_data = Z;
		19'b0111011110110010110: color_data = Z;
		19'b0111011110110010111: color_data = Z;
		19'b0111011110110011000: color_data = Z;
		19'b0111011110110011001: color_data = Z;
		19'b0111011110110011010: color_data = Z;
		19'b0111011110110011011: color_data = Z;
		19'b0111011110110011100: color_data = Z;
		19'b0111011110110011101: color_data = Z;
		19'b0111011110110011110: color_data = Z;
		19'b0111011110110011111: color_data = Z;
		19'b0111011110110100000: color_data = Z;
		19'b0111011110110100001: color_data = Z;
		19'b0111011110110100010: color_data = Z;
		19'b0111011110110100011: color_data = Z;
		19'b0111011110110100100: color_data = Z;
		19'b0111011110110100101: color_data = Z;
		19'b0111011110110100110: color_data = Z;
		19'b0111011110110100111: color_data = Z;
		19'b0111011110110101000: color_data = Z;
		19'b0111011110110101001: color_data = Z;
		19'b0111011110110101010: color_data = Z;
		19'b0111011110110101011: color_data = Z;
		19'b0111011110110101100: color_data = Z;
		19'b0111011110110101101: color_data = Z;
		19'b0111011110110101110: color_data = Z;
		19'b0111011110110101111: color_data = Z;
		19'b0111011110110110000: color_data = Z;
		19'b0111011110110110001: color_data = Z;
		19'b0111011110110110010: color_data = Z;
		19'b0111011110110110011: color_data = Z;
		19'b0111011110110110100: color_data = Z;
		19'b0111011110110110101: color_data = Z;
		19'b0111011110110110110: color_data = Z;
		19'b0111011110110110111: color_data = Z;
		19'b0111011110110111000: color_data = Z;
		19'b0111011110110111001: color_data = Z;
		19'b0111011110110111010: color_data = Z;
		19'b0111011110110111011: color_data = Z;
		19'b0111011110110111100: color_data = Z;
		19'b0111011110110111101: color_data = Z;
		19'b0111011110110111110: color_data = Z;
		19'b0111011110110111111: color_data = Z;
		19'b0111011110111000000: color_data = Z;
		19'b0111011110111000001: color_data = Z;
		19'b0111011110111000010: color_data = Z;
		19'b0111011110111000011: color_data = Z;
		19'b0111011110111000100: color_data = Z;
		19'b0111011110111000101: color_data = Z;
		19'b0111100000010101101: color_data = Z;
		19'b0111100000010101110: color_data = Z;
		19'b0111100000010101111: color_data = Z;
		19'b0111100000010110000: color_data = Z;
		19'b0111100000010110001: color_data = Z;
		19'b0111100000010110010: color_data = Z;
		19'b0111100000010110011: color_data = Z;
		19'b0111100000010110100: color_data = Z;
		19'b0111100000010110101: color_data = Z;
		19'b0111100000010110110: color_data = Z;
		19'b0111100000010110111: color_data = Z;
		19'b0111100000010111000: color_data = Z;
		19'b0111100000010111001: color_data = Z;
		19'b0111100000010111010: color_data = Z;
		19'b0111100000010111011: color_data = Z;
		19'b0111100000011000100: color_data = Z;
		19'b0111100000011000101: color_data = Z;
		19'b0111100000011000110: color_data = Z;
		19'b0111100000011000111: color_data = Z;
		19'b0111100000011001000: color_data = Z;
		19'b0111100000011001001: color_data = Z;
		19'b0111100000011001010: color_data = Z;
		19'b0111100000011001011: color_data = Z;
		19'b0111100000011001100: color_data = Z;
		19'b0111100000011001101: color_data = Z;
		19'b0111100000011001110: color_data = Z;
		19'b0111100000011001111: color_data = Z;
		19'b0111100000011010000: color_data = Z;
		19'b0111100000011010001: color_data = Z;
		19'b0111100000011010010: color_data = Z;
		19'b0111100000011010011: color_data = Z;
		19'b0111100000011010100: color_data = Z;
		19'b0111100000011010101: color_data = Z;
		19'b0111100000011010110: color_data = Z;
		19'b0111100000011010111: color_data = Z;
		19'b0111100000011011000: color_data = Z;
		19'b0111100000011011001: color_data = Z;
		19'b0111100000100001010: color_data = Z;
		19'b0111100000100001111: color_data = Z;
		19'b0111100000100010000: color_data = Z;
		19'b0111100000100010001: color_data = Z;
		19'b0111100000100010010: color_data = Z;
		19'b0111100000100010011: color_data = Z;
		19'b0111100000100010110: color_data = Z;
		19'b0111100000100011000: color_data = Z;
		19'b0111100000100011001: color_data = Z;
		19'b0111100000100011010: color_data = Z;
		19'b0111100000100011011: color_data = Z;
		19'b0111100000100011100: color_data = Z;
		19'b0111100000100011101: color_data = Z;
		19'b0111100000100011110: color_data = Z;
		19'b0111100000100011111: color_data = Z;
		19'b0111100000100100000: color_data = Z;
		19'b0111100000100100001: color_data = Z;
		19'b0111100000100100010: color_data = Z;
		19'b0111100000100100011: color_data = Z;
		19'b0111100000100100100: color_data = Z;
		19'b0111100000100100101: color_data = Z;
		19'b0111100000100101000: color_data = Z;
		19'b0111100000100101001: color_data = Z;
		19'b0111100000100101010: color_data = Z;
		19'b0111100000100101011: color_data = Z;
		19'b0111100000100101100: color_data = Z;
		19'b0111100000100101101: color_data = Z;
		19'b0111100000100101110: color_data = Z;
		19'b0111100000100101111: color_data = Z;
		19'b0111100000100110000: color_data = Z;
		19'b0111100000100110001: color_data = Z;
		19'b0111100000100110010: color_data = Z;
		19'b0111100000100110011: color_data = Z;
		19'b0111100000100110100: color_data = Z;
		19'b0111100000100110110: color_data = Z;
		19'b0111100000100110111: color_data = Z;
		19'b0111100000100111000: color_data = Z;
		19'b0111100000100111001: color_data = Z;
		19'b0111100000100111010: color_data = Z;
		19'b0111100000100111011: color_data = Z;
		19'b0111100000100111100: color_data = Z;
		19'b0111100000100111101: color_data = Z;
		19'b0111100000100111110: color_data = Z;
		19'b0111100000100111111: color_data = Z;
		19'b0111100000101000000: color_data = Z;
		19'b0111100000101000001: color_data = Z;
		19'b0111100000101000010: color_data = Z;
		19'b0111100000101000011: color_data = Z;
		19'b0111100000101000100: color_data = Z;
		19'b0111100000101000101: color_data = Z;
		19'b0111100000101000110: color_data = Z;
		19'b0111100000101000111: color_data = Z;
		19'b0111100000101001000: color_data = Z;
		19'b0111100000101001001: color_data = Z;
		19'b0111100000101001010: color_data = Z;
		19'b0111100000101001011: color_data = Z;
		19'b0111100000101001100: color_data = Z;
		19'b0111100000101001101: color_data = Z;
		19'b0111100000101001110: color_data = Z;
		19'b0111100000101001111: color_data = Z;
		19'b0111100000101010000: color_data = Z;
		19'b0111100000101010001: color_data = Z;
		19'b0111100000101010010: color_data = Z;
		19'b0111100000101010011: color_data = Z;
		19'b0111100000101010100: color_data = Z;
		19'b0111100000101010101: color_data = Z;
		19'b0111100000101010110: color_data = Z;
		19'b0111100000101010111: color_data = Z;
		19'b0111100000101011000: color_data = Z;
		19'b0111100000101011001: color_data = Z;
		19'b0111100000101011010: color_data = Z;
		19'b0111100000101011011: color_data = Z;
		19'b0111100000101011100: color_data = Z;
		19'b0111100000101011101: color_data = Z;
		19'b0111100000101011110: color_data = Z;
		19'b0111100000101011111: color_data = Z;
		19'b0111100000101100000: color_data = Z;
		19'b0111100000101100001: color_data = Z;
		19'b0111100000101100010: color_data = Z;
		19'b0111100000101100011: color_data = Z;
		19'b0111100000101100100: color_data = Z;
		19'b0111100000101100101: color_data = Z;
		19'b0111100000101100110: color_data = Z;
		19'b0111100000101100111: color_data = Z;
		19'b0111100000101101000: color_data = Z;
		19'b0111100000101101001: color_data = Z;
		19'b0111100000101101010: color_data = Z;
		19'b0111100000101101011: color_data = Z;
		19'b0111100000101101100: color_data = Z;
		19'b0111100000101101101: color_data = Z;
		19'b0111100000101101110: color_data = Z;
		19'b0111100000101101111: color_data = Z;
		19'b0111100000101110000: color_data = Z;
		19'b0111100000101110001: color_data = Z;
		19'b0111100000101110010: color_data = Z;
		19'b0111100000101110011: color_data = Z;
		19'b0111100000101110100: color_data = Z;
		19'b0111100000101110101: color_data = Z;
		19'b0111100000101110110: color_data = Z;
		19'b0111100000101110111: color_data = Z;
		19'b0111100000101111000: color_data = Z;
		19'b0111100000101111001: color_data = Z;
		19'b0111100000101111010: color_data = Z;
		19'b0111100000101111011: color_data = Z;
		19'b0111100000101111100: color_data = Z;
		19'b0111100000101111101: color_data = Z;
		19'b0111100000101111110: color_data = Z;
		19'b0111100000101111111: color_data = Z;
		19'b0111100000110000000: color_data = Z;
		19'b0111100000110000001: color_data = Z;
		19'b0111100000110000010: color_data = Z;
		19'b0111100000110000011: color_data = Z;
		19'b0111100000110000100: color_data = Z;
		19'b0111100000110000101: color_data = Z;
		19'b0111100000110000110: color_data = Z;
		19'b0111100000110000111: color_data = Z;
		19'b0111100000110001000: color_data = Z;
		19'b0111100000110001001: color_data = Z;
		19'b0111100000110001010: color_data = Z;
		19'b0111100000110001011: color_data = Z;
		19'b0111100000110001110: color_data = Z;
		19'b0111100000110001111: color_data = Z;
		19'b0111100000110010000: color_data = Z;
		19'b0111100000110011000: color_data = Z;
		19'b0111100000110011001: color_data = Z;
		19'b0111100000110011010: color_data = Z;
		19'b0111100000110011011: color_data = Z;
		19'b0111100000110011100: color_data = Z;
		19'b0111100000110011101: color_data = Z;
		19'b0111100000110011110: color_data = Z;
		19'b0111100000110011111: color_data = Z;
		19'b0111100000110100000: color_data = Z;
		19'b0111100000110100001: color_data = Z;
		19'b0111100000110100010: color_data = Z;
		19'b0111100000110100011: color_data = Z;
		19'b0111100000110100100: color_data = Z;
		19'b0111100000110100101: color_data = Z;
		19'b0111100000110100110: color_data = Z;
		19'b0111100000110100111: color_data = Z;
		19'b0111100000110101000: color_data = Z;
		19'b0111100000110101001: color_data = Z;
		19'b0111100000110101010: color_data = Z;
		19'b0111100000110101011: color_data = Z;
		19'b0111100000110101100: color_data = Z;
		19'b0111100000110101101: color_data = Z;
		19'b0111100000110101110: color_data = Z;
		19'b0111100000110101111: color_data = Z;
		19'b0111100000110110000: color_data = Z;
		19'b0111100000110110001: color_data = Z;
		19'b0111100000110110010: color_data = Z;
		19'b0111100000110110011: color_data = Z;
		19'b0111100000110110100: color_data = Z;
		19'b0111100000110110101: color_data = Z;
		19'b0111100000110110110: color_data = Z;
		19'b0111100000110110111: color_data = Z;
		19'b0111100000110111000: color_data = Z;
		19'b0111100000110111001: color_data = Z;
		19'b0111100000110111010: color_data = Z;
		19'b0111100000110111011: color_data = Z;
		19'b0111100000110111100: color_data = Z;
		19'b0111100000110111101: color_data = Z;
		19'b0111100000110111110: color_data = Z;
		19'b0111100000110111111: color_data = Z;
		19'b0111100000111000000: color_data = Z;
		19'b0111100000111000001: color_data = Z;
		19'b0111100000111000010: color_data = Z;
		19'b0111100000111000011: color_data = Z;
		19'b0111100000111000100: color_data = Z;
		19'b0111100000111000101: color_data = Z;
		19'b0111100000111000110: color_data = Z;
		19'b0111100010010101101: color_data = Z;
		19'b0111100010010101110: color_data = Z;
		19'b0111100010010101111: color_data = Z;
		19'b0111100010010110000: color_data = Z;
		19'b0111100010010110001: color_data = Z;
		19'b0111100010010110010: color_data = Z;
		19'b0111100010010110011: color_data = Z;
		19'b0111100010010110100: color_data = Z;
		19'b0111100010010110101: color_data = Z;
		19'b0111100010010110110: color_data = Z;
		19'b0111100010010110111: color_data = Z;
		19'b0111100010010111000: color_data = Z;
		19'b0111100010010111001: color_data = Z;
		19'b0111100010010111010: color_data = Z;
		19'b0111100010010111011: color_data = Z;
		19'b0111100010010111100: color_data = Z;
		19'b0111100010011000101: color_data = Z;
		19'b0111100010011000110: color_data = Z;
		19'b0111100010011000111: color_data = Z;
		19'b0111100010011001000: color_data = Z;
		19'b0111100010011001001: color_data = Z;
		19'b0111100010011001010: color_data = Z;
		19'b0111100010011001011: color_data = Z;
		19'b0111100010011001100: color_data = Z;
		19'b0111100010011001101: color_data = Z;
		19'b0111100010011001110: color_data = Z;
		19'b0111100010011001111: color_data = Z;
		19'b0111100010011010000: color_data = Z;
		19'b0111100010011010001: color_data = Z;
		19'b0111100010011010010: color_data = Z;
		19'b0111100010011010011: color_data = Z;
		19'b0111100010011010100: color_data = Z;
		19'b0111100010011010101: color_data = Z;
		19'b0111100010011010110: color_data = Z;
		19'b0111100010011010111: color_data = Z;
		19'b0111100010011011000: color_data = Z;
		19'b0111100010011011001: color_data = Z;
		19'b0111100010100000010: color_data = Z;
		19'b0111100010100000011: color_data = Z;
		19'b0111100010100001111: color_data = Z;
		19'b0111100010100010000: color_data = Z;
		19'b0111100010100010001: color_data = Z;
		19'b0111100010100010010: color_data = Z;
		19'b0111100010100010110: color_data = Z;
		19'b0111100010100010111: color_data = Z;
		19'b0111100010100011000: color_data = Z;
		19'b0111100010100011001: color_data = Z;
		19'b0111100010100011010: color_data = Z;
		19'b0111100010100011011: color_data = Z;
		19'b0111100010100011100: color_data = Z;
		19'b0111100010100011101: color_data = Z;
		19'b0111100010100011110: color_data = Z;
		19'b0111100010100011111: color_data = Z;
		19'b0111100010100100000: color_data = Z;
		19'b0111100010100100001: color_data = Z;
		19'b0111100010100100010: color_data = Z;
		19'b0111100010100100011: color_data = Z;
		19'b0111100010100100100: color_data = Z;
		19'b0111100010100100101: color_data = Z;
		19'b0111100010100101000: color_data = Z;
		19'b0111100010100101001: color_data = Z;
		19'b0111100010100101010: color_data = Z;
		19'b0111100010100101011: color_data = Z;
		19'b0111100010100101100: color_data = Z;
		19'b0111100010100101101: color_data = Z;
		19'b0111100010100101110: color_data = Z;
		19'b0111100010100101111: color_data = Z;
		19'b0111100010100110000: color_data = Z;
		19'b0111100010100110001: color_data = Z;
		19'b0111100010100110010: color_data = Z;
		19'b0111100010100110011: color_data = Z;
		19'b0111100010100110111: color_data = Z;
		19'b0111100010100111000: color_data = Z;
		19'b0111100010100111001: color_data = Z;
		19'b0111100010100111010: color_data = Z;
		19'b0111100010100111011: color_data = Z;
		19'b0111100010100111100: color_data = Z;
		19'b0111100010100111101: color_data = Z;
		19'b0111100010100111110: color_data = Z;
		19'b0111100010100111111: color_data = Z;
		19'b0111100010101000000: color_data = Z;
		19'b0111100010101000001: color_data = Z;
		19'b0111100010101000010: color_data = Z;
		19'b0111100010101000011: color_data = Z;
		19'b0111100010101000100: color_data = Z;
		19'b0111100010101000101: color_data = Z;
		19'b0111100010101000110: color_data = Z;
		19'b0111100010101000111: color_data = Z;
		19'b0111100010101001000: color_data = Z;
		19'b0111100010101001001: color_data = Z;
		19'b0111100010101001010: color_data = Z;
		19'b0111100010101001011: color_data = Z;
		19'b0111100010101001100: color_data = Z;
		19'b0111100010101001101: color_data = Z;
		19'b0111100010101001110: color_data = Z;
		19'b0111100010101001111: color_data = Z;
		19'b0111100010101010000: color_data = Z;
		19'b0111100010101010001: color_data = Z;
		19'b0111100010101010010: color_data = Z;
		19'b0111100010101010011: color_data = Z;
		19'b0111100010101010100: color_data = Z;
		19'b0111100010101010101: color_data = Z;
		19'b0111100010101010110: color_data = Z;
		19'b0111100010101010111: color_data = Z;
		19'b0111100010101011000: color_data = Z;
		19'b0111100010101011001: color_data = Z;
		19'b0111100010101011010: color_data = Z;
		19'b0111100010101011011: color_data = Z;
		19'b0111100010101011100: color_data = Z;
		19'b0111100010101011101: color_data = Z;
		19'b0111100010101011110: color_data = Z;
		19'b0111100010101011111: color_data = Z;
		19'b0111100010101100000: color_data = Z;
		19'b0111100010101100001: color_data = Z;
		19'b0111100010101100011: color_data = Z;
		19'b0111100010101100100: color_data = Z;
		19'b0111100010101100101: color_data = Z;
		19'b0111100010101100110: color_data = Z;
		19'b0111100010101100111: color_data = Z;
		19'b0111100010101101000: color_data = Z;
		19'b0111100010101101001: color_data = Z;
		19'b0111100010101101010: color_data = Z;
		19'b0111100010101101011: color_data = Z;
		19'b0111100010101101100: color_data = Z;
		19'b0111100010101101101: color_data = Z;
		19'b0111100010101101110: color_data = Z;
		19'b0111100010101101111: color_data = Z;
		19'b0111100010101110000: color_data = Z;
		19'b0111100010101110001: color_data = Z;
		19'b0111100010101110010: color_data = Z;
		19'b0111100010101110011: color_data = Z;
		19'b0111100010101110100: color_data = Z;
		19'b0111100010101110101: color_data = Z;
		19'b0111100010101110110: color_data = Z;
		19'b0111100010101110111: color_data = Z;
		19'b0111100010101111000: color_data = Z;
		19'b0111100010101111001: color_data = Z;
		19'b0111100010101111010: color_data = Z;
		19'b0111100010101111011: color_data = Z;
		19'b0111100010101111100: color_data = Z;
		19'b0111100010101111101: color_data = Z;
		19'b0111100010101111110: color_data = Z;
		19'b0111100010101111111: color_data = Z;
		19'b0111100010110000000: color_data = Z;
		19'b0111100010110000001: color_data = Z;
		19'b0111100010110000010: color_data = Z;
		19'b0111100010110000011: color_data = Z;
		19'b0111100010110000100: color_data = Z;
		19'b0111100010110000101: color_data = Z;
		19'b0111100010110000110: color_data = Z;
		19'b0111100010110000111: color_data = Z;
		19'b0111100010110001000: color_data = Z;
		19'b0111100010110001001: color_data = Z;
		19'b0111100010110001010: color_data = Z;
		19'b0111100010110001011: color_data = Z;
		19'b0111100010110001100: color_data = Z;
		19'b0111100010110001110: color_data = Z;
		19'b0111100010110001111: color_data = Z;
		19'b0111100010110010000: color_data = Z;
		19'b0111100010110011010: color_data = Z;
		19'b0111100010110011011: color_data = Z;
		19'b0111100010110011100: color_data = Z;
		19'b0111100010110011101: color_data = Z;
		19'b0111100010110011110: color_data = Z;
		19'b0111100010110011111: color_data = Z;
		19'b0111100010110100000: color_data = Z;
		19'b0111100010110100001: color_data = Z;
		19'b0111100010110100010: color_data = Z;
		19'b0111100010110100011: color_data = Z;
		19'b0111100010110100100: color_data = Z;
		19'b0111100010110100101: color_data = Z;
		19'b0111100010110100110: color_data = Z;
		19'b0111100010110100111: color_data = Z;
		19'b0111100010110101000: color_data = Z;
		19'b0111100010110101001: color_data = Z;
		19'b0111100010110101010: color_data = Z;
		19'b0111100010110101011: color_data = Z;
		19'b0111100010110101100: color_data = Z;
		19'b0111100010110101101: color_data = Z;
		19'b0111100010110101110: color_data = Z;
		19'b0111100010110101111: color_data = Z;
		19'b0111100010110110000: color_data = Z;
		19'b0111100010110110001: color_data = Z;
		19'b0111100010110110010: color_data = Z;
		19'b0111100010110110011: color_data = Z;
		19'b0111100010110110100: color_data = Z;
		19'b0111100010110110101: color_data = Z;
		19'b0111100010110110110: color_data = Z;
		19'b0111100010110111000: color_data = Z;
		19'b0111100010110111001: color_data = Z;
		19'b0111100010110111010: color_data = Z;
		19'b0111100010110111011: color_data = Z;
		19'b0111100010110111100: color_data = Z;
		19'b0111100010110111101: color_data = Z;
		19'b0111100010110111110: color_data = Z;
		19'b0111100010110111111: color_data = Z;
		19'b0111100010111000000: color_data = Z;
		19'b0111100010111000001: color_data = Z;
		19'b0111100010111000010: color_data = Z;
		19'b0111100010111000011: color_data = Z;
		19'b0111100010111000100: color_data = Z;
		19'b0111100010111000101: color_data = Z;
		19'b0111100010111000110: color_data = Z;
		19'b0111100010111000111: color_data = Z;
		19'b0111100100010101110: color_data = Z;
		19'b0111100100010101111: color_data = Z;
		19'b0111100100010110000: color_data = Z;
		19'b0111100100010110001: color_data = Z;
		19'b0111100100010110010: color_data = Z;
		19'b0111100100010110011: color_data = Z;
		19'b0111100100010110100: color_data = Z;
		19'b0111100100010110101: color_data = Z;
		19'b0111100100010110110: color_data = Z;
		19'b0111100100010110111: color_data = Z;
		19'b0111100100010111000: color_data = Z;
		19'b0111100100010111001: color_data = Z;
		19'b0111100100010111010: color_data = Z;
		19'b0111100100010111011: color_data = Z;
		19'b0111100100010111100: color_data = Z;
		19'b0111100100011000110: color_data = Z;
		19'b0111100100011000111: color_data = Z;
		19'b0111100100011001000: color_data = Z;
		19'b0111100100011001001: color_data = Z;
		19'b0111100100011001010: color_data = Z;
		19'b0111100100011001011: color_data = Z;
		19'b0111100100011001100: color_data = Z;
		19'b0111100100011001101: color_data = Z;
		19'b0111100100011001110: color_data = Z;
		19'b0111100100011001111: color_data = Z;
		19'b0111100100011010000: color_data = Z;
		19'b0111100100011010001: color_data = Z;
		19'b0111100100011010010: color_data = Z;
		19'b0111100100011010011: color_data = Z;
		19'b0111100100011010100: color_data = Z;
		19'b0111100100011010101: color_data = Z;
		19'b0111100100011010110: color_data = Z;
		19'b0111100100011010111: color_data = Z;
		19'b0111100100011011000: color_data = Z;
		19'b0111100100011011001: color_data = Z;
		19'b0111100100100000000: color_data = Z;
		19'b0111100100100000001: color_data = Z;
		19'b0111100100100000010: color_data = Z;
		19'b0111100100100000011: color_data = Z;
		19'b0111100100100000100: color_data = Z;
		19'b0111100100100000101: color_data = Z;
		19'b0111100100100001110: color_data = Z;
		19'b0111100100100001111: color_data = Z;
		19'b0111100100100010000: color_data = Z;
		19'b0111100100100010001: color_data = Z;
		19'b0111100100100010010: color_data = Z;
		19'b0111100100100010101: color_data = Z;
		19'b0111100100100010110: color_data = Z;
		19'b0111100100100010111: color_data = Z;
		19'b0111100100100011000: color_data = Z;
		19'b0111100100100011001: color_data = Z;
		19'b0111100100100011010: color_data = Z;
		19'b0111100100100011011: color_data = Z;
		19'b0111100100100011100: color_data = Z;
		19'b0111100100100011101: color_data = Z;
		19'b0111100100100011110: color_data = Z;
		19'b0111100100100011111: color_data = Z;
		19'b0111100100100100000: color_data = Z;
		19'b0111100100100100001: color_data = Z;
		19'b0111100100100100010: color_data = Z;
		19'b0111100100100100011: color_data = Z;
		19'b0111100100100100100: color_data = Z;
		19'b0111100100100100101: color_data = Z;
		19'b0111100100100100110: color_data = Z;
		19'b0111100100100100111: color_data = Z;
		19'b0111100100100101000: color_data = Z;
		19'b0111100100100101001: color_data = Z;
		19'b0111100100100101010: color_data = Z;
		19'b0111100100100101011: color_data = Z;
		19'b0111100100100101100: color_data = Z;
		19'b0111100100100101101: color_data = Z;
		19'b0111100100100101110: color_data = Z;
		19'b0111100100100101111: color_data = Z;
		19'b0111100100100110000: color_data = Z;
		19'b0111100100100110001: color_data = Z;
		19'b0111100100100110010: color_data = Z;
		19'b0111100100100110111: color_data = Z;
		19'b0111100100100111000: color_data = Z;
		19'b0111100100100111001: color_data = Z;
		19'b0111100100100111010: color_data = Z;
		19'b0111100100100111011: color_data = Z;
		19'b0111100100100111100: color_data = Z;
		19'b0111100100100111101: color_data = Z;
		19'b0111100100100111110: color_data = Z;
		19'b0111100100100111111: color_data = Z;
		19'b0111100100101000000: color_data = Z;
		19'b0111100100101000001: color_data = Z;
		19'b0111100100101000010: color_data = Z;
		19'b0111100100101000011: color_data = Z;
		19'b0111100100101000100: color_data = Z;
		19'b0111100100101000101: color_data = Z;
		19'b0111100100101000110: color_data = Z;
		19'b0111100100101000111: color_data = Z;
		19'b0111100100101001000: color_data = Z;
		19'b0111100100101001001: color_data = Z;
		19'b0111100100101001010: color_data = Z;
		19'b0111100100101001011: color_data = Z;
		19'b0111100100101001100: color_data = Z;
		19'b0111100100101001101: color_data = Z;
		19'b0111100100101001110: color_data = Z;
		19'b0111100100101001111: color_data = Z;
		19'b0111100100101010000: color_data = Z;
		19'b0111100100101010001: color_data = Z;
		19'b0111100100101010010: color_data = Z;
		19'b0111100100101010011: color_data = Z;
		19'b0111100100101010100: color_data = Z;
		19'b0111100100101010101: color_data = Z;
		19'b0111100100101010110: color_data = Z;
		19'b0111100100101010111: color_data = Z;
		19'b0111100100101011000: color_data = Z;
		19'b0111100100101011001: color_data = Z;
		19'b0111100100101011010: color_data = Z;
		19'b0111100100101011011: color_data = Z;
		19'b0111100100101011100: color_data = Z;
		19'b0111100100101011101: color_data = Z;
		19'b0111100100101011110: color_data = Z;
		19'b0111100100101011111: color_data = Z;
		19'b0111100100101100000: color_data = Z;
		19'b0111100100101100001: color_data = Z;
		19'b0111100100101100010: color_data = Z;
		19'b0111100100101100100: color_data = Z;
		19'b0111100100101100101: color_data = Z;
		19'b0111100100101100110: color_data = Z;
		19'b0111100100101100111: color_data = Z;
		19'b0111100100101101000: color_data = Z;
		19'b0111100100101101001: color_data = Z;
		19'b0111100100101101010: color_data = Z;
		19'b0111100100101101011: color_data = Z;
		19'b0111100100101101100: color_data = Z;
		19'b0111100100101101101: color_data = Z;
		19'b0111100100101101110: color_data = Z;
		19'b0111100100101101111: color_data = Z;
		19'b0111100100101110000: color_data = Z;
		19'b0111100100101110001: color_data = Z;
		19'b0111100100101110010: color_data = Z;
		19'b0111100100101110011: color_data = Z;
		19'b0111100100101110100: color_data = Z;
		19'b0111100100101110101: color_data = Z;
		19'b0111100100101110110: color_data = Z;
		19'b0111100100101110111: color_data = Z;
		19'b0111100100101111000: color_data = Z;
		19'b0111100100101111001: color_data = Z;
		19'b0111100100101111010: color_data = Z;
		19'b0111100100101111011: color_data = Z;
		19'b0111100100101111100: color_data = Z;
		19'b0111100100101111101: color_data = Z;
		19'b0111100100101111110: color_data = Z;
		19'b0111100100101111111: color_data = Z;
		19'b0111100100110000000: color_data = Z;
		19'b0111100100110000001: color_data = Z;
		19'b0111100100110000010: color_data = Z;
		19'b0111100100110000011: color_data = Z;
		19'b0111100100110000100: color_data = Z;
		19'b0111100100110000101: color_data = Z;
		19'b0111100100110000110: color_data = Z;
		19'b0111100100110000111: color_data = Z;
		19'b0111100100110001000: color_data = Z;
		19'b0111100100110001001: color_data = Z;
		19'b0111100100110001010: color_data = Z;
		19'b0111100100110001011: color_data = Z;
		19'b0111100100110001100: color_data = Z;
		19'b0111100100110001110: color_data = Z;
		19'b0111100100110001111: color_data = Z;
		19'b0111100100110010000: color_data = Z;
		19'b0111100100110010001: color_data = Z;
		19'b0111100100110010100: color_data = Z;
		19'b0111100100110010101: color_data = Z;
		19'b0111100100110011101: color_data = Z;
		19'b0111100100110011110: color_data = Z;
		19'b0111100100110011111: color_data = Z;
		19'b0111100100110100000: color_data = Z;
		19'b0111100100110100001: color_data = Z;
		19'b0111100100110100010: color_data = Z;
		19'b0111100100110100011: color_data = Z;
		19'b0111100100110100100: color_data = Z;
		19'b0111100100110100101: color_data = Z;
		19'b0111100100110100110: color_data = Z;
		19'b0111100100110100111: color_data = Z;
		19'b0111100100110101000: color_data = Z;
		19'b0111100100110101001: color_data = Z;
		19'b0111100100110101010: color_data = Z;
		19'b0111100100110101011: color_data = Z;
		19'b0111100100110101100: color_data = Z;
		19'b0111100100110101101: color_data = Z;
		19'b0111100100110101110: color_data = Z;
		19'b0111100100110101111: color_data = Z;
		19'b0111100100110110000: color_data = Z;
		19'b0111100100110110001: color_data = Z;
		19'b0111100100110110010: color_data = Z;
		19'b0111100100110110011: color_data = Z;
		19'b0111100100110110100: color_data = Z;
		19'b0111100100110110101: color_data = Z;
		19'b0111100100110110110: color_data = Z;
		19'b0111100100110111001: color_data = Z;
		19'b0111100100110111010: color_data = Z;
		19'b0111100100110111011: color_data = Z;
		19'b0111100100110111100: color_data = Z;
		19'b0111100100110111101: color_data = Z;
		19'b0111100100110111110: color_data = Z;
		19'b0111100100110111111: color_data = Z;
		19'b0111100100111000000: color_data = Z;
		19'b0111100100111000001: color_data = Z;
		19'b0111100100111000010: color_data = Z;
		19'b0111100100111000011: color_data = Z;
		19'b0111100100111000100: color_data = Z;
		19'b0111100100111000101: color_data = Z;
		19'b0111100100111000110: color_data = Z;
		19'b0111100100111000111: color_data = Z;
		19'b0111100110010101110: color_data = Z;
		19'b0111100110010101111: color_data = Z;
		19'b0111100110010110000: color_data = Z;
		19'b0111100110010110001: color_data = Z;
		19'b0111100110010110010: color_data = Z;
		19'b0111100110010110011: color_data = Z;
		19'b0111100110010110100: color_data = Z;
		19'b0111100110010110101: color_data = Z;
		19'b0111100110010110110: color_data = Z;
		19'b0111100110010110111: color_data = Z;
		19'b0111100110010111000: color_data = Z;
		19'b0111100110010111001: color_data = Z;
		19'b0111100110010111010: color_data = Z;
		19'b0111100110010111011: color_data = Z;
		19'b0111100110010111100: color_data = Z;
		19'b0111100110010111101: color_data = Z;
		19'b0111100110011000111: color_data = Z;
		19'b0111100110011001000: color_data = Z;
		19'b0111100110011001001: color_data = Z;
		19'b0111100110011001010: color_data = Z;
		19'b0111100110011001011: color_data = Z;
		19'b0111100110011001100: color_data = Z;
		19'b0111100110011001101: color_data = Z;
		19'b0111100110011001110: color_data = Z;
		19'b0111100110011001111: color_data = Z;
		19'b0111100110011010000: color_data = Z;
		19'b0111100110011010001: color_data = Z;
		19'b0111100110011010010: color_data = Z;
		19'b0111100110011010011: color_data = Z;
		19'b0111100110011010100: color_data = Z;
		19'b0111100110011010101: color_data = Z;
		19'b0111100110011010110: color_data = Z;
		19'b0111100110011010111: color_data = Z;
		19'b0111100110011011000: color_data = Z;
		19'b0111100110011011001: color_data = Z;
		19'b0111100110011011010: color_data = Z;
		19'b0111100110011111101: color_data = Z;
		19'b0111100110011111110: color_data = Z;
		19'b0111100110011111111: color_data = Z;
		19'b0111100110100000000: color_data = Z;
		19'b0111100110100000001: color_data = Z;
		19'b0111100110100000010: color_data = Z;
		19'b0111100110100000011: color_data = Z;
		19'b0111100110100000100: color_data = Z;
		19'b0111100110100000101: color_data = Z;
		19'b0111100110100001111: color_data = Z;
		19'b0111100110100010000: color_data = Z;
		19'b0111100110100010001: color_data = Z;
		19'b0111100110100010100: color_data = Z;
		19'b0111100110100010101: color_data = Z;
		19'b0111100110100010110: color_data = Z;
		19'b0111100110100010111: color_data = Z;
		19'b0111100110100011000: color_data = Z;
		19'b0111100110100011001: color_data = Z;
		19'b0111100110100011010: color_data = Z;
		19'b0111100110100011011: color_data = Z;
		19'b0111100110100011100: color_data = Z;
		19'b0111100110100011101: color_data = Z;
		19'b0111100110100011110: color_data = Z;
		19'b0111100110100011111: color_data = Z;
		19'b0111100110100100000: color_data = Z;
		19'b0111100110100100001: color_data = Z;
		19'b0111100110100100010: color_data = Z;
		19'b0111100110100100011: color_data = Z;
		19'b0111100110100100100: color_data = Z;
		19'b0111100110100100101: color_data = Z;
		19'b0111100110100100110: color_data = Z;
		19'b0111100110100100111: color_data = Z;
		19'b0111100110100101000: color_data = Z;
		19'b0111100110100101001: color_data = Z;
		19'b0111100110100101010: color_data = Z;
		19'b0111100110100101011: color_data = Z;
		19'b0111100110100101100: color_data = Z;
		19'b0111100110100101101: color_data = Z;
		19'b0111100110100101110: color_data = Z;
		19'b0111100110100101111: color_data = Z;
		19'b0111100110100110000: color_data = Z;
		19'b0111100110100110001: color_data = Z;
		19'b0111100110100110111: color_data = Z;
		19'b0111100110100111000: color_data = Z;
		19'b0111100110100111001: color_data = Z;
		19'b0111100110100111010: color_data = Z;
		19'b0111100110100111011: color_data = Z;
		19'b0111100110100111100: color_data = Z;
		19'b0111100110100111101: color_data = Z;
		19'b0111100110100111110: color_data = Z;
		19'b0111100110100111111: color_data = Z;
		19'b0111100110101000000: color_data = Z;
		19'b0111100110101000001: color_data = Z;
		19'b0111100110101000010: color_data = Z;
		19'b0111100110101000011: color_data = Z;
		19'b0111100110101000100: color_data = Z;
		19'b0111100110101000101: color_data = Z;
		19'b0111100110101000110: color_data = Z;
		19'b0111100110101000111: color_data = Z;
		19'b0111100110101001000: color_data = Z;
		19'b0111100110101001001: color_data = Z;
		19'b0111100110101001010: color_data = Z;
		19'b0111100110101001011: color_data = Z;
		19'b0111100110101001100: color_data = Z;
		19'b0111100110101001101: color_data = Z;
		19'b0111100110101001110: color_data = Z;
		19'b0111100110101001111: color_data = Z;
		19'b0111100110101010000: color_data = Z;
		19'b0111100110101010001: color_data = Z;
		19'b0111100110101010010: color_data = Z;
		19'b0111100110101010011: color_data = Z;
		19'b0111100110101010100: color_data = Z;
		19'b0111100110101010101: color_data = Z;
		19'b0111100110101010110: color_data = Z;
		19'b0111100110101010111: color_data = Z;
		19'b0111100110101011000: color_data = Z;
		19'b0111100110101011001: color_data = Z;
		19'b0111100110101011010: color_data = Z;
		19'b0111100110101011011: color_data = Z;
		19'b0111100110101011100: color_data = Z;
		19'b0111100110101011101: color_data = Z;
		19'b0111100110101011110: color_data = Z;
		19'b0111100110101011111: color_data = Z;
		19'b0111100110101100000: color_data = Z;
		19'b0111100110101100001: color_data = Z;
		19'b0111100110101100010: color_data = Z;
		19'b0111100110101100100: color_data = Z;
		19'b0111100110101100101: color_data = Z;
		19'b0111100110101100110: color_data = Z;
		19'b0111100110101100111: color_data = Z;
		19'b0111100110101101000: color_data = Z;
		19'b0111100110101101001: color_data = Z;
		19'b0111100110101101010: color_data = Z;
		19'b0111100110101101011: color_data = Z;
		19'b0111100110101101100: color_data = Z;
		19'b0111100110101101101: color_data = Z;
		19'b0111100110101101110: color_data = Z;
		19'b0111100110101101111: color_data = Z;
		19'b0111100110101110000: color_data = Z;
		19'b0111100110101110001: color_data = Z;
		19'b0111100110101110010: color_data = Z;
		19'b0111100110101110011: color_data = Z;
		19'b0111100110101110100: color_data = Z;
		19'b0111100110101110101: color_data = Z;
		19'b0111100110101110110: color_data = Z;
		19'b0111100110101110111: color_data = Z;
		19'b0111100110101111000: color_data = Z;
		19'b0111100110101111001: color_data = Z;
		19'b0111100110101111010: color_data = Z;
		19'b0111100110101111011: color_data = Z;
		19'b0111100110101111100: color_data = Z;
		19'b0111100110101111101: color_data = Z;
		19'b0111100110101111110: color_data = Z;
		19'b0111100110101111111: color_data = Z;
		19'b0111100110110000000: color_data = Z;
		19'b0111100110110000001: color_data = Z;
		19'b0111100110110000010: color_data = Z;
		19'b0111100110110000011: color_data = Z;
		19'b0111100110110000100: color_data = Z;
		19'b0111100110110000101: color_data = Z;
		19'b0111100110110000110: color_data = Z;
		19'b0111100110110000111: color_data = Z;
		19'b0111100110110001000: color_data = Z;
		19'b0111100110110001001: color_data = Z;
		19'b0111100110110001010: color_data = Z;
		19'b0111100110110001011: color_data = Z;
		19'b0111100110110001110: color_data = Z;
		19'b0111100110110001111: color_data = Z;
		19'b0111100110110010000: color_data = Z;
		19'b0111100110110010001: color_data = Z;
		19'b0111100110110010110: color_data = Z;
		19'b0111100110110010111: color_data = Z;
		19'b0111100110110011000: color_data = Z;
		19'b0111100110110100000: color_data = Z;
		19'b0111100110110100001: color_data = Z;
		19'b0111100110110100010: color_data = Z;
		19'b0111100110110100011: color_data = Z;
		19'b0111100110110100100: color_data = Z;
		19'b0111100110110100101: color_data = Z;
		19'b0111100110110100110: color_data = Z;
		19'b0111100110110100111: color_data = Z;
		19'b0111100110110101000: color_data = Z;
		19'b0111100110110101001: color_data = Z;
		19'b0111100110110101010: color_data = Z;
		19'b0111100110110101011: color_data = Z;
		19'b0111100110110101100: color_data = Z;
		19'b0111100110110101101: color_data = Z;
		19'b0111100110110101110: color_data = Z;
		19'b0111100110110101111: color_data = Z;
		19'b0111100110110110000: color_data = Z;
		19'b0111100110110110001: color_data = Z;
		19'b0111100110110110010: color_data = Z;
		19'b0111100110110110011: color_data = Z;
		19'b0111100110110110100: color_data = Z;
		19'b0111100110110110101: color_data = Z;
		19'b0111100110110110110: color_data = Z;
		19'b0111100110110110111: color_data = Z;
		19'b0111100110110111001: color_data = Z;
		19'b0111100110110111010: color_data = Z;
		19'b0111100110110111011: color_data = Z;
		19'b0111100110110111100: color_data = Z;
		19'b0111100110110111101: color_data = Z;
		19'b0111100110110111110: color_data = Z;
		19'b0111100110110111111: color_data = Z;
		19'b0111100110111000000: color_data = Z;
		19'b0111100110111000001: color_data = Z;
		19'b0111100110111000010: color_data = Z;
		19'b0111100110111000011: color_data = Z;
		19'b0111100110111000100: color_data = Z;
		19'b0111100110111000101: color_data = Z;
		19'b0111100110111000110: color_data = Z;
		19'b0111100110111000111: color_data = Z;
		19'b0111100110111001000: color_data = Z;
		19'b0111101000010101110: color_data = Z;
		19'b0111101000010101111: color_data = Z;
		19'b0111101000010110000: color_data = Z;
		19'b0111101000010110001: color_data = Z;
		19'b0111101000010110010: color_data = Z;
		19'b0111101000010110011: color_data = Z;
		19'b0111101000010110100: color_data = Z;
		19'b0111101000010110101: color_data = Z;
		19'b0111101000010110110: color_data = Z;
		19'b0111101000010110111: color_data = Z;
		19'b0111101000010111000: color_data = Z;
		19'b0111101000010111001: color_data = Z;
		19'b0111101000010111010: color_data = Z;
		19'b0111101000010111011: color_data = Z;
		19'b0111101000010111100: color_data = Z;
		19'b0111101000010111101: color_data = Z;
		19'b0111101000010111110: color_data = Z;
		19'b0111101000011001000: color_data = Z;
		19'b0111101000011001001: color_data = Z;
		19'b0111101000011001010: color_data = Z;
		19'b0111101000011001011: color_data = Z;
		19'b0111101000011001100: color_data = Z;
		19'b0111101000011001101: color_data = Z;
		19'b0111101000011001110: color_data = Z;
		19'b0111101000011001111: color_data = Z;
		19'b0111101000011010000: color_data = Z;
		19'b0111101000011010001: color_data = Z;
		19'b0111101000011010010: color_data = Z;
		19'b0111101000011010011: color_data = Z;
		19'b0111101000011010100: color_data = Z;
		19'b0111101000011010101: color_data = Z;
		19'b0111101000011010110: color_data = Z;
		19'b0111101000011010111: color_data = Z;
		19'b0111101000011011000: color_data = Z;
		19'b0111101000011011001: color_data = Z;
		19'b0111101000011011010: color_data = Z;
		19'b0111101000011011011: color_data = Z;
		19'b0111101000011011100: color_data = Z;
		19'b0111101000011110011: color_data = Z;
		19'b0111101000011110100: color_data = Z;
		19'b0111101000011110101: color_data = Z;
		19'b0111101000011110110: color_data = Z;
		19'b0111101000011110111: color_data = Z;
		19'b0111101000011111001: color_data = Z;
		19'b0111101000011111010: color_data = Z;
		19'b0111101000011111011: color_data = Z;
		19'b0111101000011111100: color_data = Z;
		19'b0111101000011111101: color_data = Z;
		19'b0111101000011111110: color_data = Z;
		19'b0111101000011111111: color_data = Z;
		19'b0111101000100000000: color_data = Z;
		19'b0111101000100000001: color_data = Z;
		19'b0111101000100000010: color_data = Z;
		19'b0111101000100000011: color_data = Z;
		19'b0111101000100000100: color_data = Z;
		19'b0111101000100000101: color_data = Z;
		19'b0111101000100001110: color_data = Z;
		19'b0111101000100001111: color_data = Z;
		19'b0111101000100010000: color_data = Z;
		19'b0111101000100010011: color_data = Z;
		19'b0111101000100010100: color_data = Z;
		19'b0111101000100010101: color_data = Z;
		19'b0111101000100010110: color_data = Z;
		19'b0111101000100010111: color_data = Z;
		19'b0111101000100011000: color_data = Z;
		19'b0111101000100011001: color_data = Z;
		19'b0111101000100011010: color_data = Z;
		19'b0111101000100011011: color_data = Z;
		19'b0111101000100011100: color_data = Z;
		19'b0111101000100011101: color_data = Z;
		19'b0111101000100011110: color_data = Z;
		19'b0111101000100011111: color_data = Z;
		19'b0111101000100100000: color_data = Z;
		19'b0111101000100100001: color_data = Z;
		19'b0111101000100100010: color_data = Z;
		19'b0111101000100100011: color_data = Z;
		19'b0111101000100100100: color_data = Z;
		19'b0111101000100100101: color_data = Z;
		19'b0111101000100100110: color_data = Z;
		19'b0111101000100100111: color_data = Z;
		19'b0111101000100101000: color_data = Z;
		19'b0111101000100101001: color_data = Z;
		19'b0111101000100101010: color_data = Z;
		19'b0111101000100101011: color_data = Z;
		19'b0111101000100101100: color_data = Z;
		19'b0111101000100101101: color_data = Z;
		19'b0111101000100101110: color_data = Z;
		19'b0111101000100101111: color_data = Z;
		19'b0111101000100110000: color_data = Z;
		19'b0111101000100110001: color_data = Z;
		19'b0111101000100110110: color_data = Z;
		19'b0111101000100110111: color_data = Z;
		19'b0111101000100111000: color_data = Z;
		19'b0111101000100111001: color_data = Z;
		19'b0111101000100111010: color_data = Z;
		19'b0111101000100111011: color_data = Z;
		19'b0111101000100111100: color_data = Z;
		19'b0111101000100111101: color_data = Z;
		19'b0111101000100111110: color_data = Z;
		19'b0111101000100111111: color_data = Z;
		19'b0111101000101000000: color_data = Z;
		19'b0111101000101000001: color_data = Z;
		19'b0111101000101000010: color_data = Z;
		19'b0111101000101000011: color_data = Z;
		19'b0111101000101000100: color_data = Z;
		19'b0111101000101000101: color_data = Z;
		19'b0111101000101000110: color_data = Z;
		19'b0111101000101000111: color_data = Z;
		19'b0111101000101001000: color_data = Z;
		19'b0111101000101001001: color_data = Z;
		19'b0111101000101001010: color_data = Z;
		19'b0111101000101001011: color_data = Z;
		19'b0111101000101001100: color_data = Z;
		19'b0111101000101001101: color_data = Z;
		19'b0111101000101001110: color_data = Z;
		19'b0111101000101001111: color_data = Z;
		19'b0111101000101010000: color_data = Z;
		19'b0111101000101010001: color_data = Z;
		19'b0111101000101010010: color_data = Z;
		19'b0111101000101010011: color_data = Z;
		19'b0111101000101010100: color_data = Z;
		19'b0111101000101010101: color_data = Z;
		19'b0111101000101010110: color_data = Z;
		19'b0111101000101010111: color_data = Z;
		19'b0111101000101011000: color_data = Z;
		19'b0111101000101011001: color_data = Z;
		19'b0111101000101011010: color_data = Z;
		19'b0111101000101011011: color_data = Z;
		19'b0111101000101011100: color_data = Z;
		19'b0111101000101011101: color_data = Z;
		19'b0111101000101011110: color_data = Z;
		19'b0111101000101011111: color_data = Z;
		19'b0111101000101100000: color_data = Z;
		19'b0111101000101100001: color_data = Z;
		19'b0111101000101100010: color_data = Z;
		19'b0111101000101100011: color_data = Z;
		19'b0111101000101100101: color_data = Z;
		19'b0111101000101100110: color_data = Z;
		19'b0111101000101100111: color_data = Z;
		19'b0111101000101101000: color_data = Z;
		19'b0111101000101101001: color_data = Z;
		19'b0111101000101101010: color_data = Z;
		19'b0111101000101101011: color_data = Z;
		19'b0111101000101101100: color_data = Z;
		19'b0111101000101101101: color_data = Z;
		19'b0111101000101101110: color_data = Z;
		19'b0111101000101101111: color_data = Z;
		19'b0111101000101110000: color_data = Z;
		19'b0111101000101110001: color_data = Z;
		19'b0111101000101110010: color_data = Z;
		19'b0111101000101110011: color_data = Z;
		19'b0111101000101110100: color_data = Z;
		19'b0111101000101110101: color_data = Z;
		19'b0111101000101110110: color_data = Z;
		19'b0111101000101110111: color_data = Z;
		19'b0111101000101111000: color_data = Z;
		19'b0111101000101111001: color_data = Z;
		19'b0111101000101111010: color_data = Z;
		19'b0111101000101111011: color_data = Z;
		19'b0111101000101111100: color_data = Z;
		19'b0111101000101111101: color_data = Z;
		19'b0111101000101111110: color_data = Z;
		19'b0111101000101111111: color_data = Z;
		19'b0111101000110000000: color_data = Z;
		19'b0111101000110000001: color_data = Z;
		19'b0111101000110000010: color_data = Z;
		19'b0111101000110000011: color_data = Z;
		19'b0111101000110000100: color_data = Z;
		19'b0111101000110000101: color_data = Z;
		19'b0111101000110000110: color_data = Z;
		19'b0111101000110000111: color_data = Z;
		19'b0111101000110001000: color_data = Z;
		19'b0111101000110001001: color_data = Z;
		19'b0111101000110001010: color_data = Z;
		19'b0111101000110001110: color_data = Z;
		19'b0111101000110001111: color_data = Z;
		19'b0111101000110010000: color_data = Z;
		19'b0111101000110010001: color_data = Z;
		19'b0111101000110010010: color_data = Z;
		19'b0111101000110011000: color_data = Z;
		19'b0111101000110011001: color_data = Z;
		19'b0111101000110011010: color_data = Z;
		19'b0111101000110011011: color_data = Z;
		19'b0111101000110100111: color_data = Z;
		19'b0111101000110101000: color_data = Z;
		19'b0111101000110101001: color_data = Z;
		19'b0111101000110101010: color_data = Z;
		19'b0111101000110101011: color_data = Z;
		19'b0111101000110101100: color_data = Z;
		19'b0111101000110101101: color_data = Z;
		19'b0111101000110101110: color_data = Z;
		19'b0111101000110101111: color_data = Z;
		19'b0111101000110110000: color_data = Z;
		19'b0111101000110110001: color_data = Z;
		19'b0111101000110110010: color_data = Z;
		19'b0111101000110110011: color_data = Z;
		19'b0111101000110110100: color_data = Z;
		19'b0111101000110110101: color_data = Z;
		19'b0111101000110110110: color_data = Z;
		19'b0111101000110110111: color_data = Z;
		19'b0111101000110111000: color_data = Z;
		19'b0111101000110111010: color_data = Z;
		19'b0111101000110111011: color_data = Z;
		19'b0111101000110111100: color_data = Z;
		19'b0111101000110111101: color_data = Z;
		19'b0111101000110111110: color_data = Z;
		19'b0111101000110111111: color_data = Z;
		19'b0111101000111000000: color_data = Z;
		19'b0111101000111000001: color_data = Z;
		19'b0111101000111000010: color_data = Z;
		19'b0111101000111000011: color_data = Z;
		19'b0111101000111000100: color_data = Z;
		19'b0111101000111000101: color_data = Z;
		19'b0111101000111000110: color_data = Z;
		19'b0111101000111000111: color_data = Z;
		19'b0111101000111001000: color_data = Z;
		19'b0111101010010101111: color_data = Z;
		19'b0111101010010110000: color_data = Z;
		19'b0111101010010110001: color_data = Z;
		19'b0111101010010110010: color_data = Z;
		19'b0111101010010110011: color_data = Z;
		19'b0111101010010110100: color_data = Z;
		19'b0111101010010110101: color_data = Z;
		19'b0111101010010110110: color_data = Z;
		19'b0111101010010110111: color_data = Z;
		19'b0111101010010111000: color_data = Z;
		19'b0111101010010111001: color_data = Z;
		19'b0111101010010111010: color_data = Z;
		19'b0111101010010111011: color_data = Z;
		19'b0111101010010111100: color_data = Z;
		19'b0111101010010111101: color_data = Z;
		19'b0111101010010111110: color_data = Z;
		19'b0111101010010111111: color_data = Z;
		19'b0111101010011001010: color_data = Z;
		19'b0111101010011001011: color_data = Z;
		19'b0111101010011001100: color_data = Z;
		19'b0111101010011001101: color_data = Z;
		19'b0111101010011001110: color_data = Z;
		19'b0111101010011001111: color_data = Z;
		19'b0111101010011010000: color_data = Z;
		19'b0111101010011010001: color_data = Z;
		19'b0111101010011010010: color_data = Z;
		19'b0111101010011010011: color_data = Z;
		19'b0111101010011010100: color_data = Z;
		19'b0111101010011010101: color_data = Z;
		19'b0111101010011010110: color_data = Z;
		19'b0111101010011010111: color_data = Z;
		19'b0111101010011011000: color_data = Z;
		19'b0111101010011011001: color_data = Z;
		19'b0111101010011011010: color_data = Z;
		19'b0111101010011011011: color_data = Z;
		19'b0111101010011011100: color_data = Z;
		19'b0111101010011011101: color_data = Z;
		19'b0111101010011011110: color_data = Z;
		19'b0111101010011101110: color_data = Z;
		19'b0111101010011101111: color_data = Z;
		19'b0111101010011110000: color_data = Z;
		19'b0111101010011110001: color_data = Z;
		19'b0111101010011110010: color_data = Z;
		19'b0111101010011110011: color_data = Z;
		19'b0111101010011110100: color_data = Z;
		19'b0111101010011110101: color_data = Z;
		19'b0111101010011110110: color_data = Z;
		19'b0111101010011110111: color_data = Z;
		19'b0111101010011111000: color_data = Z;
		19'b0111101010011111001: color_data = Z;
		19'b0111101010011111010: color_data = Z;
		19'b0111101010011111011: color_data = Z;
		19'b0111101010011111100: color_data = Z;
		19'b0111101010011111101: color_data = Z;
		19'b0111101010011111110: color_data = Z;
		19'b0111101010011111111: color_data = Z;
		19'b0111101010100000000: color_data = Z;
		19'b0111101010100000001: color_data = Z;
		19'b0111101010100000010: color_data = Z;
		19'b0111101010100000011: color_data = Z;
		19'b0111101010100000100: color_data = Z;
		19'b0111101010100001101: color_data = Z;
		19'b0111101010100001110: color_data = Z;
		19'b0111101010100001111: color_data = Z;
		19'b0111101010100010000: color_data = Z;
		19'b0111101010100010001: color_data = Z;
		19'b0111101010100010010: color_data = Z;
		19'b0111101010100010011: color_data = Z;
		19'b0111101010100010100: color_data = Z;
		19'b0111101010100010101: color_data = Z;
		19'b0111101010100010110: color_data = Z;
		19'b0111101010100010111: color_data = Z;
		19'b0111101010100011000: color_data = Z;
		19'b0111101010100011001: color_data = Z;
		19'b0111101010100011010: color_data = Z;
		19'b0111101010100011011: color_data = Z;
		19'b0111101010100011100: color_data = Z;
		19'b0111101010100011101: color_data = Z;
		19'b0111101010100011110: color_data = Z;
		19'b0111101010100011111: color_data = Z;
		19'b0111101010100100000: color_data = Z;
		19'b0111101010100100001: color_data = Z;
		19'b0111101010100100010: color_data = Z;
		19'b0111101010100100011: color_data = Z;
		19'b0111101010100100100: color_data = Z;
		19'b0111101010100100101: color_data = Z;
		19'b0111101010100100110: color_data = Z;
		19'b0111101010100100111: color_data = Z;
		19'b0111101010100101000: color_data = Z;
		19'b0111101010100101001: color_data = Z;
		19'b0111101010100101010: color_data = Z;
		19'b0111101010100101011: color_data = Z;
		19'b0111101010100101100: color_data = Z;
		19'b0111101010100101101: color_data = Z;
		19'b0111101010100101110: color_data = Z;
		19'b0111101010100101111: color_data = Z;
		19'b0111101010100110000: color_data = Z;
		19'b0111101010100110001: color_data = Z;
		19'b0111101010100110110: color_data = Z;
		19'b0111101010100110111: color_data = Z;
		19'b0111101010100111000: color_data = Z;
		19'b0111101010100111001: color_data = Z;
		19'b0111101010100111010: color_data = Z;
		19'b0111101010100111011: color_data = Z;
		19'b0111101010100111100: color_data = Z;
		19'b0111101010100111101: color_data = Z;
		19'b0111101010100111110: color_data = Z;
		19'b0111101010100111111: color_data = Z;
		19'b0111101010101000000: color_data = Z;
		19'b0111101010101000001: color_data = Z;
		19'b0111101010101000010: color_data = Z;
		19'b0111101010101000011: color_data = Z;
		19'b0111101010101000100: color_data = Z;
		19'b0111101010101000101: color_data = Z;
		19'b0111101010101000110: color_data = Z;
		19'b0111101010101000111: color_data = Z;
		19'b0111101010101001000: color_data = Z;
		19'b0111101010101001001: color_data = Z;
		19'b0111101010101001010: color_data = Z;
		19'b0111101010101001011: color_data = Z;
		19'b0111101010101001100: color_data = Z;
		19'b0111101010101001101: color_data = Z;
		19'b0111101010101001110: color_data = Z;
		19'b0111101010101001111: color_data = Z;
		19'b0111101010101010000: color_data = Z;
		19'b0111101010101010001: color_data = Z;
		19'b0111101010101010010: color_data = Z;
		19'b0111101010101010011: color_data = Z;
		19'b0111101010101010100: color_data = Z;
		19'b0111101010101010101: color_data = Z;
		19'b0111101010101010110: color_data = Z;
		19'b0111101010101010111: color_data = Z;
		19'b0111101010101011000: color_data = Z;
		19'b0111101010101011001: color_data = Z;
		19'b0111101010101011010: color_data = Z;
		19'b0111101010101011011: color_data = Z;
		19'b0111101010101011100: color_data = Z;
		19'b0111101010101011101: color_data = Z;
		19'b0111101010101011110: color_data = Z;
		19'b0111101010101011111: color_data = Z;
		19'b0111101010101100000: color_data = Z;
		19'b0111101010101100001: color_data = Z;
		19'b0111101010101100010: color_data = Z;
		19'b0111101010101100011: color_data = Z;
		19'b0111101010101100100: color_data = Z;
		19'b0111101010101100110: color_data = Z;
		19'b0111101010101100111: color_data = Z;
		19'b0111101010101101000: color_data = Z;
		19'b0111101010101101001: color_data = Z;
		19'b0111101010101101010: color_data = Z;
		19'b0111101010101101011: color_data = Z;
		19'b0111101010101101100: color_data = Z;
		19'b0111101010101101101: color_data = Z;
		19'b0111101010101101110: color_data = Z;
		19'b0111101010101101111: color_data = Z;
		19'b0111101010101110000: color_data = Z;
		19'b0111101010101110001: color_data = Z;
		19'b0111101010101110010: color_data = Z;
		19'b0111101010101110011: color_data = Z;
		19'b0111101010101110100: color_data = Z;
		19'b0111101010101110101: color_data = Z;
		19'b0111101010101110110: color_data = Z;
		19'b0111101010101110111: color_data = Z;
		19'b0111101010101111000: color_data = Z;
		19'b0111101010101111001: color_data = Z;
		19'b0111101010101111010: color_data = Z;
		19'b0111101010101111011: color_data = Z;
		19'b0111101010101111100: color_data = Z;
		19'b0111101010101111101: color_data = Z;
		19'b0111101010101111110: color_data = Z;
		19'b0111101010101111111: color_data = Z;
		19'b0111101010110000000: color_data = Z;
		19'b0111101010110000001: color_data = Z;
		19'b0111101010110000010: color_data = Z;
		19'b0111101010110000011: color_data = Z;
		19'b0111101010110000100: color_data = Z;
		19'b0111101010110000101: color_data = Z;
		19'b0111101010110000110: color_data = Z;
		19'b0111101010110000111: color_data = Z;
		19'b0111101010110001000: color_data = Z;
		19'b0111101010110001001: color_data = Z;
		19'b0111101010110001110: color_data = Z;
		19'b0111101010110001111: color_data = Z;
		19'b0111101010110010000: color_data = Z;
		19'b0111101010110010001: color_data = Z;
		19'b0111101010110010010: color_data = Z;
		19'b0111101010110010011: color_data = Z;
		19'b0111101010110011001: color_data = Z;
		19'b0111101010110011010: color_data = Z;
		19'b0111101010110011011: color_data = Z;
		19'b0111101010110011100: color_data = Z;
		19'b0111101010110011101: color_data = Z;
		19'b0111101010110011110: color_data = Z;
		19'b0111101010110101000: color_data = Z;
		19'b0111101010110101001: color_data = Z;
		19'b0111101010110101010: color_data = Z;
		19'b0111101010110101011: color_data = Z;
		19'b0111101010110101100: color_data = Z;
		19'b0111101010110101101: color_data = Z;
		19'b0111101010110101110: color_data = Z;
		19'b0111101010110101111: color_data = Z;
		19'b0111101010110110000: color_data = Z;
		19'b0111101010110110001: color_data = Z;
		19'b0111101010110110010: color_data = Z;
		19'b0111101010110110011: color_data = Z;
		19'b0111101010110110100: color_data = Z;
		19'b0111101010110110101: color_data = Z;
		19'b0111101010110110110: color_data = Z;
		19'b0111101010110110111: color_data = Z;
		19'b0111101010110111010: color_data = Z;
		19'b0111101010110111011: color_data = Z;
		19'b0111101010110111100: color_data = Z;
		19'b0111101010110111101: color_data = Z;
		19'b0111101010110111110: color_data = Z;
		19'b0111101010110111111: color_data = Z;
		19'b0111101010111000000: color_data = Z;
		19'b0111101010111000001: color_data = Z;
		19'b0111101010111000010: color_data = Z;
		19'b0111101010111000011: color_data = Z;
		19'b0111101010111000100: color_data = Z;
		19'b0111101010111000101: color_data = Z;
		19'b0111101010111000110: color_data = Z;
		19'b0111101010111000111: color_data = Z;
		19'b0111101100010110000: color_data = Z;
		19'b0111101100010110001: color_data = Z;
		19'b0111101100010110010: color_data = Z;
		19'b0111101100010110011: color_data = Z;
		19'b0111101100010110100: color_data = Z;
		19'b0111101100010110101: color_data = Z;
		19'b0111101100010110110: color_data = Z;
		19'b0111101100010110111: color_data = Z;
		19'b0111101100010111000: color_data = Z;
		19'b0111101100010111001: color_data = Z;
		19'b0111101100010111010: color_data = Z;
		19'b0111101100010111011: color_data = Z;
		19'b0111101100010111100: color_data = Z;
		19'b0111101100010111101: color_data = Z;
		19'b0111101100010111110: color_data = Z;
		19'b0111101100010111111: color_data = Z;
		19'b0111101100011001010: color_data = Z;
		19'b0111101100011001011: color_data = Z;
		19'b0111101100011001100: color_data = Z;
		19'b0111101100011001101: color_data = Z;
		19'b0111101100011001110: color_data = Z;
		19'b0111101100011001111: color_data = Z;
		19'b0111101100011010000: color_data = Z;
		19'b0111101100011010001: color_data = Z;
		19'b0111101100011010010: color_data = Z;
		19'b0111101100011010011: color_data = Z;
		19'b0111101100011010100: color_data = Z;
		19'b0111101100011010101: color_data = Z;
		19'b0111101100011010110: color_data = Z;
		19'b0111101100011010111: color_data = Z;
		19'b0111101100011011000: color_data = Z;
		19'b0111101100011011001: color_data = Z;
		19'b0111101100011011010: color_data = Z;
		19'b0111101100011011011: color_data = Z;
		19'b0111101100011011100: color_data = Z;
		19'b0111101100011011101: color_data = Z;
		19'b0111101100011011110: color_data = Z;
		19'b0111101100011011111: color_data = Z;
		19'b0111101100011100000: color_data = Z;
		19'b0111101100011100001: color_data = Z;
		19'b0111101100011100010: color_data = Z;
		19'b0111101100011100011: color_data = Z;
		19'b0111101100011100100: color_data = Z;
		19'b0111101100011100101: color_data = Z;
		19'b0111101100011100110: color_data = Z;
		19'b0111101100011100111: color_data = Z;
		19'b0111101100011101000: color_data = Z;
		19'b0111101100011101001: color_data = Z;
		19'b0111101100011101010: color_data = Z;
		19'b0111101100011101011: color_data = Z;
		19'b0111101100011101100: color_data = Z;
		19'b0111101100011101101: color_data = Z;
		19'b0111101100011101110: color_data = Z;
		19'b0111101100011101111: color_data = Z;
		19'b0111101100011110000: color_data = Z;
		19'b0111101100011110001: color_data = Z;
		19'b0111101100011110010: color_data = Z;
		19'b0111101100011110011: color_data = Z;
		19'b0111101100011110100: color_data = Z;
		19'b0111101100011110101: color_data = Z;
		19'b0111101100011110110: color_data = Z;
		19'b0111101100011110111: color_data = Z;
		19'b0111101100011111000: color_data = Z;
		19'b0111101100011111110: color_data = Z;
		19'b0111101100011111111: color_data = Z;
		19'b0111101100100000000: color_data = Z;
		19'b0111101100100000001: color_data = Z;
		19'b0111101100100000010: color_data = Z;
		19'b0111101100100000011: color_data = Z;
		19'b0111101100100001100: color_data = Z;
		19'b0111101100100001101: color_data = Z;
		19'b0111101100100001110: color_data = Z;
		19'b0111101100100001111: color_data = Z;
		19'b0111101100100010000: color_data = Z;
		19'b0111101100100010001: color_data = Z;
		19'b0111101100100010010: color_data = Z;
		19'b0111101100100010011: color_data = Z;
		19'b0111101100100010100: color_data = Z;
		19'b0111101100100010101: color_data = Z;
		19'b0111101100100010110: color_data = Z;
		19'b0111101100100010111: color_data = Z;
		19'b0111101100100011000: color_data = Z;
		19'b0111101100100011001: color_data = Z;
		19'b0111101100100011010: color_data = Z;
		19'b0111101100100011011: color_data = Z;
		19'b0111101100100011100: color_data = Z;
		19'b0111101100100011101: color_data = Z;
		19'b0111101100100011110: color_data = Z;
		19'b0111101100100011111: color_data = Z;
		19'b0111101100100100000: color_data = Z;
		19'b0111101100100100001: color_data = Z;
		19'b0111101100100100010: color_data = Z;
		19'b0111101100100100011: color_data = Z;
		19'b0111101100100100100: color_data = Z;
		19'b0111101100100100101: color_data = Z;
		19'b0111101100100100110: color_data = Z;
		19'b0111101100100100111: color_data = Z;
		19'b0111101100100101000: color_data = Z;
		19'b0111101100100101001: color_data = Z;
		19'b0111101100100101010: color_data = Z;
		19'b0111101100100101011: color_data = Z;
		19'b0111101100100101100: color_data = Z;
		19'b0111101100100101101: color_data = Z;
		19'b0111101100100101110: color_data = Z;
		19'b0111101100100101111: color_data = Z;
		19'b0111101100100110000: color_data = Z;
		19'b0111101100100110101: color_data = Z;
		19'b0111101100100110110: color_data = Z;
		19'b0111101100100110111: color_data = Z;
		19'b0111101100100111000: color_data = Z;
		19'b0111101100100111001: color_data = Z;
		19'b0111101100100111010: color_data = Z;
		19'b0111101100100111011: color_data = Z;
		19'b0111101100100111100: color_data = Z;
		19'b0111101100100111101: color_data = Z;
		19'b0111101100100111110: color_data = Z;
		19'b0111101100100111111: color_data = Z;
		19'b0111101100101000000: color_data = Z;
		19'b0111101100101000001: color_data = Z;
		19'b0111101100101000010: color_data = Z;
		19'b0111101100101000011: color_data = Z;
		19'b0111101100101000100: color_data = Z;
		19'b0111101100101000101: color_data = Z;
		19'b0111101100101000110: color_data = Z;
		19'b0111101100101000111: color_data = Z;
		19'b0111101100101001000: color_data = Z;
		19'b0111101100101001001: color_data = Z;
		19'b0111101100101001010: color_data = Z;
		19'b0111101100101001011: color_data = Z;
		19'b0111101100101001100: color_data = Z;
		19'b0111101100101001101: color_data = Z;
		19'b0111101100101001110: color_data = Z;
		19'b0111101100101001111: color_data = Z;
		19'b0111101100101010000: color_data = Z;
		19'b0111101100101010001: color_data = Z;
		19'b0111101100101010010: color_data = Z;
		19'b0111101100101010011: color_data = Z;
		19'b0111101100101010100: color_data = Z;
		19'b0111101100101010101: color_data = Z;
		19'b0111101100101010110: color_data = Z;
		19'b0111101100101010111: color_data = Z;
		19'b0111101100101011000: color_data = Z;
		19'b0111101100101011001: color_data = Z;
		19'b0111101100101011010: color_data = Z;
		19'b0111101100101011011: color_data = Z;
		19'b0111101100101011100: color_data = Z;
		19'b0111101100101011101: color_data = Z;
		19'b0111101100101011110: color_data = Z;
		19'b0111101100101011111: color_data = Z;
		19'b0111101100101100000: color_data = Z;
		19'b0111101100101100001: color_data = Z;
		19'b0111101100101100010: color_data = Z;
		19'b0111101100101100011: color_data = Z;
		19'b0111101100101100100: color_data = Z;
		19'b0111101100101100101: color_data = Z;
		19'b0111101100101100110: color_data = Z;
		19'b0111101100101100111: color_data = Z;
		19'b0111101100101101000: color_data = Z;
		19'b0111101100101101001: color_data = Z;
		19'b0111101100101101010: color_data = Z;
		19'b0111101100101101011: color_data = Z;
		19'b0111101100101101100: color_data = Z;
		19'b0111101100101101101: color_data = Z;
		19'b0111101100101101110: color_data = Z;
		19'b0111101100101101111: color_data = Z;
		19'b0111101100101110000: color_data = Z;
		19'b0111101100101110001: color_data = Z;
		19'b0111101100101110010: color_data = Z;
		19'b0111101100101110011: color_data = Z;
		19'b0111101100101110100: color_data = Z;
		19'b0111101100101110101: color_data = Z;
		19'b0111101100101110110: color_data = Z;
		19'b0111101100101110111: color_data = Z;
		19'b0111101100101111000: color_data = Z;
		19'b0111101100101111001: color_data = Z;
		19'b0111101100101111010: color_data = Z;
		19'b0111101100101111011: color_data = Z;
		19'b0111101100101111100: color_data = Z;
		19'b0111101100101111101: color_data = Z;
		19'b0111101100101111110: color_data = Z;
		19'b0111101100101111111: color_data = Z;
		19'b0111101100110000000: color_data = Z;
		19'b0111101100110000001: color_data = Z;
		19'b0111101100110000010: color_data = Z;
		19'b0111101100110000011: color_data = Z;
		19'b0111101100110000100: color_data = Z;
		19'b0111101100110000101: color_data = Z;
		19'b0111101100110000110: color_data = Z;
		19'b0111101100110000111: color_data = Z;
		19'b0111101100110001110: color_data = Z;
		19'b0111101100110001111: color_data = Z;
		19'b0111101100110010000: color_data = Z;
		19'b0111101100110010001: color_data = Z;
		19'b0111101100110010010: color_data = Z;
		19'b0111101100110010011: color_data = Z;
		19'b0111101100110010100: color_data = Z;
		19'b0111101100110011001: color_data = Z;
		19'b0111101100110011010: color_data = Z;
		19'b0111101100110011011: color_data = Z;
		19'b0111101100110011100: color_data = Z;
		19'b0111101100110011101: color_data = Z;
		19'b0111101100110011110: color_data = Z;
		19'b0111101100110011111: color_data = Z;
		19'b0111101100110100000: color_data = Z;
		19'b0111101100110100001: color_data = Z;
		19'b0111101100110100010: color_data = Z;
		19'b0111101100110100011: color_data = Z;
		19'b0111101100110100100: color_data = Z;
		19'b0111101100110100110: color_data = Z;
		19'b0111101100110100111: color_data = Z;
		19'b0111101100110101000: color_data = Z;
		19'b0111101100110101001: color_data = Z;
		19'b0111101100110101010: color_data = Z;
		19'b0111101100110101011: color_data = Z;
		19'b0111101100110101100: color_data = Z;
		19'b0111101100110101101: color_data = Z;
		19'b0111101100110101110: color_data = Z;
		19'b0111101100110101111: color_data = Z;
		19'b0111101100110110000: color_data = Z;
		19'b0111101100110110001: color_data = Z;
		19'b0111101100110110010: color_data = Z;
		19'b0111101100110110011: color_data = Z;
		19'b0111101100110110100: color_data = Z;
		19'b0111101100110110101: color_data = Z;
		19'b0111101100110111001: color_data = Z;
		19'b0111101100110111010: color_data = Z;
		19'b0111101100110111011: color_data = Z;
		19'b0111101100110111100: color_data = Z;
		19'b0111101100110111101: color_data = Z;
		19'b0111101100110111110: color_data = Z;
		19'b0111101100110111111: color_data = Z;
		19'b0111101100111000000: color_data = Z;
		19'b0111101100111000001: color_data = Z;
		19'b0111101100111000010: color_data = Z;
		19'b0111101100111000011: color_data = Z;
		19'b0111101100111000100: color_data = Z;
		19'b0111101100111000101: color_data = Z;
		19'b0111101100111000110: color_data = Z;
		19'b0111101100111000111: color_data = Z;
		19'b0111101110010110000: color_data = Z;
		19'b0111101110010110001: color_data = Z;
		19'b0111101110010110010: color_data = Z;
		19'b0111101110010110011: color_data = Z;
		19'b0111101110010110100: color_data = Z;
		19'b0111101110010110101: color_data = Z;
		19'b0111101110010110110: color_data = Z;
		19'b0111101110010110111: color_data = Z;
		19'b0111101110010111000: color_data = Z;
		19'b0111101110010111001: color_data = Z;
		19'b0111101110010111010: color_data = Z;
		19'b0111101110010111011: color_data = Z;
		19'b0111101110010111100: color_data = Z;
		19'b0111101110010111101: color_data = Z;
		19'b0111101110010111110: color_data = Z;
		19'b0111101110010111111: color_data = Z;
		19'b0111101110011000000: color_data = Z;
		19'b0111101110011001011: color_data = Z;
		19'b0111101110011001100: color_data = Z;
		19'b0111101110011001101: color_data = Z;
		19'b0111101110011001110: color_data = Z;
		19'b0111101110011001111: color_data = Z;
		19'b0111101110011010010: color_data = Z;
		19'b0111101110011010011: color_data = Z;
		19'b0111101110011010100: color_data = Z;
		19'b0111101110011010101: color_data = Z;
		19'b0111101110011010110: color_data = Z;
		19'b0111101110011010111: color_data = Z;
		19'b0111101110011011000: color_data = Z;
		19'b0111101110011011001: color_data = Z;
		19'b0111101110011011010: color_data = Z;
		19'b0111101110011011011: color_data = Z;
		19'b0111101110011011100: color_data = Z;
		19'b0111101110011011101: color_data = Z;
		19'b0111101110011011110: color_data = Z;
		19'b0111101110011011111: color_data = Z;
		19'b0111101110011100000: color_data = Z;
		19'b0111101110011100001: color_data = Z;
		19'b0111101110011100010: color_data = Z;
		19'b0111101110011100011: color_data = Z;
		19'b0111101110011100100: color_data = Z;
		19'b0111101110011100101: color_data = Z;
		19'b0111101110011100110: color_data = Z;
		19'b0111101110011100111: color_data = Z;
		19'b0111101110011101000: color_data = Z;
		19'b0111101110011101001: color_data = Z;
		19'b0111101110011101010: color_data = Z;
		19'b0111101110011101011: color_data = Z;
		19'b0111101110011101100: color_data = Z;
		19'b0111101110011101101: color_data = Z;
		19'b0111101110011101110: color_data = Z;
		19'b0111101110011101111: color_data = Z;
		19'b0111101110011110000: color_data = Z;
		19'b0111101110011110001: color_data = Z;
		19'b0111101110011110010: color_data = Z;
		19'b0111101110011110011: color_data = Z;
		19'b0111101110011110100: color_data = Z;
		19'b0111101110011110101: color_data = Z;
		19'b0111101110011110110: color_data = Z;
		19'b0111101110011110111: color_data = Z;
		19'b0111101110011111110: color_data = Z;
		19'b0111101110011111111: color_data = Z;
		19'b0111101110100000000: color_data = Z;
		19'b0111101110100000001: color_data = Z;
		19'b0111101110100001100: color_data = Z;
		19'b0111101110100001101: color_data = Z;
		19'b0111101110100001110: color_data = Z;
		19'b0111101110100001111: color_data = Z;
		19'b0111101110100010000: color_data = Z;
		19'b0111101110100010001: color_data = Z;
		19'b0111101110100010010: color_data = Z;
		19'b0111101110100010011: color_data = Z;
		19'b0111101110100010100: color_data = Z;
		19'b0111101110100010101: color_data = Z;
		19'b0111101110100010110: color_data = Z;
		19'b0111101110100010111: color_data = Z;
		19'b0111101110100011000: color_data = Z;
		19'b0111101110100011001: color_data = Z;
		19'b0111101110100011010: color_data = Z;
		19'b0111101110100011011: color_data = Z;
		19'b0111101110100011100: color_data = Z;
		19'b0111101110100011101: color_data = Z;
		19'b0111101110100011110: color_data = Z;
		19'b0111101110100011111: color_data = Z;
		19'b0111101110100100000: color_data = Z;
		19'b0111101110100100001: color_data = Z;
		19'b0111101110100100010: color_data = Z;
		19'b0111101110100100011: color_data = Z;
		19'b0111101110100100100: color_data = Z;
		19'b0111101110100100101: color_data = Z;
		19'b0111101110100100110: color_data = Z;
		19'b0111101110100100111: color_data = Z;
		19'b0111101110100101000: color_data = Z;
		19'b0111101110100101001: color_data = Z;
		19'b0111101110100101010: color_data = Z;
		19'b0111101110100101011: color_data = Z;
		19'b0111101110100101100: color_data = Z;
		19'b0111101110100101101: color_data = Z;
		19'b0111101110100101110: color_data = Z;
		19'b0111101110100101111: color_data = Z;
		19'b0111101110100110000: color_data = Z;
		19'b0111101110100110101: color_data = Z;
		19'b0111101110100110110: color_data = Z;
		19'b0111101110100110111: color_data = Z;
		19'b0111101110100111000: color_data = Z;
		19'b0111101110100111001: color_data = Z;
		19'b0111101110100111010: color_data = Z;
		19'b0111101110100111011: color_data = Z;
		19'b0111101110100111100: color_data = Z;
		19'b0111101110100111101: color_data = Z;
		19'b0111101110100111110: color_data = Z;
		19'b0111101110100111111: color_data = Z;
		19'b0111101110101000000: color_data = Z;
		19'b0111101110101000001: color_data = Z;
		19'b0111101110101000010: color_data = Z;
		19'b0111101110101000011: color_data = Z;
		19'b0111101110101000100: color_data = Z;
		19'b0111101110101000101: color_data = Z;
		19'b0111101110101000110: color_data = Z;
		19'b0111101110101000111: color_data = Z;
		19'b0111101110101001000: color_data = Z;
		19'b0111101110101001001: color_data = Z;
		19'b0111101110101001010: color_data = Z;
		19'b0111101110101001011: color_data = Z;
		19'b0111101110101001100: color_data = Z;
		19'b0111101110101001101: color_data = Z;
		19'b0111101110101001110: color_data = Z;
		19'b0111101110101001111: color_data = Z;
		19'b0111101110101010000: color_data = Z;
		19'b0111101110101010001: color_data = Z;
		19'b0111101110101010010: color_data = Z;
		19'b0111101110101010011: color_data = Z;
		19'b0111101110101010100: color_data = Z;
		19'b0111101110101010101: color_data = Z;
		19'b0111101110101010110: color_data = Z;
		19'b0111101110101010111: color_data = Z;
		19'b0111101110101011000: color_data = Z;
		19'b0111101110101011001: color_data = Z;
		19'b0111101110101011010: color_data = Z;
		19'b0111101110101011011: color_data = Z;
		19'b0111101110101011100: color_data = Z;
		19'b0111101110101011101: color_data = Z;
		19'b0111101110101011110: color_data = Z;
		19'b0111101110101011111: color_data = Z;
		19'b0111101110101100000: color_data = Z;
		19'b0111101110101100001: color_data = Z;
		19'b0111101110101100010: color_data = Z;
		19'b0111101110101100011: color_data = Z;
		19'b0111101110101100100: color_data = Z;
		19'b0111101110101100101: color_data = Z;
		19'b0111101110101101000: color_data = Z;
		19'b0111101110101101001: color_data = Z;
		19'b0111101110101101010: color_data = Z;
		19'b0111101110101101011: color_data = Z;
		19'b0111101110101101100: color_data = Z;
		19'b0111101110101101101: color_data = Z;
		19'b0111101110101101110: color_data = Z;
		19'b0111101110101101111: color_data = Z;
		19'b0111101110101110000: color_data = Z;
		19'b0111101110101110001: color_data = Z;
		19'b0111101110101110010: color_data = Z;
		19'b0111101110101110011: color_data = Z;
		19'b0111101110101110100: color_data = Z;
		19'b0111101110101110101: color_data = Z;
		19'b0111101110101110110: color_data = Z;
		19'b0111101110101110111: color_data = Z;
		19'b0111101110101111000: color_data = Z;
		19'b0111101110101111001: color_data = Z;
		19'b0111101110101111010: color_data = Z;
		19'b0111101110101111011: color_data = Z;
		19'b0111101110101111100: color_data = Z;
		19'b0111101110101111101: color_data = Z;
		19'b0111101110101111110: color_data = Z;
		19'b0111101110101111111: color_data = Z;
		19'b0111101110110000000: color_data = Z;
		19'b0111101110110000001: color_data = Z;
		19'b0111101110110000010: color_data = Z;
		19'b0111101110110000011: color_data = Z;
		19'b0111101110110000100: color_data = Z;
		19'b0111101110110000101: color_data = Z;
		19'b0111101110110000110: color_data = Z;
		19'b0111101110110000111: color_data = Z;
		19'b0111101110110001110: color_data = Z;
		19'b0111101110110010000: color_data = Z;
		19'b0111101110110010001: color_data = Z;
		19'b0111101110110010010: color_data = Z;
		19'b0111101110110010011: color_data = Z;
		19'b0111101110110010100: color_data = Z;
		19'b0111101110110010101: color_data = Z;
		19'b0111101110110010110: color_data = Z;
		19'b0111101110110011000: color_data = Z;
		19'b0111101110110011001: color_data = Z;
		19'b0111101110110011010: color_data = Z;
		19'b0111101110110011011: color_data = Z;
		19'b0111101110110011100: color_data = Z;
		19'b0111101110110011101: color_data = Z;
		19'b0111101110110011110: color_data = Z;
		19'b0111101110110011111: color_data = Z;
		19'b0111101110110100000: color_data = Z;
		19'b0111101110110100001: color_data = Z;
		19'b0111101110110100010: color_data = Z;
		19'b0111101110110100011: color_data = Z;
		19'b0111101110110100100: color_data = Z;
		19'b0111101110110100101: color_data = Z;
		19'b0111101110110100110: color_data = Z;
		19'b0111101110110100111: color_data = Z;
		19'b0111101110110101000: color_data = Z;
		19'b0111101110110101001: color_data = Z;
		19'b0111101110110101010: color_data = Z;
		19'b0111101110110101011: color_data = Z;
		19'b0111101110110101100: color_data = Z;
		19'b0111101110110101101: color_data = Z;
		19'b0111101110110101110: color_data = Z;
		19'b0111101110110101111: color_data = Z;
		19'b0111101110110110000: color_data = Z;
		19'b0111101110110110001: color_data = Z;
		19'b0111101110110110010: color_data = Z;
		19'b0111101110110110011: color_data = Z;
		19'b0111101110110111001: color_data = Z;
		19'b0111101110110111010: color_data = Z;
		19'b0111101110110111011: color_data = Z;
		19'b0111101110110111100: color_data = Z;
		19'b0111101110110111101: color_data = Z;
		19'b0111101110110111110: color_data = Z;
		19'b0111101110110111111: color_data = Z;
		19'b0111101110111000000: color_data = Z;
		19'b0111101110111000001: color_data = Z;
		19'b0111101110111000010: color_data = Z;
		19'b0111101110111000011: color_data = Z;
		19'b0111101110111000100: color_data = Z;
		19'b0111101110111000101: color_data = Z;
		19'b0111101110111000110: color_data = Z;
		19'b0111101110111000111: color_data = Z;
		19'b0111110000010110000: color_data = Z;
		19'b0111110000010110001: color_data = Z;
		19'b0111110000010110010: color_data = Z;
		19'b0111110000010110011: color_data = Z;
		19'b0111110000010110100: color_data = Z;
		19'b0111110000010110101: color_data = Z;
		19'b0111110000010110110: color_data = Z;
		19'b0111110000010110111: color_data = Z;
		19'b0111110000010111000: color_data = Z;
		19'b0111110000010111001: color_data = Z;
		19'b0111110000010111010: color_data = Z;
		19'b0111110000010111011: color_data = Z;
		19'b0111110000010111100: color_data = Z;
		19'b0111110000010111101: color_data = Z;
		19'b0111110000010111110: color_data = Z;
		19'b0111110000010111111: color_data = Z;
		19'b0111110000011000000: color_data = Z;
		19'b0111110000011001100: color_data = Z;
		19'b0111110000011001101: color_data = Z;
		19'b0111110000011001110: color_data = Z;
		19'b0111110000011001111: color_data = Z;
		19'b0111110000011010000: color_data = Z;
		19'b0111110000011010011: color_data = Z;
		19'b0111110000011010100: color_data = Z;
		19'b0111110000011010101: color_data = Z;
		19'b0111110000011010110: color_data = Z;
		19'b0111110000011010111: color_data = Z;
		19'b0111110000011011000: color_data = Z;
		19'b0111110000011011001: color_data = Z;
		19'b0111110000011011010: color_data = Z;
		19'b0111110000011011011: color_data = Z;
		19'b0111110000011011100: color_data = Z;
		19'b0111110000011011101: color_data = Z;
		19'b0111110000011011110: color_data = Z;
		19'b0111110000011011111: color_data = Z;
		19'b0111110000011100000: color_data = Z;
		19'b0111110000011100001: color_data = Z;
		19'b0111110000011100010: color_data = Z;
		19'b0111110000011100011: color_data = Z;
		19'b0111110000011100100: color_data = Z;
		19'b0111110000011100101: color_data = Z;
		19'b0111110000011100110: color_data = Z;
		19'b0111110000011100111: color_data = Z;
		19'b0111110000011101000: color_data = Z;
		19'b0111110000011101001: color_data = Z;
		19'b0111110000011101010: color_data = Z;
		19'b0111110000011101011: color_data = Z;
		19'b0111110000011101100: color_data = Z;
		19'b0111110000011101101: color_data = Z;
		19'b0111110000011101110: color_data = Z;
		19'b0111110000011101111: color_data = Z;
		19'b0111110000011110000: color_data = Z;
		19'b0111110000011110001: color_data = Z;
		19'b0111110000011110010: color_data = Z;
		19'b0111110000011110011: color_data = Z;
		19'b0111110000011110101: color_data = Z;
		19'b0111110000011110110: color_data = Z;
		19'b0111110000011111110: color_data = Z;
		19'b0111110000011111111: color_data = Z;
		19'b0111110000100000000: color_data = Z;
		19'b0111110000100000001: color_data = Z;
		19'b0111110000100000010: color_data = Z;
		19'b0111110000100001100: color_data = Z;
		19'b0111110000100001101: color_data = Z;
		19'b0111110000100001110: color_data = Z;
		19'b0111110000100001111: color_data = Z;
		19'b0111110000100010000: color_data = Z;
		19'b0111110000100010001: color_data = Z;
		19'b0111110000100010010: color_data = Z;
		19'b0111110000100010011: color_data = Z;
		19'b0111110000100010100: color_data = Z;
		19'b0111110000100010101: color_data = Z;
		19'b0111110000100010110: color_data = Z;
		19'b0111110000100010111: color_data = Z;
		19'b0111110000100011000: color_data = Z;
		19'b0111110000100011001: color_data = Z;
		19'b0111110000100011010: color_data = Z;
		19'b0111110000100011011: color_data = Z;
		19'b0111110000100011100: color_data = Z;
		19'b0111110000100011101: color_data = Z;
		19'b0111110000100011110: color_data = Z;
		19'b0111110000100011111: color_data = Z;
		19'b0111110000100100000: color_data = Z;
		19'b0111110000100100001: color_data = Z;
		19'b0111110000100100010: color_data = Z;
		19'b0111110000100100011: color_data = Z;
		19'b0111110000100100100: color_data = Z;
		19'b0111110000100100101: color_data = Z;
		19'b0111110000100100110: color_data = Z;
		19'b0111110000100100111: color_data = Z;
		19'b0111110000100101000: color_data = Z;
		19'b0111110000100101001: color_data = Z;
		19'b0111110000100101010: color_data = Z;
		19'b0111110000100101011: color_data = Z;
		19'b0111110000100101100: color_data = Z;
		19'b0111110000100101101: color_data = Z;
		19'b0111110000100101110: color_data = Z;
		19'b0111110000100101111: color_data = Z;
		19'b0111110000100110100: color_data = Z;
		19'b0111110000100110101: color_data = Z;
		19'b0111110000100110110: color_data = Z;
		19'b0111110000100110111: color_data = Z;
		19'b0111110000100111000: color_data = Z;
		19'b0111110000100111001: color_data = Z;
		19'b0111110000100111010: color_data = Z;
		19'b0111110000100111011: color_data = Z;
		19'b0111110000100111100: color_data = Z;
		19'b0111110000100111101: color_data = Z;
		19'b0111110000100111110: color_data = Z;
		19'b0111110000100111111: color_data = Z;
		19'b0111110000101000010: color_data = Z;
		19'b0111110000101000011: color_data = Z;
		19'b0111110000101000100: color_data = Z;
		19'b0111110000101000101: color_data = Z;
		19'b0111110000101000110: color_data = Z;
		19'b0111110000101000111: color_data = Z;
		19'b0111110000101001000: color_data = Z;
		19'b0111110000101001001: color_data = Z;
		19'b0111110000101001010: color_data = Z;
		19'b0111110000101001011: color_data = Z;
		19'b0111110000101001100: color_data = Z;
		19'b0111110000101001101: color_data = Z;
		19'b0111110000101001110: color_data = Z;
		19'b0111110000101001111: color_data = Z;
		19'b0111110000101010000: color_data = Z;
		19'b0111110000101010001: color_data = Z;
		19'b0111110000101010010: color_data = Z;
		19'b0111110000101010011: color_data = Z;
		19'b0111110000101010100: color_data = Z;
		19'b0111110000101010101: color_data = Z;
		19'b0111110000101010110: color_data = Z;
		19'b0111110000101010111: color_data = Z;
		19'b0111110000101011000: color_data = Z;
		19'b0111110000101011010: color_data = Z;
		19'b0111110000101011011: color_data = Z;
		19'b0111110000101011100: color_data = Z;
		19'b0111110000101011101: color_data = Z;
		19'b0111110000101011110: color_data = Z;
		19'b0111110000101011111: color_data = Z;
		19'b0111110000101100000: color_data = Z;
		19'b0111110000101100001: color_data = Z;
		19'b0111110000101100010: color_data = Z;
		19'b0111110000101100011: color_data = Z;
		19'b0111110000101100100: color_data = Z;
		19'b0111110000101100101: color_data = Z;
		19'b0111110000101100110: color_data = Z;
		19'b0111110000101101000: color_data = Z;
		19'b0111110000101101001: color_data = Z;
		19'b0111110000101101010: color_data = Z;
		19'b0111110000101101011: color_data = Z;
		19'b0111110000101101100: color_data = Z;
		19'b0111110000101101101: color_data = Z;
		19'b0111110000101101110: color_data = Z;
		19'b0111110000101101111: color_data = Z;
		19'b0111110000101110000: color_data = Z;
		19'b0111110000101110001: color_data = Z;
		19'b0111110000101110010: color_data = Z;
		19'b0111110000101110011: color_data = Z;
		19'b0111110000101110100: color_data = Z;
		19'b0111110000101110101: color_data = Z;
		19'b0111110000101110110: color_data = Z;
		19'b0111110000101110111: color_data = Z;
		19'b0111110000101111000: color_data = Z;
		19'b0111110000101111001: color_data = Z;
		19'b0111110000101111010: color_data = Z;
		19'b0111110000101111011: color_data = Z;
		19'b0111110000101111100: color_data = Z;
		19'b0111110000101111101: color_data = Z;
		19'b0111110000101111110: color_data = Z;
		19'b0111110000101111111: color_data = Z;
		19'b0111110000110000000: color_data = Z;
		19'b0111110000110000001: color_data = Z;
		19'b0111110000110000010: color_data = Z;
		19'b0111110000110000011: color_data = Z;
		19'b0111110000110000100: color_data = Z;
		19'b0111110000110000101: color_data = Z;
		19'b0111110000110000110: color_data = Z;
		19'b0111110000110000111: color_data = Z;
		19'b0111110000110010001: color_data = Z;
		19'b0111110000110010010: color_data = Z;
		19'b0111110000110010011: color_data = Z;
		19'b0111110000110010100: color_data = Z;
		19'b0111110000110010101: color_data = Z;
		19'b0111110000110010110: color_data = Z;
		19'b0111110000110010111: color_data = Z;
		19'b0111110000110011000: color_data = Z;
		19'b0111110000110011001: color_data = Z;
		19'b0111110000110011010: color_data = Z;
		19'b0111110000110011011: color_data = Z;
		19'b0111110000110011100: color_data = Z;
		19'b0111110000110011101: color_data = Z;
		19'b0111110000110011110: color_data = Z;
		19'b0111110000110011111: color_data = Z;
		19'b0111110000110100000: color_data = Z;
		19'b0111110000110100001: color_data = Z;
		19'b0111110000110100010: color_data = Z;
		19'b0111110000110100011: color_data = Z;
		19'b0111110000110100100: color_data = Z;
		19'b0111110000110100101: color_data = Z;
		19'b0111110000110100110: color_data = Z;
		19'b0111110000110100111: color_data = Z;
		19'b0111110000110101000: color_data = Z;
		19'b0111110000110101001: color_data = Z;
		19'b0111110000110101010: color_data = Z;
		19'b0111110000110101011: color_data = Z;
		19'b0111110000110101100: color_data = Z;
		19'b0111110000110101101: color_data = Z;
		19'b0111110000110101110: color_data = Z;
		19'b0111110000110101111: color_data = Z;
		19'b0111110000110110000: color_data = Z;
		19'b0111110000110110001: color_data = Z;
		19'b0111110000110111000: color_data = Z;
		19'b0111110000110111001: color_data = Z;
		19'b0111110000110111010: color_data = Z;
		19'b0111110000110111011: color_data = Z;
		19'b0111110000110111100: color_data = Z;
		19'b0111110000111000000: color_data = Z;
		19'b0111110000111000001: color_data = Z;
		19'b0111110000111000010: color_data = Z;
		19'b0111110000111000011: color_data = Z;
		19'b0111110000111000100: color_data = Z;
		19'b0111110000111000101: color_data = Z;
		19'b0111110000111000110: color_data = Z;
		19'b0111110000111000111: color_data = Z;
		19'b0111110000111001000: color_data = Z;
		19'b0111110010010110001: color_data = Z;
		19'b0111110010010110010: color_data = Z;
		19'b0111110010010110011: color_data = Z;
		19'b0111110010010110100: color_data = Z;
		19'b0111110010010110101: color_data = Z;
		19'b0111110010010110110: color_data = Z;
		19'b0111110010010110111: color_data = Z;
		19'b0111110010010111000: color_data = Z;
		19'b0111110010010111001: color_data = Z;
		19'b0111110010010111010: color_data = Z;
		19'b0111110010010111011: color_data = Z;
		19'b0111110010010111100: color_data = Z;
		19'b0111110010010111101: color_data = Z;
		19'b0111110010010111110: color_data = Z;
		19'b0111110010010111111: color_data = Z;
		19'b0111110010011000000: color_data = Z;
		19'b0111110010011000001: color_data = Z;
		19'b0111110010011001101: color_data = Z;
		19'b0111110010011001110: color_data = Z;
		19'b0111110010011001111: color_data = Z;
		19'b0111110010011010000: color_data = Z;
		19'b0111110010011010100: color_data = Z;
		19'b0111110010011010101: color_data = Z;
		19'b0111110010011010110: color_data = Z;
		19'b0111110010011010111: color_data = Z;
		19'b0111110010011011000: color_data = Z;
		19'b0111110010011011001: color_data = Z;
		19'b0111110010011011010: color_data = Z;
		19'b0111110010011011011: color_data = Z;
		19'b0111110010011011100: color_data = Z;
		19'b0111110010011011101: color_data = Z;
		19'b0111110010011011110: color_data = Z;
		19'b0111110010011011111: color_data = Z;
		19'b0111110010011100000: color_data = Z;
		19'b0111110010011100001: color_data = Z;
		19'b0111110010011100010: color_data = Z;
		19'b0111110010011100011: color_data = Z;
		19'b0111110010011100100: color_data = Z;
		19'b0111110010011100101: color_data = Z;
		19'b0111110010011100110: color_data = Z;
		19'b0111110010011100111: color_data = Z;
		19'b0111110010011101000: color_data = Z;
		19'b0111110010011101001: color_data = Z;
		19'b0111110010011101010: color_data = Z;
		19'b0111110010011101011: color_data = Z;
		19'b0111110010011101100: color_data = Z;
		19'b0111110010011101101: color_data = Z;
		19'b0111110010011101110: color_data = Z;
		19'b0111110010011110100: color_data = Z;
		19'b0111110010011110101: color_data = Z;
		19'b0111110010011110110: color_data = Z;
		19'b0111110010011110111: color_data = Z;
		19'b0111110010011111000: color_data = Z;
		19'b0111110010011111001: color_data = Z;
		19'b0111110010011111101: color_data = Z;
		19'b0111110010011111110: color_data = Z;
		19'b0111110010011111111: color_data = Z;
		19'b0111110010100000000: color_data = Z;
		19'b0111110010100000001: color_data = Z;
		19'b0111110010100001101: color_data = Z;
		19'b0111110010100001110: color_data = Z;
		19'b0111110010100001111: color_data = Z;
		19'b0111110010100010000: color_data = Z;
		19'b0111110010100010001: color_data = Z;
		19'b0111110010100010010: color_data = Z;
		19'b0111110010100010011: color_data = Z;
		19'b0111110010100010100: color_data = Z;
		19'b0111110010100010101: color_data = Z;
		19'b0111110010100010110: color_data = Z;
		19'b0111110010100010111: color_data = Z;
		19'b0111110010100011000: color_data = Z;
		19'b0111110010100011001: color_data = Z;
		19'b0111110010100011010: color_data = Z;
		19'b0111110010100011011: color_data = Z;
		19'b0111110010100011100: color_data = Z;
		19'b0111110010100011101: color_data = Z;
		19'b0111110010100011110: color_data = Z;
		19'b0111110010100011111: color_data = Z;
		19'b0111110010100100000: color_data = Z;
		19'b0111110010100100001: color_data = Z;
		19'b0111110010100100010: color_data = Z;
		19'b0111110010100100011: color_data = Z;
		19'b0111110010100100100: color_data = Z;
		19'b0111110010100100101: color_data = Z;
		19'b0111110010100100110: color_data = Z;
		19'b0111110010100100111: color_data = Z;
		19'b0111110010100101000: color_data = Z;
		19'b0111110010100101001: color_data = Z;
		19'b0111110010100101010: color_data = Z;
		19'b0111110010100101011: color_data = Z;
		19'b0111110010100101100: color_data = Z;
		19'b0111110010100101101: color_data = Z;
		19'b0111110010100101110: color_data = Z;
		19'b0111110010100101111: color_data = Z;
		19'b0111110010100110100: color_data = Z;
		19'b0111110010100110110: color_data = Z;
		19'b0111110010100110111: color_data = Z;
		19'b0111110010100111000: color_data = Z;
		19'b0111110010100111001: color_data = Z;
		19'b0111110010100111010: color_data = Z;
		19'b0111110010100111011: color_data = Z;
		19'b0111110010100111100: color_data = Z;
		19'b0111110010100111101: color_data = Z;
		19'b0111110010100111110: color_data = Z;
		19'b0111110010100111111: color_data = Z;
		19'b0111110010101000010: color_data = Z;
		19'b0111110010101000011: color_data = Z;
		19'b0111110010101000100: color_data = Z;
		19'b0111110010101000101: color_data = Z;
		19'b0111110010101000110: color_data = Z;
		19'b0111110010101000111: color_data = Z;
		19'b0111110010101001000: color_data = Z;
		19'b0111110010101001001: color_data = Z;
		19'b0111110010101001010: color_data = Z;
		19'b0111110010101001011: color_data = Z;
		19'b0111110010101001100: color_data = Z;
		19'b0111110010101001101: color_data = Z;
		19'b0111110010101001110: color_data = Z;
		19'b0111110010101001111: color_data = Z;
		19'b0111110010101010000: color_data = Z;
		19'b0111110010101010001: color_data = Z;
		19'b0111110010101010010: color_data = Z;
		19'b0111110010101010011: color_data = Z;
		19'b0111110010101010100: color_data = Z;
		19'b0111110010101010101: color_data = Z;
		19'b0111110010101010110: color_data = Z;
		19'b0111110010101010111: color_data = Z;
		19'b0111110010101011000: color_data = Z;
		19'b0111110010101011010: color_data = Z;
		19'b0111110010101011011: color_data = Z;
		19'b0111110010101011100: color_data = Z;
		19'b0111110010101011101: color_data = Z;
		19'b0111110010101011110: color_data = Z;
		19'b0111110010101011111: color_data = Z;
		19'b0111110010101100000: color_data = Z;
		19'b0111110010101100001: color_data = Z;
		19'b0111110010101100010: color_data = Z;
		19'b0111110010101100011: color_data = Z;
		19'b0111110010101100100: color_data = Z;
		19'b0111110010101100101: color_data = Z;
		19'b0111110010101100110: color_data = Z;
		19'b0111110010101101001: color_data = Z;
		19'b0111110010101101010: color_data = Z;
		19'b0111110010101101011: color_data = Z;
		19'b0111110010101101100: color_data = Z;
		19'b0111110010101101101: color_data = Z;
		19'b0111110010101101110: color_data = Z;
		19'b0111110010101101111: color_data = Z;
		19'b0111110010101110000: color_data = Z;
		19'b0111110010101110001: color_data = Z;
		19'b0111110010101110010: color_data = Z;
		19'b0111110010101110011: color_data = Z;
		19'b0111110010101110100: color_data = Z;
		19'b0111110010101110101: color_data = Z;
		19'b0111110010101110110: color_data = Z;
		19'b0111110010101110111: color_data = Z;
		19'b0111110010101111000: color_data = Z;
		19'b0111110010101111001: color_data = Z;
		19'b0111110010101111010: color_data = Z;
		19'b0111110010101111011: color_data = Z;
		19'b0111110010101111100: color_data = Z;
		19'b0111110010101111101: color_data = Z;
		19'b0111110010101111110: color_data = Z;
		19'b0111110010101111111: color_data = Z;
		19'b0111110010110000000: color_data = Z;
		19'b0111110010110000001: color_data = Z;
		19'b0111110010110000010: color_data = Z;
		19'b0111110010110000011: color_data = Z;
		19'b0111110010110000100: color_data = Z;
		19'b0111110010110000101: color_data = Z;
		19'b0111110010110000110: color_data = Z;
		19'b0111110010110000111: color_data = Z;
		19'b0111110010110001000: color_data = Z;
		19'b0111110010110010001: color_data = Z;
		19'b0111110010110010010: color_data = Z;
		19'b0111110010110010011: color_data = Z;
		19'b0111110010110010100: color_data = Z;
		19'b0111110010110010101: color_data = Z;
		19'b0111110010110010110: color_data = Z;
		19'b0111110010110010111: color_data = Z;
		19'b0111110010110011000: color_data = Z;
		19'b0111110010110011001: color_data = Z;
		19'b0111110010110011010: color_data = Z;
		19'b0111110010110011011: color_data = Z;
		19'b0111110010110011100: color_data = Z;
		19'b0111110010110011101: color_data = Z;
		19'b0111110010110011110: color_data = Z;
		19'b0111110010110011111: color_data = Z;
		19'b0111110010110100000: color_data = Z;
		19'b0111110010110100001: color_data = Z;
		19'b0111110010110100010: color_data = Z;
		19'b0111110010110100011: color_data = Z;
		19'b0111110010110100100: color_data = Z;
		19'b0111110010110100101: color_data = Z;
		19'b0111110010110100110: color_data = Z;
		19'b0111110010110100111: color_data = Z;
		19'b0111110010110101000: color_data = Z;
		19'b0111110010110101001: color_data = Z;
		19'b0111110010110101010: color_data = Z;
		19'b0111110010110101011: color_data = Z;
		19'b0111110010110101100: color_data = Z;
		19'b0111110010110101101: color_data = Z;
		19'b0111110010110101110: color_data = Z;
		19'b0111110010110101111: color_data = Z;
		19'b0111110010110110111: color_data = Z;
		19'b0111110010110111000: color_data = Z;
		19'b0111110010110111001: color_data = Z;
		19'b0111110010110111010: color_data = Z;
		19'b0111110010110111011: color_data = Z;
		19'b0111110010110111100: color_data = Z;
		19'b0111110010111000000: color_data = Z;
		19'b0111110010111000001: color_data = Z;
		19'b0111110010111000010: color_data = Z;
		19'b0111110010111000011: color_data = Z;
		19'b0111110010111000100: color_data = Z;
		19'b0111110010111000101: color_data = Z;
		19'b0111110010111000110: color_data = Z;
		19'b0111110010111000111: color_data = Z;
		19'b0111110100010110001: color_data = Z;
		19'b0111110100010110010: color_data = Z;
		19'b0111110100010110011: color_data = Z;
		19'b0111110100010110100: color_data = Z;
		19'b0111110100010110101: color_data = Z;
		19'b0111110100010110110: color_data = Z;
		19'b0111110100010110111: color_data = Z;
		19'b0111110100010111000: color_data = Z;
		19'b0111110100010111001: color_data = Z;
		19'b0111110100010111010: color_data = Z;
		19'b0111110100010111011: color_data = Z;
		19'b0111110100010111100: color_data = Z;
		19'b0111110100010111101: color_data = Z;
		19'b0111110100010111110: color_data = Z;
		19'b0111110100010111111: color_data = Z;
		19'b0111110100011000000: color_data = Z;
		19'b0111110100011000001: color_data = Z;
		19'b0111110100011000010: color_data = Z;
		19'b0111110100011001111: color_data = Z;
		19'b0111110100011010000: color_data = Z;
		19'b0111110100011010100: color_data = Z;
		19'b0111110100011010101: color_data = Z;
		19'b0111110100011010110: color_data = Z;
		19'b0111110100011010111: color_data = Z;
		19'b0111110100011011000: color_data = Z;
		19'b0111110100011011001: color_data = Z;
		19'b0111110100011011010: color_data = Z;
		19'b0111110100011011011: color_data = Z;
		19'b0111110100011011100: color_data = Z;
		19'b0111110100011011101: color_data = Z;
		19'b0111110100011011110: color_data = Z;
		19'b0111110100011011111: color_data = Z;
		19'b0111110100011100000: color_data = Z;
		19'b0111110100011100001: color_data = Z;
		19'b0111110100011100010: color_data = Z;
		19'b0111110100011100011: color_data = Z;
		19'b0111110100011100100: color_data = Z;
		19'b0111110100011100101: color_data = Z;
		19'b0111110100011100110: color_data = Z;
		19'b0111110100011100111: color_data = Z;
		19'b0111110100011101000: color_data = Z;
		19'b0111110100011101001: color_data = Z;
		19'b0111110100011101010: color_data = Z;
		19'b0111110100011101011: color_data = Z;
		19'b0111110100011110010: color_data = Z;
		19'b0111110100011110011: color_data = Z;
		19'b0111110100011110100: color_data = Z;
		19'b0111110100011110101: color_data = Z;
		19'b0111110100011110110: color_data = Z;
		19'b0111110100011110111: color_data = Z;
		19'b0111110100011111000: color_data = Z;
		19'b0111110100011111001: color_data = Z;
		19'b0111110100011111100: color_data = Z;
		19'b0111110100011111101: color_data = Z;
		19'b0111110100011111110: color_data = Z;
		19'b0111110100100001100: color_data = Z;
		19'b0111110100100001101: color_data = Z;
		19'b0111110100100001110: color_data = Z;
		19'b0111110100100001111: color_data = Z;
		19'b0111110100100010000: color_data = Z;
		19'b0111110100100010001: color_data = Z;
		19'b0111110100100010010: color_data = Z;
		19'b0111110100100010011: color_data = Z;
		19'b0111110100100010100: color_data = Z;
		19'b0111110100100010101: color_data = Z;
		19'b0111110100100010110: color_data = Z;
		19'b0111110100100010111: color_data = Z;
		19'b0111110100100011000: color_data = Z;
		19'b0111110100100011001: color_data = Z;
		19'b0111110100100011010: color_data = Z;
		19'b0111110100100011011: color_data = Z;
		19'b0111110100100011100: color_data = Z;
		19'b0111110100100011101: color_data = Z;
		19'b0111110100100011110: color_data = Z;
		19'b0111110100100011111: color_data = Z;
		19'b0111110100100100000: color_data = Z;
		19'b0111110100100100001: color_data = Z;
		19'b0111110100100100010: color_data = Z;
		19'b0111110100100100011: color_data = Z;
		19'b0111110100100100100: color_data = Z;
		19'b0111110100100100101: color_data = Z;
		19'b0111110100100100110: color_data = Z;
		19'b0111110100100100111: color_data = Z;
		19'b0111110100100101000: color_data = Z;
		19'b0111110100100101001: color_data = Z;
		19'b0111110100100101010: color_data = Z;
		19'b0111110100100101011: color_data = Z;
		19'b0111110100100101100: color_data = Z;
		19'b0111110100100101101: color_data = Z;
		19'b0111110100100101110: color_data = Z;
		19'b0111110100100101111: color_data = Z;
		19'b0111110100100110110: color_data = Z;
		19'b0111110100100110111: color_data = Z;
		19'b0111110100100111000: color_data = Z;
		19'b0111110100100111001: color_data = Z;
		19'b0111110100100111010: color_data = Z;
		19'b0111110100100111011: color_data = Z;
		19'b0111110100100111100: color_data = Z;
		19'b0111110100100111101: color_data = Z;
		19'b0111110100100111110: color_data = Z;
		19'b0111110100100111111: color_data = Z;
		19'b0111110100101000010: color_data = Z;
		19'b0111110100101000011: color_data = Z;
		19'b0111110100101000100: color_data = Z;
		19'b0111110100101000101: color_data = Z;
		19'b0111110100101000110: color_data = Z;
		19'b0111110100101000111: color_data = Z;
		19'b0111110100101001000: color_data = Z;
		19'b0111110100101001001: color_data = Z;
		19'b0111110100101001010: color_data = Z;
		19'b0111110100101001011: color_data = Z;
		19'b0111110100101001100: color_data = Z;
		19'b0111110100101001101: color_data = Z;
		19'b0111110100101001110: color_data = Z;
		19'b0111110100101001111: color_data = Z;
		19'b0111110100101010000: color_data = Z;
		19'b0111110100101010001: color_data = Z;
		19'b0111110100101010010: color_data = Z;
		19'b0111110100101010011: color_data = Z;
		19'b0111110100101010100: color_data = Z;
		19'b0111110100101010101: color_data = Z;
		19'b0111110100101010110: color_data = Z;
		19'b0111110100101010111: color_data = Z;
		19'b0111110100101011000: color_data = Z;
		19'b0111110100101011010: color_data = Z;
		19'b0111110100101011011: color_data = Z;
		19'b0111110100101011100: color_data = Z;
		19'b0111110100101011101: color_data = Z;
		19'b0111110100101011110: color_data = Z;
		19'b0111110100101011111: color_data = Z;
		19'b0111110100101100000: color_data = Z;
		19'b0111110100101100001: color_data = Z;
		19'b0111110100101100010: color_data = Z;
		19'b0111110100101100011: color_data = Z;
		19'b0111110100101100100: color_data = Z;
		19'b0111110100101100101: color_data = Z;
		19'b0111110100101100110: color_data = Z;
		19'b0111110100101101010: color_data = Z;
		19'b0111110100101101011: color_data = Z;
		19'b0111110100101101100: color_data = Z;
		19'b0111110100101101101: color_data = Z;
		19'b0111110100101101110: color_data = Z;
		19'b0111110100101101111: color_data = Z;
		19'b0111110100101110000: color_data = Z;
		19'b0111110100101110001: color_data = Z;
		19'b0111110100101110010: color_data = Z;
		19'b0111110100101110011: color_data = Z;
		19'b0111110100101110100: color_data = Z;
		19'b0111110100101110101: color_data = Z;
		19'b0111110100101110110: color_data = Z;
		19'b0111110100101110111: color_data = Z;
		19'b0111110100101111000: color_data = Z;
		19'b0111110100101111001: color_data = Z;
		19'b0111110100101111010: color_data = Z;
		19'b0111110100101111011: color_data = Z;
		19'b0111110100101111100: color_data = Z;
		19'b0111110100101111101: color_data = Z;
		19'b0111110100101111110: color_data = Z;
		19'b0111110100101111111: color_data = Z;
		19'b0111110100110000000: color_data = Z;
		19'b0111110100110000001: color_data = Z;
		19'b0111110100110000010: color_data = Z;
		19'b0111110100110000011: color_data = Z;
		19'b0111110100110000100: color_data = Z;
		19'b0111110100110000101: color_data = Z;
		19'b0111110100110000110: color_data = Z;
		19'b0111110100110000111: color_data = Z;
		19'b0111110100110001000: color_data = Z;
		19'b0111110100110001001: color_data = Z;
		19'b0111110100110001010: color_data = Z;
		19'b0111110100110010010: color_data = Z;
		19'b0111110100110010011: color_data = Z;
		19'b0111110100110010100: color_data = Z;
		19'b0111110100110010101: color_data = Z;
		19'b0111110100110010110: color_data = Z;
		19'b0111110100110010111: color_data = Z;
		19'b0111110100110011000: color_data = Z;
		19'b0111110100110011001: color_data = Z;
		19'b0111110100110011010: color_data = Z;
		19'b0111110100110011011: color_data = Z;
		19'b0111110100110011100: color_data = Z;
		19'b0111110100110011101: color_data = Z;
		19'b0111110100110011110: color_data = Z;
		19'b0111110100110011111: color_data = Z;
		19'b0111110100110100000: color_data = Z;
		19'b0111110100110100001: color_data = Z;
		19'b0111110100110100010: color_data = Z;
		19'b0111110100110100011: color_data = Z;
		19'b0111110100110100100: color_data = Z;
		19'b0111110100110100101: color_data = Z;
		19'b0111110100110100110: color_data = Z;
		19'b0111110100110100111: color_data = Z;
		19'b0111110100110101000: color_data = Z;
		19'b0111110100110101001: color_data = Z;
		19'b0111110100110101010: color_data = Z;
		19'b0111110100110101011: color_data = Z;
		19'b0111110100110101100: color_data = Z;
		19'b0111110100110101101: color_data = Z;
		19'b0111110100110101110: color_data = Z;
		19'b0111110100110110010: color_data = Z;
		19'b0111110100110110100: color_data = Z;
		19'b0111110100110110101: color_data = Z;
		19'b0111110100110110110: color_data = Z;
		19'b0111110100110110111: color_data = Z;
		19'b0111110100110111000: color_data = Z;
		19'b0111110100110111001: color_data = Z;
		19'b0111110100110111010: color_data = Z;
		19'b0111110100110111011: color_data = Z;
		19'b0111110100110111100: color_data = Z;
		19'b0111110100111000000: color_data = Z;
		19'b0111110100111000001: color_data = Z;
		19'b0111110100111000010: color_data = Z;
		19'b0111110100111000011: color_data = Z;
		19'b0111110100111000100: color_data = Z;
		19'b0111110100111000101: color_data = Z;
		19'b0111110100111000110: color_data = Z;
		19'b0111110100111000111: color_data = Z;
		19'b0111110110010110010: color_data = Z;
		19'b0111110110010110011: color_data = Z;
		19'b0111110110010110100: color_data = Z;
		19'b0111110110010110101: color_data = Z;
		19'b0111110110010110110: color_data = Z;
		19'b0111110110010110111: color_data = Z;
		19'b0111110110010111000: color_data = Z;
		19'b0111110110010111001: color_data = Z;
		19'b0111110110010111010: color_data = Z;
		19'b0111110110010111011: color_data = Z;
		19'b0111110110010111100: color_data = Z;
		19'b0111110110010111101: color_data = Z;
		19'b0111110110010111110: color_data = Z;
		19'b0111110110010111111: color_data = Z;
		19'b0111110110011000000: color_data = Z;
		19'b0111110110011000001: color_data = Z;
		19'b0111110110011000010: color_data = Z;
		19'b0111110110011010101: color_data = Z;
		19'b0111110110011010110: color_data = Z;
		19'b0111110110011010111: color_data = Z;
		19'b0111110110011011000: color_data = Z;
		19'b0111110110011011001: color_data = Z;
		19'b0111110110011011010: color_data = Z;
		19'b0111110110011011011: color_data = Z;
		19'b0111110110011011111: color_data = Z;
		19'b0111110110011100000: color_data = Z;
		19'b0111110110011100001: color_data = Z;
		19'b0111110110011100010: color_data = Z;
		19'b0111110110011100011: color_data = Z;
		19'b0111110110011110000: color_data = Z;
		19'b0111110110011110001: color_data = Z;
		19'b0111110110011110010: color_data = Z;
		19'b0111110110011110011: color_data = Z;
		19'b0111110110011110100: color_data = Z;
		19'b0111110110011110101: color_data = Z;
		19'b0111110110011110110: color_data = Z;
		19'b0111110110011110111: color_data = Z;
		19'b0111110110011111000: color_data = Z;
		19'b0111110110011111001: color_data = Z;
		19'b0111110110011111010: color_data = Z;
		19'b0111110110011111011: color_data = Z;
		19'b0111110110011111100: color_data = Z;
		19'b0111110110100001100: color_data = Z;
		19'b0111110110100001101: color_data = Z;
		19'b0111110110100001110: color_data = Z;
		19'b0111110110100001111: color_data = Z;
		19'b0111110110100010000: color_data = Z;
		19'b0111110110100010001: color_data = Z;
		19'b0111110110100010010: color_data = Z;
		19'b0111110110100010011: color_data = Z;
		19'b0111110110100010100: color_data = Z;
		19'b0111110110100010101: color_data = Z;
		19'b0111110110100010110: color_data = Z;
		19'b0111110110100010111: color_data = Z;
		19'b0111110110100011000: color_data = Z;
		19'b0111110110100011001: color_data = Z;
		19'b0111110110100011010: color_data = Z;
		19'b0111110110100011011: color_data = Z;
		19'b0111110110100011100: color_data = Z;
		19'b0111110110100011101: color_data = Z;
		19'b0111110110100011110: color_data = Z;
		19'b0111110110100011111: color_data = Z;
		19'b0111110110100100000: color_data = Z;
		19'b0111110110100100001: color_data = Z;
		19'b0111110110100100010: color_data = Z;
		19'b0111110110100100011: color_data = Z;
		19'b0111110110100100100: color_data = Z;
		19'b0111110110100100101: color_data = Z;
		19'b0111110110100100110: color_data = Z;
		19'b0111110110100100111: color_data = Z;
		19'b0111110110100101000: color_data = Z;
		19'b0111110110100101001: color_data = Z;
		19'b0111110110100101010: color_data = Z;
		19'b0111110110100101011: color_data = Z;
		19'b0111110110100101100: color_data = Z;
		19'b0111110110100101101: color_data = Z;
		19'b0111110110100101110: color_data = Z;
		19'b0111110110100101111: color_data = Z;
		19'b0111110110100110110: color_data = Z;
		19'b0111110110100110111: color_data = Z;
		19'b0111110110100111000: color_data = Z;
		19'b0111110110100111001: color_data = Z;
		19'b0111110110100111010: color_data = Z;
		19'b0111110110100111011: color_data = Z;
		19'b0111110110100111100: color_data = Z;
		19'b0111110110100111101: color_data = Z;
		19'b0111110110100111110: color_data = Z;
		19'b0111110110100111111: color_data = Z;
		19'b0111110110101000010: color_data = Z;
		19'b0111110110101000011: color_data = Z;
		19'b0111110110101000100: color_data = Z;
		19'b0111110110101000101: color_data = Z;
		19'b0111110110101000110: color_data = Z;
		19'b0111110110101000111: color_data = Z;
		19'b0111110110101001000: color_data = Z;
		19'b0111110110101001001: color_data = Z;
		19'b0111110110101001010: color_data = Z;
		19'b0111110110101001011: color_data = Z;
		19'b0111110110101001100: color_data = Z;
		19'b0111110110101001101: color_data = Z;
		19'b0111110110101001110: color_data = Z;
		19'b0111110110101001111: color_data = Z;
		19'b0111110110101010000: color_data = Z;
		19'b0111110110101010001: color_data = Z;
		19'b0111110110101010010: color_data = Z;
		19'b0111110110101010011: color_data = Z;
		19'b0111110110101010100: color_data = Z;
		19'b0111110110101010101: color_data = Z;
		19'b0111110110101010110: color_data = Z;
		19'b0111110110101010111: color_data = Z;
		19'b0111110110101011000: color_data = Z;
		19'b0111110110101011010: color_data = Z;
		19'b0111110110101011011: color_data = Z;
		19'b0111110110101011100: color_data = Z;
		19'b0111110110101011101: color_data = Z;
		19'b0111110110101011110: color_data = Z;
		19'b0111110110101011111: color_data = Z;
		19'b0111110110101100000: color_data = Z;
		19'b0111110110101100001: color_data = Z;
		19'b0111110110101100010: color_data = Z;
		19'b0111110110101100011: color_data = Z;
		19'b0111110110101100100: color_data = Z;
		19'b0111110110101100101: color_data = Z;
		19'b0111110110101100110: color_data = Z;
		19'b0111110110101101010: color_data = Z;
		19'b0111110110101101011: color_data = Z;
		19'b0111110110101101100: color_data = Z;
		19'b0111110110101101101: color_data = Z;
		19'b0111110110101101110: color_data = Z;
		19'b0111110110101101111: color_data = Z;
		19'b0111110110101110000: color_data = Z;
		19'b0111110110101110001: color_data = Z;
		19'b0111110110101110010: color_data = Z;
		19'b0111110110101110011: color_data = Z;
		19'b0111110110101110100: color_data = Z;
		19'b0111110110101110101: color_data = Z;
		19'b0111110110101110110: color_data = Z;
		19'b0111110110101110111: color_data = Z;
		19'b0111110110101111000: color_data = Z;
		19'b0111110110101111001: color_data = Z;
		19'b0111110110101111010: color_data = Z;
		19'b0111110110101111011: color_data = Z;
		19'b0111110110101111100: color_data = Z;
		19'b0111110110101111101: color_data = Z;
		19'b0111110110101111110: color_data = Z;
		19'b0111110110101111111: color_data = Z;
		19'b0111110110110000000: color_data = Z;
		19'b0111110110110000001: color_data = Z;
		19'b0111110110110000010: color_data = Z;
		19'b0111110110110000011: color_data = Z;
		19'b0111110110110000100: color_data = Z;
		19'b0111110110110000101: color_data = Z;
		19'b0111110110110000110: color_data = Z;
		19'b0111110110110000111: color_data = Z;
		19'b0111110110110001000: color_data = Z;
		19'b0111110110110001001: color_data = Z;
		19'b0111110110110001010: color_data = Z;
		19'b0111110110110001011: color_data = Z;
		19'b0111110110110001100: color_data = Z;
		19'b0111110110110001101: color_data = Z;
		19'b0111110110110010010: color_data = Z;
		19'b0111110110110010011: color_data = Z;
		19'b0111110110110010100: color_data = Z;
		19'b0111110110110010101: color_data = Z;
		19'b0111110110110010110: color_data = Z;
		19'b0111110110110010111: color_data = Z;
		19'b0111110110110011000: color_data = Z;
		19'b0111110110110011001: color_data = Z;
		19'b0111110110110011010: color_data = Z;
		19'b0111110110110011011: color_data = Z;
		19'b0111110110110011100: color_data = Z;
		19'b0111110110110011101: color_data = Z;
		19'b0111110110110011110: color_data = Z;
		19'b0111110110110011111: color_data = Z;
		19'b0111110110110100000: color_data = Z;
		19'b0111110110110100001: color_data = Z;
		19'b0111110110110100010: color_data = Z;
		19'b0111110110110100011: color_data = Z;
		19'b0111110110110100100: color_data = Z;
		19'b0111110110110100101: color_data = Z;
		19'b0111110110110100110: color_data = Z;
		19'b0111110110110100111: color_data = Z;
		19'b0111110110110101000: color_data = Z;
		19'b0111110110110101001: color_data = Z;
		19'b0111110110110101010: color_data = Z;
		19'b0111110110110101011: color_data = Z;
		19'b0111110110110101100: color_data = Z;
		19'b0111110110110101101: color_data = Z;
		19'b0111110110110101110: color_data = Z;
		19'b0111110110110101111: color_data = Z;
		19'b0111110110110110000: color_data = Z;
		19'b0111110110110110001: color_data = Z;
		19'b0111110110110110010: color_data = Z;
		19'b0111110110110110011: color_data = Z;
		19'b0111110110110110100: color_data = Z;
		19'b0111110110110110101: color_data = Z;
		19'b0111110110110110110: color_data = Z;
		19'b0111110110110110111: color_data = Z;
		19'b0111110110110111000: color_data = Z;
		19'b0111110110110111001: color_data = Z;
		19'b0111110110110111010: color_data = Z;
		19'b0111110110110111011: color_data = Z;
		19'b0111110110110111100: color_data = Z;
		19'b0111110110111000000: color_data = Z;
		19'b0111110110111000001: color_data = Z;
		19'b0111110110111000010: color_data = Z;
		19'b0111110110111000011: color_data = Z;
		19'b0111110110111000100: color_data = Z;
		19'b0111110110111000101: color_data = Z;
		19'b0111110110111000110: color_data = Z;
		19'b0111110110111000111: color_data = Z;
		19'b0111111000010110010: color_data = Z;
		19'b0111111000010110011: color_data = Z;
		19'b0111111000010110100: color_data = Z;
		19'b0111111000010110101: color_data = Z;
		19'b0111111000010110110: color_data = Z;
		19'b0111111000010110111: color_data = Z;
		19'b0111111000010111000: color_data = Z;
		19'b0111111000010111001: color_data = Z;
		19'b0111111000010111010: color_data = Z;
		19'b0111111000010111011: color_data = Z;
		19'b0111111000010111100: color_data = Z;
		19'b0111111000010111101: color_data = Z;
		19'b0111111000010111110: color_data = Z;
		19'b0111111000010111111: color_data = Z;
		19'b0111111000011000000: color_data = Z;
		19'b0111111000011000001: color_data = Z;
		19'b0111111000011000010: color_data = Z;
		19'b0111111000011000011: color_data = Z;
		19'b0111111000011001010: color_data = Z;
		19'b0111111000011010110: color_data = Z;
		19'b0111111000011010111: color_data = Z;
		19'b0111111000011011000: color_data = Z;
		19'b0111111000011011001: color_data = Z;
		19'b0111111000011011010: color_data = Z;
		19'b0111111000011110000: color_data = Z;
		19'b0111111000011110001: color_data = Z;
		19'b0111111000011110010: color_data = Z;
		19'b0111111000011110011: color_data = Z;
		19'b0111111000011110100: color_data = Z;
		19'b0111111000011110101: color_data = Z;
		19'b0111111000011110110: color_data = Z;
		19'b0111111000011110111: color_data = Z;
		19'b0111111000011111000: color_data = Z;
		19'b0111111000011111001: color_data = Z;
		19'b0111111000011111010: color_data = Z;
		19'b0111111000011111011: color_data = Z;
		19'b0111111000011111100: color_data = Z;
		19'b0111111000100001011: color_data = Z;
		19'b0111111000100001100: color_data = Z;
		19'b0111111000100001101: color_data = Z;
		19'b0111111000100001110: color_data = Z;
		19'b0111111000100001111: color_data = Z;
		19'b0111111000100010000: color_data = Z;
		19'b0111111000100010001: color_data = Z;
		19'b0111111000100010010: color_data = Z;
		19'b0111111000100010011: color_data = Z;
		19'b0111111000100010100: color_data = Z;
		19'b0111111000100010101: color_data = Z;
		19'b0111111000100010110: color_data = Z;
		19'b0111111000100010111: color_data = Z;
		19'b0111111000100011000: color_data = Z;
		19'b0111111000100011001: color_data = Z;
		19'b0111111000100011010: color_data = Z;
		19'b0111111000100011011: color_data = Z;
		19'b0111111000100011100: color_data = Z;
		19'b0111111000100011101: color_data = Z;
		19'b0111111000100011110: color_data = Z;
		19'b0111111000100011111: color_data = Z;
		19'b0111111000100100000: color_data = Z;
		19'b0111111000100100001: color_data = Z;
		19'b0111111000100100010: color_data = Z;
		19'b0111111000100100011: color_data = Z;
		19'b0111111000100100100: color_data = Z;
		19'b0111111000100100101: color_data = Z;
		19'b0111111000100100110: color_data = Z;
		19'b0111111000100100111: color_data = Z;
		19'b0111111000100101000: color_data = Z;
		19'b0111111000100101001: color_data = Z;
		19'b0111111000100101010: color_data = Z;
		19'b0111111000100101011: color_data = Z;
		19'b0111111000100101100: color_data = Z;
		19'b0111111000100101101: color_data = Z;
		19'b0111111000100101110: color_data = Z;
		19'b0111111000100110110: color_data = Z;
		19'b0111111000100110111: color_data = Z;
		19'b0111111000100111000: color_data = Z;
		19'b0111111000100111001: color_data = Z;
		19'b0111111000100111010: color_data = Z;
		19'b0111111000100111011: color_data = Z;
		19'b0111111000100111100: color_data = Z;
		19'b0111111000100111101: color_data = Z;
		19'b0111111000100111110: color_data = Z;
		19'b0111111000100111111: color_data = Z;
		19'b0111111000101000011: color_data = Z;
		19'b0111111000101000100: color_data = Z;
		19'b0111111000101000101: color_data = Z;
		19'b0111111000101000110: color_data = Z;
		19'b0111111000101000111: color_data = Z;
		19'b0111111000101001000: color_data = Z;
		19'b0111111000101001001: color_data = Z;
		19'b0111111000101001010: color_data = Z;
		19'b0111111000101001011: color_data = Z;
		19'b0111111000101001100: color_data = Z;
		19'b0111111000101001101: color_data = Z;
		19'b0111111000101001110: color_data = Z;
		19'b0111111000101001111: color_data = Z;
		19'b0111111000101010000: color_data = Z;
		19'b0111111000101010001: color_data = Z;
		19'b0111111000101010010: color_data = Z;
		19'b0111111000101010011: color_data = Z;
		19'b0111111000101010100: color_data = Z;
		19'b0111111000101010101: color_data = Z;
		19'b0111111000101010110: color_data = Z;
		19'b0111111000101010111: color_data = Z;
		19'b0111111000101011000: color_data = Z;
		19'b0111111000101011011: color_data = Z;
		19'b0111111000101011100: color_data = Z;
		19'b0111111000101011101: color_data = Z;
		19'b0111111000101011110: color_data = Z;
		19'b0111111000101011111: color_data = Z;
		19'b0111111000101100000: color_data = Z;
		19'b0111111000101100001: color_data = Z;
		19'b0111111000101100010: color_data = Z;
		19'b0111111000101100011: color_data = Z;
		19'b0111111000101100100: color_data = Z;
		19'b0111111000101100101: color_data = Z;
		19'b0111111000101101010: color_data = Z;
		19'b0111111000101101011: color_data = Z;
		19'b0111111000101101100: color_data = Z;
		19'b0111111000101101101: color_data = Z;
		19'b0111111000101101110: color_data = Z;
		19'b0111111000101101111: color_data = Z;
		19'b0111111000101110000: color_data = Z;
		19'b0111111000101110001: color_data = Z;
		19'b0111111000101110010: color_data = Z;
		19'b0111111000101110011: color_data = Z;
		19'b0111111000101110100: color_data = Z;
		19'b0111111000101110101: color_data = Z;
		19'b0111111000101110110: color_data = Z;
		19'b0111111000101110111: color_data = Z;
		19'b0111111000101111000: color_data = Z;
		19'b0111111000101111001: color_data = Z;
		19'b0111111000101111010: color_data = Z;
		19'b0111111000101111011: color_data = Z;
		19'b0111111000101111100: color_data = Z;
		19'b0111111000101111101: color_data = Z;
		19'b0111111000101111110: color_data = Z;
		19'b0111111000101111111: color_data = Z;
		19'b0111111000110000000: color_data = Z;
		19'b0111111000110000001: color_data = Z;
		19'b0111111000110000010: color_data = Z;
		19'b0111111000110000011: color_data = Z;
		19'b0111111000110000100: color_data = Z;
		19'b0111111000110000101: color_data = Z;
		19'b0111111000110000110: color_data = Z;
		19'b0111111000110000111: color_data = Z;
		19'b0111111000110001000: color_data = Z;
		19'b0111111000110001001: color_data = Z;
		19'b0111111000110001010: color_data = Z;
		19'b0111111000110001100: color_data = Z;
		19'b0111111000110001101: color_data = Z;
		19'b0111111000110001110: color_data = Z;
		19'b0111111000110001111: color_data = Z;
		19'b0111111000110010000: color_data = Z;
		19'b0111111000110010001: color_data = Z;
		19'b0111111000110010101: color_data = Z;
		19'b0111111000110010110: color_data = Z;
		19'b0111111000110010111: color_data = Z;
		19'b0111111000110011000: color_data = Z;
		19'b0111111000110011001: color_data = Z;
		19'b0111111000110011010: color_data = Z;
		19'b0111111000110011011: color_data = Z;
		19'b0111111000110011100: color_data = Z;
		19'b0111111000110011101: color_data = Z;
		19'b0111111000110011110: color_data = Z;
		19'b0111111000110011111: color_data = Z;
		19'b0111111000110100000: color_data = Z;
		19'b0111111000110100001: color_data = Z;
		19'b0111111000110100010: color_data = Z;
		19'b0111111000110100011: color_data = Z;
		19'b0111111000110100100: color_data = Z;
		19'b0111111000110100101: color_data = Z;
		19'b0111111000110100110: color_data = Z;
		19'b0111111000110100111: color_data = Z;
		19'b0111111000110101000: color_data = Z;
		19'b0111111000110101001: color_data = Z;
		19'b0111111000110101010: color_data = Z;
		19'b0111111000110101011: color_data = Z;
		19'b0111111000110101100: color_data = Z;
		19'b0111111000110101101: color_data = Z;
		19'b0111111000110101110: color_data = Z;
		19'b0111111000110101111: color_data = Z;
		19'b0111111000110110000: color_data = Z;
		19'b0111111000110110001: color_data = Z;
		19'b0111111000110110010: color_data = Z;
		19'b0111111000110110011: color_data = Z;
		19'b0111111000110110100: color_data = Z;
		19'b0111111000110110101: color_data = Z;
		19'b0111111000110110110: color_data = Z;
		19'b0111111000110110111: color_data = Z;
		19'b0111111000110111000: color_data = Z;
		19'b0111111000110111001: color_data = Z;
		19'b0111111000110111010: color_data = Z;
		19'b0111111000110111011: color_data = Z;
		19'b0111111000110111100: color_data = Z;
		19'b0111111000111000000: color_data = Z;
		19'b0111111000111000001: color_data = Z;
		19'b0111111000111000010: color_data = Z;
		19'b0111111000111000011: color_data = Z;
		19'b0111111000111000100: color_data = Z;
		19'b0111111000111000101: color_data = Z;
		19'b0111111000111000110: color_data = Z;
		19'b0111111000111000111: color_data = Z;
		19'b0111111000111001000: color_data = Z;
		19'b0111111010010110011: color_data = Z;
		19'b0111111010010110100: color_data = Z;
		19'b0111111010010110101: color_data = Z;
		19'b0111111010010110110: color_data = Z;
		19'b0111111010010110111: color_data = Z;
		19'b0111111010010111000: color_data = Z;
		19'b0111111010010111001: color_data = Z;
		19'b0111111010010111010: color_data = Z;
		19'b0111111010010111011: color_data = Z;
		19'b0111111010010111100: color_data = Z;
		19'b0111111010010111101: color_data = Z;
		19'b0111111010010111110: color_data = Z;
		19'b0111111010010111111: color_data = Z;
		19'b0111111010011000000: color_data = Z;
		19'b0111111010011000001: color_data = Z;
		19'b0111111010011000010: color_data = Z;
		19'b0111111010011000011: color_data = Z;
		19'b0111111010011000100: color_data = Z;
		19'b0111111010011001100: color_data = Z;
		19'b0111111010011010110: color_data = Z;
		19'b0111111010011010111: color_data = Z;
		19'b0111111010011011000: color_data = Z;
		19'b0111111010011011001: color_data = Z;
		19'b0111111010011011010: color_data = Z;
		19'b0111111010011011011: color_data = Z;
		19'b0111111010011101111: color_data = Z;
		19'b0111111010011110000: color_data = Z;
		19'b0111111010011110001: color_data = Z;
		19'b0111111010011110010: color_data = Z;
		19'b0111111010011110011: color_data = Z;
		19'b0111111010011110100: color_data = Z;
		19'b0111111010011110101: color_data = Z;
		19'b0111111010011110110: color_data = Z;
		19'b0111111010011110111: color_data = Z;
		19'b0111111010011111000: color_data = Z;
		19'b0111111010011111001: color_data = Z;
		19'b0111111010011111010: color_data = Z;
		19'b0111111010011111011: color_data = Z;
		19'b0111111010100001010: color_data = Z;
		19'b0111111010100001011: color_data = Z;
		19'b0111111010100001100: color_data = Z;
		19'b0111111010100001101: color_data = Z;
		19'b0111111010100001110: color_data = Z;
		19'b0111111010100001111: color_data = Z;
		19'b0111111010100010000: color_data = Z;
		19'b0111111010100010001: color_data = Z;
		19'b0111111010100010010: color_data = Z;
		19'b0111111010100010011: color_data = Z;
		19'b0111111010100010100: color_data = Z;
		19'b0111111010100010101: color_data = Z;
		19'b0111111010100010110: color_data = Z;
		19'b0111111010100010111: color_data = Z;
		19'b0111111010100011000: color_data = Z;
		19'b0111111010100011001: color_data = Z;
		19'b0111111010100011010: color_data = Z;
		19'b0111111010100011011: color_data = Z;
		19'b0111111010100011100: color_data = Z;
		19'b0111111010100011101: color_data = Z;
		19'b0111111010100011110: color_data = Z;
		19'b0111111010100011111: color_data = Z;
		19'b0111111010100100000: color_data = Z;
		19'b0111111010100100001: color_data = Z;
		19'b0111111010100100010: color_data = Z;
		19'b0111111010100100011: color_data = Z;
		19'b0111111010100100100: color_data = Z;
		19'b0111111010100100101: color_data = Z;
		19'b0111111010100100110: color_data = Z;
		19'b0111111010100100111: color_data = Z;
		19'b0111111010100101000: color_data = Z;
		19'b0111111010100101001: color_data = Z;
		19'b0111111010100101010: color_data = Z;
		19'b0111111010100101011: color_data = Z;
		19'b0111111010100101100: color_data = Z;
		19'b0111111010100101101: color_data = Z;
		19'b0111111010100101110: color_data = Z;
		19'b0111111010100110110: color_data = Z;
		19'b0111111010100110111: color_data = Z;
		19'b0111111010100111000: color_data = Z;
		19'b0111111010100111001: color_data = Z;
		19'b0111111010100111010: color_data = Z;
		19'b0111111010100111011: color_data = Z;
		19'b0111111010100111100: color_data = Z;
		19'b0111111010100111101: color_data = Z;
		19'b0111111010100111110: color_data = Z;
		19'b0111111010100111111: color_data = Z;
		19'b0111111010101000011: color_data = Z;
		19'b0111111010101000100: color_data = Z;
		19'b0111111010101000101: color_data = Z;
		19'b0111111010101000110: color_data = Z;
		19'b0111111010101000111: color_data = Z;
		19'b0111111010101001000: color_data = Z;
		19'b0111111010101001001: color_data = Z;
		19'b0111111010101001010: color_data = Z;
		19'b0111111010101001011: color_data = Z;
		19'b0111111010101001100: color_data = Z;
		19'b0111111010101001101: color_data = Z;
		19'b0111111010101001110: color_data = Z;
		19'b0111111010101001111: color_data = Z;
		19'b0111111010101010000: color_data = Z;
		19'b0111111010101010001: color_data = Z;
		19'b0111111010101010010: color_data = Z;
		19'b0111111010101010011: color_data = Z;
		19'b0111111010101010100: color_data = Z;
		19'b0111111010101010101: color_data = Z;
		19'b0111111010101010110: color_data = Z;
		19'b0111111010101010111: color_data = Z;
		19'b0111111010101011000: color_data = Z;
		19'b0111111010101011011: color_data = Z;
		19'b0111111010101011100: color_data = Z;
		19'b0111111010101011101: color_data = Z;
		19'b0111111010101011110: color_data = Z;
		19'b0111111010101011111: color_data = Z;
		19'b0111111010101100000: color_data = Z;
		19'b0111111010101100001: color_data = Z;
		19'b0111111010101100010: color_data = Z;
		19'b0111111010101100011: color_data = Z;
		19'b0111111010101100100: color_data = Z;
		19'b0111111010101100101: color_data = Z;
		19'b0111111010101100110: color_data = Z;
		19'b0111111010101101010: color_data = Z;
		19'b0111111010101101011: color_data = Z;
		19'b0111111010101101100: color_data = Z;
		19'b0111111010101101101: color_data = Z;
		19'b0111111010101101110: color_data = Z;
		19'b0111111010101101111: color_data = Z;
		19'b0111111010101110000: color_data = Z;
		19'b0111111010101110001: color_data = Z;
		19'b0111111010101110010: color_data = Z;
		19'b0111111010101110011: color_data = Z;
		19'b0111111010101110100: color_data = Z;
		19'b0111111010101110101: color_data = Z;
		19'b0111111010101110110: color_data = Z;
		19'b0111111010101110111: color_data = Z;
		19'b0111111010101111000: color_data = Z;
		19'b0111111010101111001: color_data = Z;
		19'b0111111010101111010: color_data = Z;
		19'b0111111010101111011: color_data = Z;
		19'b0111111010101111100: color_data = Z;
		19'b0111111010101111101: color_data = Z;
		19'b0111111010101111110: color_data = Z;
		19'b0111111010101111111: color_data = Z;
		19'b0111111010110000000: color_data = Z;
		19'b0111111010110000001: color_data = Z;
		19'b0111111010110000010: color_data = Z;
		19'b0111111010110000011: color_data = Z;
		19'b0111111010110000100: color_data = Z;
		19'b0111111010110000101: color_data = Z;
		19'b0111111010110000110: color_data = Z;
		19'b0111111010110000111: color_data = Z;
		19'b0111111010110001000: color_data = Z;
		19'b0111111010110001001: color_data = Z;
		19'b0111111010110001010: color_data = Z;
		19'b0111111010110001011: color_data = Z;
		19'b0111111010110001100: color_data = Z;
		19'b0111111010110001101: color_data = Z;
		19'b0111111010110001110: color_data = Z;
		19'b0111111010110001111: color_data = Z;
		19'b0111111010110010000: color_data = Z;
		19'b0111111010110010001: color_data = Z;
		19'b0111111010110010010: color_data = Z;
		19'b0111111010110010011: color_data = Z;
		19'b0111111010110010111: color_data = Z;
		19'b0111111010110011000: color_data = Z;
		19'b0111111010110011001: color_data = Z;
		19'b0111111010110011010: color_data = Z;
		19'b0111111010110011011: color_data = Z;
		19'b0111111010110011100: color_data = Z;
		19'b0111111010110011101: color_data = Z;
		19'b0111111010110011110: color_data = Z;
		19'b0111111010110011111: color_data = Z;
		19'b0111111010110100000: color_data = Z;
		19'b0111111010110100001: color_data = Z;
		19'b0111111010110100010: color_data = Z;
		19'b0111111010110100011: color_data = Z;
		19'b0111111010110100100: color_data = Z;
		19'b0111111010110100101: color_data = Z;
		19'b0111111010110100110: color_data = Z;
		19'b0111111010110100111: color_data = Z;
		19'b0111111010110101000: color_data = Z;
		19'b0111111010110101001: color_data = Z;
		19'b0111111010110101010: color_data = Z;
		19'b0111111010110101011: color_data = Z;
		19'b0111111010110101100: color_data = Z;
		19'b0111111010110101101: color_data = Z;
		19'b0111111010110101110: color_data = Z;
		19'b0111111010110101111: color_data = Z;
		19'b0111111010110110000: color_data = Z;
		19'b0111111010110110001: color_data = Z;
		19'b0111111010110110010: color_data = Z;
		19'b0111111010110110011: color_data = Z;
		19'b0111111010110110100: color_data = Z;
		19'b0111111010110110101: color_data = Z;
		19'b0111111010110110110: color_data = Z;
		19'b0111111010110110111: color_data = Z;
		19'b0111111010110111000: color_data = Z;
		19'b0111111010110111001: color_data = Z;
		19'b0111111010110111010: color_data = Z;
		19'b0111111010110111011: color_data = Z;
		19'b0111111010110111100: color_data = Z;
		19'b0111111010111000000: color_data = Z;
		19'b0111111010111000001: color_data = Z;
		19'b0111111010111000010: color_data = Z;
		19'b0111111010111000011: color_data = Z;
		19'b0111111010111000100: color_data = Z;
		19'b0111111010111000101: color_data = Z;
		19'b0111111010111000110: color_data = Z;
		19'b0111111010111000111: color_data = Z;
		19'b0111111010111001000: color_data = Z;
		19'b0111111100010110011: color_data = Z;
		19'b0111111100010110100: color_data = Z;
		19'b0111111100010110101: color_data = Z;
		19'b0111111100010110110: color_data = Z;
		19'b0111111100010110111: color_data = Z;
		19'b0111111100010111000: color_data = Z;
		19'b0111111100010111001: color_data = Z;
		19'b0111111100010111010: color_data = Z;
		19'b0111111100010111011: color_data = Z;
		19'b0111111100010111100: color_data = Z;
		19'b0111111100010111101: color_data = Z;
		19'b0111111100010111110: color_data = Z;
		19'b0111111100010111111: color_data = Z;
		19'b0111111100011000000: color_data = Z;
		19'b0111111100011000001: color_data = Z;
		19'b0111111100011000010: color_data = Z;
		19'b0111111100011000011: color_data = Z;
		19'b0111111100011000100: color_data = Z;
		19'b0111111100011000101: color_data = Z;
		19'b0111111100011001100: color_data = Z;
		19'b0111111100011001101: color_data = Z;
		19'b0111111100011010101: color_data = Z;
		19'b0111111100011010110: color_data = Z;
		19'b0111111100011010111: color_data = Z;
		19'b0111111100011011000: color_data = Z;
		19'b0111111100011011001: color_data = Z;
		19'b0111111100011011010: color_data = Z;
		19'b0111111100011011011: color_data = Z;
		19'b0111111100011011100: color_data = Z;
		19'b0111111100011011101: color_data = Z;
		19'b0111111100011101110: color_data = Z;
		19'b0111111100011101111: color_data = Z;
		19'b0111111100011110000: color_data = Z;
		19'b0111111100011110001: color_data = Z;
		19'b0111111100011110010: color_data = Z;
		19'b0111111100011110011: color_data = Z;
		19'b0111111100011110100: color_data = Z;
		19'b0111111100011110101: color_data = Z;
		19'b0111111100011110110: color_data = Z;
		19'b0111111100011110111: color_data = Z;
		19'b0111111100011111000: color_data = Z;
		19'b0111111100011111001: color_data = Z;
		19'b0111111100011111010: color_data = Z;
		19'b0111111100011111011: color_data = Z;
		19'b0111111100011111100: color_data = Z;
		19'b0111111100100001001: color_data = Z;
		19'b0111111100100001010: color_data = Z;
		19'b0111111100100001011: color_data = Z;
		19'b0111111100100001100: color_data = Z;
		19'b0111111100100001101: color_data = Z;
		19'b0111111100100001110: color_data = Z;
		19'b0111111100100001111: color_data = Z;
		19'b0111111100100010000: color_data = Z;
		19'b0111111100100010001: color_data = Z;
		19'b0111111100100010010: color_data = Z;
		19'b0111111100100010011: color_data = Z;
		19'b0111111100100010100: color_data = Z;
		19'b0111111100100010101: color_data = Z;
		19'b0111111100100010110: color_data = Z;
		19'b0111111100100010111: color_data = Z;
		19'b0111111100100011000: color_data = Z;
		19'b0111111100100011001: color_data = Z;
		19'b0111111100100011010: color_data = Z;
		19'b0111111100100011011: color_data = Z;
		19'b0111111100100011100: color_data = Z;
		19'b0111111100100011101: color_data = Z;
		19'b0111111100100011110: color_data = Z;
		19'b0111111100100011111: color_data = Z;
		19'b0111111100100100000: color_data = Z;
		19'b0111111100100100001: color_data = Z;
		19'b0111111100100100010: color_data = Z;
		19'b0111111100100100011: color_data = Z;
		19'b0111111100100100100: color_data = Z;
		19'b0111111100100100101: color_data = Z;
		19'b0111111100100100110: color_data = Z;
		19'b0111111100100100111: color_data = Z;
		19'b0111111100100101000: color_data = Z;
		19'b0111111100100101001: color_data = Z;
		19'b0111111100100101010: color_data = Z;
		19'b0111111100100101011: color_data = Z;
		19'b0111111100100101100: color_data = Z;
		19'b0111111100100101101: color_data = Z;
		19'b0111111100100101110: color_data = Z;
		19'b0111111100100110110: color_data = Z;
		19'b0111111100100110111: color_data = Z;
		19'b0111111100100111000: color_data = Z;
		19'b0111111100100111001: color_data = Z;
		19'b0111111100100111010: color_data = Z;
		19'b0111111100100111011: color_data = Z;
		19'b0111111100100111100: color_data = Z;
		19'b0111111100100111101: color_data = Z;
		19'b0111111100100111110: color_data = Z;
		19'b0111111100100111111: color_data = Z;
		19'b0111111100101000100: color_data = Z;
		19'b0111111100101000101: color_data = Z;
		19'b0111111100101000110: color_data = Z;
		19'b0111111100101000111: color_data = Z;
		19'b0111111100101001000: color_data = Z;
		19'b0111111100101001001: color_data = Z;
		19'b0111111100101001010: color_data = Z;
		19'b0111111100101001011: color_data = Z;
		19'b0111111100101001100: color_data = Z;
		19'b0111111100101001101: color_data = Z;
		19'b0111111100101001110: color_data = Z;
		19'b0111111100101001111: color_data = Z;
		19'b0111111100101010000: color_data = Z;
		19'b0111111100101010001: color_data = Z;
		19'b0111111100101010010: color_data = Z;
		19'b0111111100101010011: color_data = Z;
		19'b0111111100101010100: color_data = Z;
		19'b0111111100101010101: color_data = Z;
		19'b0111111100101010110: color_data = Z;
		19'b0111111100101010111: color_data = Z;
		19'b0111111100101011000: color_data = Z;
		19'b0111111100101011100: color_data = Z;
		19'b0111111100101011101: color_data = Z;
		19'b0111111100101011110: color_data = Z;
		19'b0111111100101011111: color_data = Z;
		19'b0111111100101100000: color_data = Z;
		19'b0111111100101100001: color_data = Z;
		19'b0111111100101100010: color_data = Z;
		19'b0111111100101100011: color_data = Z;
		19'b0111111100101100100: color_data = Z;
		19'b0111111100101100101: color_data = Z;
		19'b0111111100101101010: color_data = Z;
		19'b0111111100101101011: color_data = Z;
		19'b0111111100101101100: color_data = Z;
		19'b0111111100101101101: color_data = Z;
		19'b0111111100101101110: color_data = Z;
		19'b0111111100101101111: color_data = Z;
		19'b0111111100101110000: color_data = Z;
		19'b0111111100101110001: color_data = Z;
		19'b0111111100101110010: color_data = Z;
		19'b0111111100101110011: color_data = Z;
		19'b0111111100101110100: color_data = Z;
		19'b0111111100101110101: color_data = Z;
		19'b0111111100101110110: color_data = Z;
		19'b0111111100101110111: color_data = Z;
		19'b0111111100101111000: color_data = Z;
		19'b0111111100101111001: color_data = Z;
		19'b0111111100101111010: color_data = Z;
		19'b0111111100101111011: color_data = Z;
		19'b0111111100101111100: color_data = Z;
		19'b0111111100101111101: color_data = Z;
		19'b0111111100101111110: color_data = Z;
		19'b0111111100101111111: color_data = Z;
		19'b0111111100110000000: color_data = Z;
		19'b0111111100110000001: color_data = Z;
		19'b0111111100110000010: color_data = Z;
		19'b0111111100110000011: color_data = Z;
		19'b0111111100110000100: color_data = Z;
		19'b0111111100110000101: color_data = Z;
		19'b0111111100110000110: color_data = Z;
		19'b0111111100110000111: color_data = Z;
		19'b0111111100110001000: color_data = Z;
		19'b0111111100110001001: color_data = Z;
		19'b0111111100110001010: color_data = Z;
		19'b0111111100110001011: color_data = Z;
		19'b0111111100110001100: color_data = Z;
		19'b0111111100110001101: color_data = Z;
		19'b0111111100110001110: color_data = Z;
		19'b0111111100110001111: color_data = Z;
		19'b0111111100110010000: color_data = Z;
		19'b0111111100110010001: color_data = Z;
		19'b0111111100110010010: color_data = Z;
		19'b0111111100110010011: color_data = Z;
		19'b0111111100110010100: color_data = Z;
		19'b0111111100110010101: color_data = Z;
		19'b0111111100110011000: color_data = Z;
		19'b0111111100110011001: color_data = Z;
		19'b0111111100110011010: color_data = Z;
		19'b0111111100110011011: color_data = Z;
		19'b0111111100110011100: color_data = Z;
		19'b0111111100110011101: color_data = Z;
		19'b0111111100110011110: color_data = Z;
		19'b0111111100110011111: color_data = Z;
		19'b0111111100110100000: color_data = Z;
		19'b0111111100110100001: color_data = Z;
		19'b0111111100110100010: color_data = Z;
		19'b0111111100110100011: color_data = Z;
		19'b0111111100110100100: color_data = Z;
		19'b0111111100110100101: color_data = Z;
		19'b0111111100110100110: color_data = Z;
		19'b0111111100110100111: color_data = Z;
		19'b0111111100110101000: color_data = Z;
		19'b0111111100110101001: color_data = Z;
		19'b0111111100110101010: color_data = Z;
		19'b0111111100110101011: color_data = Z;
		19'b0111111100110101100: color_data = Z;
		19'b0111111100110101101: color_data = Z;
		19'b0111111100110101110: color_data = Z;
		19'b0111111100110101111: color_data = Z;
		19'b0111111100110110000: color_data = Z;
		19'b0111111100110110001: color_data = Z;
		19'b0111111100110110010: color_data = Z;
		19'b0111111100110110011: color_data = Z;
		19'b0111111100110110100: color_data = Z;
		19'b0111111100110110101: color_data = Z;
		19'b0111111100110110110: color_data = Z;
		19'b0111111100110110111: color_data = Z;
		19'b0111111100110111000: color_data = Z;
		19'b0111111100110111001: color_data = Z;
		19'b0111111100110111010: color_data = Z;
		19'b0111111100110111011: color_data = Z;
		19'b0111111100110111100: color_data = Z;
		19'b0111111100111000000: color_data = Z;
		19'b0111111100111000001: color_data = Z;
		19'b0111111100111000010: color_data = Z;
		19'b0111111100111000011: color_data = Z;
		19'b0111111100111000100: color_data = Z;
		19'b0111111100111000101: color_data = Z;
		19'b0111111100111000110: color_data = Z;
		19'b0111111100111000111: color_data = Z;
		19'b0111111100111001000: color_data = Z;
		19'b0111111110010110100: color_data = Z;
		19'b0111111110010110101: color_data = Z;
		19'b0111111110010110110: color_data = Z;
		19'b0111111110010110111: color_data = Z;
		19'b0111111110010111000: color_data = Z;
		19'b0111111110010111001: color_data = Z;
		19'b0111111110010111010: color_data = Z;
		19'b0111111110010111011: color_data = Z;
		19'b0111111110010111100: color_data = Z;
		19'b0111111110010111101: color_data = Z;
		19'b0111111110010111110: color_data = Z;
		19'b0111111110010111111: color_data = Z;
		19'b0111111110011000000: color_data = Z;
		19'b0111111110011000001: color_data = Z;
		19'b0111111110011000010: color_data = Z;
		19'b0111111110011000011: color_data = Z;
		19'b0111111110011000100: color_data = Z;
		19'b0111111110011000101: color_data = Z;
		19'b0111111110011000110: color_data = Z;
		19'b0111111110011001101: color_data = Z;
		19'b0111111110011001110: color_data = Z;
		19'b0111111110011010010: color_data = Z;
		19'b0111111110011010011: color_data = Z;
		19'b0111111110011010100: color_data = Z;
		19'b0111111110011010101: color_data = Z;
		19'b0111111110011010110: color_data = Z;
		19'b0111111110011010111: color_data = Z;
		19'b0111111110011011000: color_data = Z;
		19'b0111111110011011001: color_data = Z;
		19'b0111111110011011010: color_data = Z;
		19'b0111111110011011011: color_data = Z;
		19'b0111111110011011100: color_data = Z;
		19'b0111111110011011101: color_data = Z;
		19'b0111111110011101100: color_data = Z;
		19'b0111111110011101101: color_data = Z;
		19'b0111111110011101110: color_data = Z;
		19'b0111111110011101111: color_data = Z;
		19'b0111111110011110000: color_data = Z;
		19'b0111111110011110001: color_data = Z;
		19'b0111111110011110010: color_data = Z;
		19'b0111111110011110011: color_data = Z;
		19'b0111111110011110100: color_data = Z;
		19'b0111111110011110101: color_data = Z;
		19'b0111111110011110110: color_data = Z;
		19'b0111111110011110111: color_data = Z;
		19'b0111111110011111000: color_data = Z;
		19'b0111111110011111001: color_data = Z;
		19'b0111111110011111010: color_data = Z;
		19'b0111111110011111011: color_data = Z;
		19'b0111111110011111100: color_data = Z;
		19'b0111111110011111101: color_data = Z;
		19'b0111111110100001000: color_data = Z;
		19'b0111111110100001001: color_data = Z;
		19'b0111111110100001010: color_data = Z;
		19'b0111111110100001011: color_data = Z;
		19'b0111111110100001100: color_data = Z;
		19'b0111111110100001101: color_data = Z;
		19'b0111111110100001110: color_data = Z;
		19'b0111111110100001111: color_data = Z;
		19'b0111111110100010000: color_data = Z;
		19'b0111111110100010001: color_data = Z;
		19'b0111111110100010010: color_data = Z;
		19'b0111111110100010011: color_data = Z;
		19'b0111111110100010100: color_data = Z;
		19'b0111111110100010101: color_data = Z;
		19'b0111111110100010110: color_data = Z;
		19'b0111111110100010111: color_data = Z;
		19'b0111111110100011000: color_data = Z;
		19'b0111111110100011001: color_data = Z;
		19'b0111111110100011010: color_data = Z;
		19'b0111111110100011011: color_data = Z;
		19'b0111111110100011100: color_data = Z;
		19'b0111111110100011101: color_data = Z;
		19'b0111111110100011110: color_data = Z;
		19'b0111111110100011111: color_data = Z;
		19'b0111111110100100000: color_data = Z;
		19'b0111111110100100001: color_data = Z;
		19'b0111111110100100010: color_data = Z;
		19'b0111111110100100011: color_data = Z;
		19'b0111111110100100100: color_data = Z;
		19'b0111111110100100101: color_data = Z;
		19'b0111111110100100110: color_data = Z;
		19'b0111111110100100111: color_data = Z;
		19'b0111111110100101000: color_data = Z;
		19'b0111111110100101001: color_data = Z;
		19'b0111111110100101010: color_data = Z;
		19'b0111111110100101011: color_data = Z;
		19'b0111111110100101100: color_data = Z;
		19'b0111111110100101101: color_data = Z;
		19'b0111111110100101110: color_data = Z;
		19'b0111111110100110110: color_data = Z;
		19'b0111111110100110111: color_data = Z;
		19'b0111111110100111000: color_data = Z;
		19'b0111111110100111001: color_data = Z;
		19'b0111111110100111010: color_data = Z;
		19'b0111111110100111011: color_data = Z;
		19'b0111111110100111100: color_data = Z;
		19'b0111111110100111101: color_data = Z;
		19'b0111111110100111110: color_data = Z;
		19'b0111111110100111111: color_data = Z;
		19'b0111111110101000100: color_data = Z;
		19'b0111111110101000101: color_data = Z;
		19'b0111111110101000110: color_data = Z;
		19'b0111111110101000111: color_data = Z;
		19'b0111111110101001000: color_data = Z;
		19'b0111111110101001001: color_data = Z;
		19'b0111111110101001010: color_data = Z;
		19'b0111111110101001011: color_data = Z;
		19'b0111111110101001100: color_data = Z;
		19'b0111111110101001101: color_data = Z;
		19'b0111111110101001110: color_data = Z;
		19'b0111111110101001111: color_data = Z;
		19'b0111111110101010000: color_data = Z;
		19'b0111111110101010001: color_data = Z;
		19'b0111111110101010010: color_data = Z;
		19'b0111111110101010011: color_data = Z;
		19'b0111111110101010100: color_data = Z;
		19'b0111111110101010101: color_data = Z;
		19'b0111111110101010110: color_data = Z;
		19'b0111111110101010111: color_data = Z;
		19'b0111111110101011100: color_data = Z;
		19'b0111111110101011101: color_data = Z;
		19'b0111111110101011110: color_data = Z;
		19'b0111111110101011111: color_data = Z;
		19'b0111111110101100000: color_data = Z;
		19'b0111111110101100001: color_data = Z;
		19'b0111111110101100010: color_data = Z;
		19'b0111111110101100011: color_data = Z;
		19'b0111111110101100100: color_data = Z;
		19'b0111111110101100101: color_data = Z;
		19'b0111111110101101011: color_data = Z;
		19'b0111111110101101100: color_data = Z;
		19'b0111111110101101101: color_data = Z;
		19'b0111111110101101110: color_data = Z;
		19'b0111111110101101111: color_data = Z;
		19'b0111111110101110000: color_data = Z;
		19'b0111111110101110001: color_data = Z;
		19'b0111111110101110010: color_data = Z;
		19'b0111111110101110011: color_data = Z;
		19'b0111111110101110100: color_data = Z;
		19'b0111111110101110101: color_data = Z;
		19'b0111111110101110110: color_data = Z;
		19'b0111111110101110111: color_data = Z;
		19'b0111111110101111000: color_data = Z;
		19'b0111111110101111001: color_data = Z;
		19'b0111111110101111010: color_data = Z;
		19'b0111111110101111011: color_data = Z;
		19'b0111111110101111100: color_data = Z;
		19'b0111111110101111101: color_data = Z;
		19'b0111111110101111110: color_data = Z;
		19'b0111111110101111111: color_data = Z;
		19'b0111111110110000000: color_data = Z;
		19'b0111111110110000001: color_data = Z;
		19'b0111111110110000010: color_data = Z;
		19'b0111111110110000011: color_data = Z;
		19'b0111111110110000100: color_data = Z;
		19'b0111111110110000101: color_data = Z;
		19'b0111111110110000110: color_data = Z;
		19'b0111111110110000111: color_data = Z;
		19'b0111111110110001000: color_data = Z;
		19'b0111111110110001001: color_data = Z;
		19'b0111111110110001010: color_data = Z;
		19'b0111111110110001011: color_data = Z;
		19'b0111111110110001110: color_data = Z;
		19'b0111111110110001111: color_data = Z;
		19'b0111111110110010000: color_data = Z;
		19'b0111111110110010001: color_data = Z;
		19'b0111111110110010010: color_data = Z;
		19'b0111111110110010011: color_data = Z;
		19'b0111111110110010100: color_data = Z;
		19'b0111111110110010101: color_data = Z;
		19'b0111111110110010110: color_data = Z;
		19'b0111111110110010111: color_data = Z;
		19'b0111111110110011000: color_data = Z;
		19'b0111111110110011001: color_data = Z;
		19'b0111111110110011010: color_data = Z;
		19'b0111111110110011011: color_data = Z;
		19'b0111111110110011100: color_data = Z;
		19'b0111111110110011101: color_data = Z;
		19'b0111111110110011110: color_data = Z;
		19'b0111111110110011111: color_data = Z;
		19'b0111111110110100000: color_data = Z;
		19'b0111111110110100001: color_data = Z;
		19'b0111111110110100010: color_data = Z;
		19'b0111111110110100011: color_data = Z;
		19'b0111111110110100100: color_data = Z;
		19'b0111111110110100101: color_data = Z;
		19'b0111111110110100110: color_data = Z;
		19'b0111111110110100111: color_data = Z;
		19'b0111111110110101000: color_data = Z;
		19'b0111111110110101001: color_data = Z;
		19'b0111111110110101010: color_data = Z;
		19'b0111111110110101011: color_data = Z;
		19'b0111111110110101100: color_data = Z;
		19'b0111111110110101101: color_data = Z;
		19'b0111111110110101110: color_data = Z;
		19'b0111111110110101111: color_data = Z;
		19'b0111111110110110000: color_data = Z;
		19'b0111111110110110001: color_data = Z;
		19'b0111111110110110010: color_data = Z;
		19'b0111111110110110011: color_data = Z;
		19'b0111111110110110100: color_data = Z;
		19'b0111111110110110101: color_data = Z;
		19'b0111111110110110110: color_data = Z;
		19'b0111111110110110111: color_data = Z;
		19'b0111111110110111000: color_data = Z;
		19'b0111111110110111001: color_data = Z;
		19'b0111111110110111010: color_data = Z;
		19'b0111111110110111011: color_data = Z;
		19'b0111111110110111100: color_data = Z;
		19'b0111111110111000000: color_data = Z;
		19'b0111111110111000001: color_data = Z;
		19'b0111111110111000010: color_data = Z;
		19'b0111111110111000011: color_data = Z;
		19'b0111111110111000100: color_data = Z;
		19'b0111111110111000101: color_data = Z;
		19'b0111111110111000110: color_data = Z;
		19'b0111111110111000111: color_data = Z;
		19'b0111111110111001000: color_data = Z;
		19'b0111111110111001001: color_data = Z;
		19'b1000000000010110100: color_data = Z;
		19'b1000000000010110101: color_data = Z;
		19'b1000000000010110110: color_data = Z;
		19'b1000000000010110111: color_data = Z;
		19'b1000000000010111000: color_data = Z;
		19'b1000000000010111001: color_data = Z;
		19'b1000000000010111010: color_data = Z;
		19'b1000000000010111011: color_data = Z;
		19'b1000000000010111100: color_data = Z;
		19'b1000000000010111101: color_data = Z;
		19'b1000000000010111110: color_data = Z;
		19'b1000000000010111111: color_data = Z;
		19'b1000000000011000000: color_data = Z;
		19'b1000000000011000001: color_data = Z;
		19'b1000000000011000010: color_data = Z;
		19'b1000000000011000011: color_data = Z;
		19'b1000000000011000100: color_data = Z;
		19'b1000000000011000101: color_data = Z;
		19'b1000000000011000110: color_data = Z;
		19'b1000000000011000111: color_data = Z;
		19'b1000000000011001110: color_data = Z;
		19'b1000000000011001111: color_data = Z;
		19'b1000000000011010010: color_data = Z;
		19'b1000000000011010011: color_data = Z;
		19'b1000000000011010100: color_data = Z;
		19'b1000000000011010101: color_data = Z;
		19'b1000000000011010110: color_data = Z;
		19'b1000000000011010111: color_data = Z;
		19'b1000000000011011000: color_data = Z;
		19'b1000000000011011001: color_data = Z;
		19'b1000000000011011010: color_data = Z;
		19'b1000000000011011011: color_data = Z;
		19'b1000000000011011100: color_data = Z;
		19'b1000000000011011101: color_data = Z;
		19'b1000000000011011110: color_data = Z;
		19'b1000000000011101011: color_data = Z;
		19'b1000000000011101100: color_data = Z;
		19'b1000000000011101101: color_data = Z;
		19'b1000000000011101110: color_data = Z;
		19'b1000000000011101111: color_data = Z;
		19'b1000000000011110000: color_data = Z;
		19'b1000000000011110001: color_data = Z;
		19'b1000000000011110010: color_data = Z;
		19'b1000000000011110011: color_data = Z;
		19'b1000000000011110100: color_data = Z;
		19'b1000000000011110101: color_data = Z;
		19'b1000000000011110110: color_data = Z;
		19'b1000000000011110111: color_data = Z;
		19'b1000000000011111000: color_data = Z;
		19'b1000000000011111001: color_data = Z;
		19'b1000000000011111010: color_data = Z;
		19'b1000000000011111011: color_data = Z;
		19'b1000000000011111100: color_data = Z;
		19'b1000000000100001000: color_data = Z;
		19'b1000000000100001001: color_data = Z;
		19'b1000000000100001010: color_data = Z;
		19'b1000000000100001011: color_data = Z;
		19'b1000000000100001100: color_data = Z;
		19'b1000000000100001101: color_data = Z;
		19'b1000000000100001110: color_data = Z;
		19'b1000000000100001111: color_data = Z;
		19'b1000000000100010000: color_data = Z;
		19'b1000000000100010001: color_data = Z;
		19'b1000000000100010010: color_data = Z;
		19'b1000000000100010011: color_data = Z;
		19'b1000000000100010100: color_data = Z;
		19'b1000000000100010101: color_data = Z;
		19'b1000000000100010110: color_data = Z;
		19'b1000000000100010111: color_data = Z;
		19'b1000000000100011000: color_data = Z;
		19'b1000000000100011001: color_data = Z;
		19'b1000000000100011010: color_data = Z;
		19'b1000000000100011011: color_data = Z;
		19'b1000000000100011100: color_data = Z;
		19'b1000000000100011101: color_data = Z;
		19'b1000000000100011110: color_data = Z;
		19'b1000000000100011111: color_data = Z;
		19'b1000000000100100000: color_data = Z;
		19'b1000000000100100001: color_data = Z;
		19'b1000000000100100010: color_data = Z;
		19'b1000000000100100011: color_data = Z;
		19'b1000000000100100100: color_data = Z;
		19'b1000000000100100101: color_data = Z;
		19'b1000000000100100110: color_data = Z;
		19'b1000000000100100111: color_data = Z;
		19'b1000000000100101000: color_data = Z;
		19'b1000000000100101001: color_data = Z;
		19'b1000000000100101010: color_data = Z;
		19'b1000000000100101011: color_data = Z;
		19'b1000000000100101100: color_data = Z;
		19'b1000000000100101101: color_data = Z;
		19'b1000000000100101110: color_data = Z;
		19'b1000000000100110111: color_data = Z;
		19'b1000000000100111000: color_data = Z;
		19'b1000000000100111001: color_data = Z;
		19'b1000000000100111010: color_data = Z;
		19'b1000000000100111011: color_data = Z;
		19'b1000000000100111100: color_data = Z;
		19'b1000000000100111101: color_data = Z;
		19'b1000000000100111110: color_data = Z;
		19'b1000000000100111111: color_data = Z;
		19'b1000000000101000101: color_data = Z;
		19'b1000000000101000110: color_data = Z;
		19'b1000000000101000111: color_data = Z;
		19'b1000000000101001000: color_data = Z;
		19'b1000000000101001001: color_data = Z;
		19'b1000000000101001010: color_data = Z;
		19'b1000000000101001011: color_data = Z;
		19'b1000000000101001100: color_data = Z;
		19'b1000000000101001101: color_data = Z;
		19'b1000000000101001110: color_data = Z;
		19'b1000000000101001111: color_data = Z;
		19'b1000000000101010000: color_data = Z;
		19'b1000000000101010001: color_data = Z;
		19'b1000000000101010010: color_data = Z;
		19'b1000000000101010011: color_data = Z;
		19'b1000000000101010100: color_data = Z;
		19'b1000000000101010101: color_data = Z;
		19'b1000000000101010110: color_data = Z;
		19'b1000000000101010111: color_data = Z;
		19'b1000000000101011100: color_data = Z;
		19'b1000000000101011101: color_data = Z;
		19'b1000000000101011110: color_data = Z;
		19'b1000000000101011111: color_data = Z;
		19'b1000000000101100000: color_data = Z;
		19'b1000000000101100001: color_data = Z;
		19'b1000000000101100010: color_data = Z;
		19'b1000000000101100011: color_data = Z;
		19'b1000000000101100100: color_data = Z;
		19'b1000000000101100101: color_data = Z;
		19'b1000000000101101010: color_data = Z;
		19'b1000000000101101011: color_data = Z;
		19'b1000000000101101100: color_data = Z;
		19'b1000000000101101101: color_data = Z;
		19'b1000000000101101110: color_data = Z;
		19'b1000000000101101111: color_data = Z;
		19'b1000000000101110000: color_data = Z;
		19'b1000000000101110001: color_data = Z;
		19'b1000000000101110010: color_data = Z;
		19'b1000000000101110011: color_data = Z;
		19'b1000000000101110100: color_data = Z;
		19'b1000000000101110101: color_data = Z;
		19'b1000000000101110110: color_data = Z;
		19'b1000000000101110111: color_data = Z;
		19'b1000000000101111000: color_data = Z;
		19'b1000000000101111001: color_data = Z;
		19'b1000000000101111010: color_data = Z;
		19'b1000000000101111011: color_data = Z;
		19'b1000000000101111100: color_data = Z;
		19'b1000000000101111101: color_data = Z;
		19'b1000000000101111110: color_data = Z;
		19'b1000000000101111111: color_data = Z;
		19'b1000000000110000000: color_data = Z;
		19'b1000000000110000001: color_data = Z;
		19'b1000000000110000010: color_data = Z;
		19'b1000000000110000011: color_data = Z;
		19'b1000000000110000100: color_data = Z;
		19'b1000000000110000101: color_data = Z;
		19'b1000000000110000110: color_data = Z;
		19'b1000000000110000111: color_data = Z;
		19'b1000000000110001000: color_data = Z;
		19'b1000000000110001001: color_data = Z;
		19'b1000000000110001010: color_data = Z;
		19'b1000000000110001011: color_data = Z;
		19'b1000000000110001100: color_data = Z;
		19'b1000000000110010000: color_data = Z;
		19'b1000000000110010001: color_data = Z;
		19'b1000000000110010010: color_data = Z;
		19'b1000000000110010011: color_data = Z;
		19'b1000000000110010100: color_data = Z;
		19'b1000000000110010101: color_data = Z;
		19'b1000000000110010110: color_data = Z;
		19'b1000000000110010111: color_data = Z;
		19'b1000000000110011000: color_data = Z;
		19'b1000000000110011001: color_data = Z;
		19'b1000000000110011010: color_data = Z;
		19'b1000000000110011011: color_data = Z;
		19'b1000000000110011100: color_data = Z;
		19'b1000000000110011101: color_data = Z;
		19'b1000000000110011110: color_data = Z;
		19'b1000000000110011111: color_data = Z;
		19'b1000000000110100000: color_data = Z;
		19'b1000000000110100001: color_data = Z;
		19'b1000000000110100010: color_data = Z;
		19'b1000000000110100011: color_data = Z;
		19'b1000000000110100100: color_data = Z;
		19'b1000000000110100101: color_data = Z;
		19'b1000000000110100110: color_data = Z;
		19'b1000000000110100111: color_data = Z;
		19'b1000000000110101000: color_data = Z;
		19'b1000000000110101001: color_data = Z;
		19'b1000000000110101010: color_data = Z;
		19'b1000000000110101011: color_data = Z;
		19'b1000000000110101100: color_data = Z;
		19'b1000000000110101101: color_data = Z;
		19'b1000000000110101110: color_data = Z;
		19'b1000000000110101111: color_data = Z;
		19'b1000000000110110000: color_data = Z;
		19'b1000000000110110001: color_data = Z;
		19'b1000000000110110010: color_data = Z;
		19'b1000000000110110011: color_data = Z;
		19'b1000000000110110100: color_data = Z;
		19'b1000000000110110101: color_data = Z;
		19'b1000000000110110110: color_data = Z;
		19'b1000000000110110111: color_data = Z;
		19'b1000000000110111000: color_data = Z;
		19'b1000000000110111001: color_data = Z;
		19'b1000000000110111010: color_data = Z;
		19'b1000000000110111011: color_data = Z;
		19'b1000000000110111100: color_data = Z;
		19'b1000000000111000001: color_data = Z;
		19'b1000000000111000010: color_data = Z;
		19'b1000000000111000011: color_data = Z;
		19'b1000000000111000100: color_data = Z;
		19'b1000000000111000101: color_data = Z;
		19'b1000000000111000110: color_data = Z;
		19'b1000000000111000111: color_data = Z;
		19'b1000000000111001000: color_data = Z;
		19'b1000000000111001001: color_data = Z;
		19'b1000000010010110101: color_data = Z;
		19'b1000000010010110110: color_data = Z;
		19'b1000000010010110111: color_data = Z;
		19'b1000000010010111000: color_data = Z;
		19'b1000000010010111001: color_data = Z;
		19'b1000000010010111010: color_data = Z;
		19'b1000000010010111011: color_data = Z;
		19'b1000000010010111100: color_data = Z;
		19'b1000000010010111101: color_data = Z;
		19'b1000000010010111110: color_data = Z;
		19'b1000000010010111111: color_data = Z;
		19'b1000000010011000000: color_data = Z;
		19'b1000000010011000001: color_data = Z;
		19'b1000000010011000010: color_data = Z;
		19'b1000000010011000011: color_data = Z;
		19'b1000000010011000100: color_data = Z;
		19'b1000000010011000101: color_data = Z;
		19'b1000000010011000110: color_data = Z;
		19'b1000000010011000111: color_data = Z;
		19'b1000000010011001000: color_data = Z;
		19'b1000000010011001111: color_data = Z;
		19'b1000000010011010000: color_data = Z;
		19'b1000000010011010001: color_data = Z;
		19'b1000000010011010010: color_data = Z;
		19'b1000000010011010011: color_data = Z;
		19'b1000000010011010100: color_data = Z;
		19'b1000000010011010101: color_data = Z;
		19'b1000000010011010110: color_data = Z;
		19'b1000000010011010111: color_data = Z;
		19'b1000000010011011000: color_data = Z;
		19'b1000000010011011001: color_data = Z;
		19'b1000000010011011010: color_data = Z;
		19'b1000000010011011011: color_data = Z;
		19'b1000000010011011100: color_data = Z;
		19'b1000000010011011101: color_data = Z;
		19'b1000000010011011110: color_data = Z;
		19'b1000000010011011111: color_data = Z;
		19'b1000000010011100000: color_data = Z;
		19'b1000000010011101011: color_data = Z;
		19'b1000000010011101100: color_data = Z;
		19'b1000000010011101101: color_data = Z;
		19'b1000000010011101110: color_data = Z;
		19'b1000000010011101111: color_data = Z;
		19'b1000000010011110000: color_data = Z;
		19'b1000000010011110001: color_data = Z;
		19'b1000000010011110010: color_data = Z;
		19'b1000000010011110011: color_data = Z;
		19'b1000000010011110100: color_data = Z;
		19'b1000000010011110101: color_data = Z;
		19'b1000000010011110110: color_data = Z;
		19'b1000000010011110111: color_data = Z;
		19'b1000000010011111000: color_data = Z;
		19'b1000000010011111001: color_data = Z;
		19'b1000000010011111010: color_data = Z;
		19'b1000000010011111011: color_data = Z;
		19'b1000000010100000111: color_data = Z;
		19'b1000000010100001000: color_data = Z;
		19'b1000000010100001001: color_data = Z;
		19'b1000000010100001010: color_data = Z;
		19'b1000000010100001011: color_data = Z;
		19'b1000000010100001100: color_data = Z;
		19'b1000000010100001101: color_data = Z;
		19'b1000000010100001110: color_data = Z;
		19'b1000000010100001111: color_data = Z;
		19'b1000000010100010000: color_data = Z;
		19'b1000000010100010001: color_data = Z;
		19'b1000000010100010010: color_data = Z;
		19'b1000000010100010011: color_data = Z;
		19'b1000000010100010100: color_data = Z;
		19'b1000000010100010101: color_data = Z;
		19'b1000000010100010110: color_data = Z;
		19'b1000000010100010111: color_data = Z;
		19'b1000000010100011000: color_data = Z;
		19'b1000000010100011001: color_data = Z;
		19'b1000000010100011010: color_data = Z;
		19'b1000000010100011011: color_data = Z;
		19'b1000000010100011100: color_data = Z;
		19'b1000000010100011101: color_data = Z;
		19'b1000000010100011110: color_data = Z;
		19'b1000000010100011111: color_data = Z;
		19'b1000000010100100000: color_data = Z;
		19'b1000000010100100001: color_data = Z;
		19'b1000000010100100010: color_data = Z;
		19'b1000000010100100011: color_data = Z;
		19'b1000000010100100100: color_data = Z;
		19'b1000000010100100101: color_data = Z;
		19'b1000000010100100110: color_data = Z;
		19'b1000000010100100111: color_data = Z;
		19'b1000000010100101000: color_data = Z;
		19'b1000000010100101001: color_data = Z;
		19'b1000000010100101010: color_data = Z;
		19'b1000000010100101011: color_data = Z;
		19'b1000000010100101100: color_data = Z;
		19'b1000000010100101101: color_data = Z;
		19'b1000000010100101110: color_data = Z;
		19'b1000000010100110111: color_data = Z;
		19'b1000000010100111000: color_data = Z;
		19'b1000000010100111001: color_data = Z;
		19'b1000000010100111010: color_data = Z;
		19'b1000000010100111011: color_data = Z;
		19'b1000000010100111100: color_data = Z;
		19'b1000000010100111101: color_data = Z;
		19'b1000000010100111110: color_data = Z;
		19'b1000000010100111111: color_data = Z;
		19'b1000000010101000110: color_data = Z;
		19'b1000000010101000111: color_data = Z;
		19'b1000000010101001000: color_data = Z;
		19'b1000000010101001001: color_data = Z;
		19'b1000000010101001010: color_data = Z;
		19'b1000000010101001011: color_data = Z;
		19'b1000000010101001100: color_data = Z;
		19'b1000000010101001101: color_data = Z;
		19'b1000000010101001110: color_data = Z;
		19'b1000000010101001111: color_data = Z;
		19'b1000000010101010000: color_data = Z;
		19'b1000000010101010001: color_data = Z;
		19'b1000000010101010010: color_data = Z;
		19'b1000000010101010011: color_data = Z;
		19'b1000000010101010100: color_data = Z;
		19'b1000000010101010101: color_data = Z;
		19'b1000000010101010110: color_data = Z;
		19'b1000000010101010111: color_data = Z;
		19'b1000000010101011101: color_data = Z;
		19'b1000000010101011110: color_data = Z;
		19'b1000000010101011111: color_data = Z;
		19'b1000000010101100000: color_data = Z;
		19'b1000000010101100001: color_data = Z;
		19'b1000000010101100010: color_data = Z;
		19'b1000000010101100011: color_data = Z;
		19'b1000000010101100100: color_data = Z;
		19'b1000000010101100101: color_data = Z;
		19'b1000000010101101010: color_data = Z;
		19'b1000000010101101011: color_data = Z;
		19'b1000000010101101100: color_data = Z;
		19'b1000000010101101101: color_data = Z;
		19'b1000000010101101110: color_data = Z;
		19'b1000000010101101111: color_data = Z;
		19'b1000000010101110000: color_data = Z;
		19'b1000000010101110001: color_data = Z;
		19'b1000000010101110010: color_data = Z;
		19'b1000000010101110011: color_data = Z;
		19'b1000000010101110100: color_data = Z;
		19'b1000000010101110101: color_data = Z;
		19'b1000000010101110110: color_data = Z;
		19'b1000000010101110111: color_data = Z;
		19'b1000000010101111000: color_data = Z;
		19'b1000000010101111001: color_data = Z;
		19'b1000000010101111010: color_data = Z;
		19'b1000000010101111011: color_data = Z;
		19'b1000000010101111100: color_data = Z;
		19'b1000000010101111101: color_data = Z;
		19'b1000000010101111110: color_data = Z;
		19'b1000000010101111111: color_data = Z;
		19'b1000000010110000000: color_data = Z;
		19'b1000000010110000001: color_data = Z;
		19'b1000000010110000010: color_data = Z;
		19'b1000000010110000011: color_data = Z;
		19'b1000000010110000100: color_data = Z;
		19'b1000000010110000101: color_data = Z;
		19'b1000000010110000110: color_data = Z;
		19'b1000000010110000111: color_data = Z;
		19'b1000000010110001000: color_data = Z;
		19'b1000000010110001001: color_data = Z;
		19'b1000000010110001010: color_data = Z;
		19'b1000000010110001011: color_data = Z;
		19'b1000000010110001100: color_data = Z;
		19'b1000000010110001101: color_data = Z;
		19'b1000000010110001110: color_data = Z;
		19'b1000000010110001111: color_data = Z;
		19'b1000000010110010000: color_data = Z;
		19'b1000000010110010001: color_data = Z;
		19'b1000000010110010010: color_data = Z;
		19'b1000000010110010011: color_data = Z;
		19'b1000000010110010100: color_data = Z;
		19'b1000000010110010101: color_data = Z;
		19'b1000000010110010110: color_data = Z;
		19'b1000000010110010111: color_data = Z;
		19'b1000000010110011000: color_data = Z;
		19'b1000000010110011001: color_data = Z;
		19'b1000000010110011010: color_data = Z;
		19'b1000000010110011011: color_data = Z;
		19'b1000000010110011100: color_data = Z;
		19'b1000000010110011101: color_data = Z;
		19'b1000000010110011110: color_data = Z;
		19'b1000000010110011111: color_data = Z;
		19'b1000000010110100000: color_data = Z;
		19'b1000000010110100001: color_data = Z;
		19'b1000000010110100010: color_data = Z;
		19'b1000000010110100011: color_data = Z;
		19'b1000000010110100100: color_data = Z;
		19'b1000000010110100101: color_data = Z;
		19'b1000000010110100110: color_data = Z;
		19'b1000000010110100111: color_data = Z;
		19'b1000000010110101000: color_data = Z;
		19'b1000000010110101001: color_data = Z;
		19'b1000000010110101010: color_data = Z;
		19'b1000000010110101011: color_data = Z;
		19'b1000000010110101100: color_data = Z;
		19'b1000000010110101101: color_data = Z;
		19'b1000000010110101110: color_data = Z;
		19'b1000000010110101111: color_data = Z;
		19'b1000000010110110000: color_data = Z;
		19'b1000000010110110001: color_data = Z;
		19'b1000000010110110010: color_data = Z;
		19'b1000000010110110011: color_data = Z;
		19'b1000000010110110100: color_data = Z;
		19'b1000000010110110101: color_data = Z;
		19'b1000000010110110110: color_data = Z;
		19'b1000000010110110111: color_data = Z;
		19'b1000000010110111000: color_data = Z;
		19'b1000000010110111001: color_data = Z;
		19'b1000000010110111010: color_data = Z;
		19'b1000000010110111011: color_data = Z;
		19'b1000000010110111100: color_data = Z;
		19'b1000000010111000001: color_data = Z;
		19'b1000000010111000010: color_data = Z;
		19'b1000000010111000011: color_data = Z;
		19'b1000000010111000100: color_data = Z;
		19'b1000000010111000101: color_data = Z;
		19'b1000000010111000110: color_data = Z;
		19'b1000000010111000111: color_data = Z;
		19'b1000000010111001000: color_data = Z;
		19'b1000000010111001001: color_data = Z;
		19'b1000000100010110101: color_data = Z;
		19'b1000000100010110110: color_data = Z;
		19'b1000000100010110111: color_data = Z;
		19'b1000000100010111000: color_data = Z;
		19'b1000000100010111001: color_data = Z;
		19'b1000000100010111010: color_data = Z;
		19'b1000000100010111011: color_data = Z;
		19'b1000000100010111100: color_data = Z;
		19'b1000000100010111101: color_data = Z;
		19'b1000000100010111110: color_data = Z;
		19'b1000000100010111111: color_data = Z;
		19'b1000000100011000000: color_data = Z;
		19'b1000000100011000001: color_data = Z;
		19'b1000000100011000010: color_data = Z;
		19'b1000000100011000011: color_data = Z;
		19'b1000000100011000100: color_data = Z;
		19'b1000000100011000101: color_data = Z;
		19'b1000000100011000110: color_data = Z;
		19'b1000000100011000111: color_data = Z;
		19'b1000000100011001000: color_data = Z;
		19'b1000000100011001001: color_data = Z;
		19'b1000000100011010000: color_data = Z;
		19'b1000000100011010001: color_data = Z;
		19'b1000000100011010010: color_data = Z;
		19'b1000000100011010011: color_data = Z;
		19'b1000000100011010100: color_data = Z;
		19'b1000000100011010101: color_data = Z;
		19'b1000000100011010110: color_data = Z;
		19'b1000000100011010111: color_data = Z;
		19'b1000000100011011000: color_data = Z;
		19'b1000000100011011001: color_data = Z;
		19'b1000000100011011010: color_data = Z;
		19'b1000000100011011011: color_data = Z;
		19'b1000000100011011100: color_data = Z;
		19'b1000000100011011101: color_data = Z;
		19'b1000000100011011110: color_data = Z;
		19'b1000000100011011111: color_data = Z;
		19'b1000000100011100000: color_data = Z;
		19'b1000000100011101011: color_data = Z;
		19'b1000000100011101100: color_data = Z;
		19'b1000000100011101101: color_data = Z;
		19'b1000000100011101110: color_data = Z;
		19'b1000000100011101111: color_data = Z;
		19'b1000000100011110000: color_data = Z;
		19'b1000000100011110001: color_data = Z;
		19'b1000000100011110010: color_data = Z;
		19'b1000000100011110011: color_data = Z;
		19'b1000000100011110100: color_data = Z;
		19'b1000000100011110101: color_data = Z;
		19'b1000000100011110110: color_data = Z;
		19'b1000000100011110111: color_data = Z;
		19'b1000000100011111000: color_data = Z;
		19'b1000000100011111001: color_data = Z;
		19'b1000000100100000110: color_data = Z;
		19'b1000000100100000111: color_data = Z;
		19'b1000000100100001000: color_data = Z;
		19'b1000000100100001001: color_data = Z;
		19'b1000000100100001010: color_data = Z;
		19'b1000000100100001011: color_data = Z;
		19'b1000000100100001100: color_data = Z;
		19'b1000000100100001101: color_data = Z;
		19'b1000000100100001110: color_data = Z;
		19'b1000000100100001111: color_data = Z;
		19'b1000000100100010000: color_data = Z;
		19'b1000000100100010001: color_data = Z;
		19'b1000000100100010010: color_data = Z;
		19'b1000000100100010011: color_data = Z;
		19'b1000000100100010100: color_data = Z;
		19'b1000000100100010101: color_data = Z;
		19'b1000000100100010110: color_data = Z;
		19'b1000000100100010111: color_data = Z;
		19'b1000000100100011000: color_data = Z;
		19'b1000000100100011001: color_data = Z;
		19'b1000000100100011010: color_data = Z;
		19'b1000000100100011011: color_data = Z;
		19'b1000000100100011100: color_data = Z;
		19'b1000000100100011101: color_data = Z;
		19'b1000000100100011110: color_data = Z;
		19'b1000000100100011111: color_data = Z;
		19'b1000000100100100000: color_data = Z;
		19'b1000000100100100001: color_data = Z;
		19'b1000000100100100010: color_data = Z;
		19'b1000000100100100011: color_data = Z;
		19'b1000000100100100100: color_data = Z;
		19'b1000000100100100101: color_data = Z;
		19'b1000000100100100110: color_data = Z;
		19'b1000000100100100111: color_data = Z;
		19'b1000000100100101000: color_data = Z;
		19'b1000000100100101001: color_data = Z;
		19'b1000000100100101010: color_data = Z;
		19'b1000000100100101011: color_data = Z;
		19'b1000000100100101100: color_data = Z;
		19'b1000000100100101101: color_data = Z;
		19'b1000000100100101110: color_data = Z;
		19'b1000000100100110111: color_data = Z;
		19'b1000000100100111000: color_data = Z;
		19'b1000000100100111001: color_data = Z;
		19'b1000000100100111010: color_data = Z;
		19'b1000000100100111011: color_data = Z;
		19'b1000000100100111100: color_data = Z;
		19'b1000000100100111101: color_data = Z;
		19'b1000000100100111110: color_data = Z;
		19'b1000000100100111111: color_data = Z;
		19'b1000000100101001000: color_data = Z;
		19'b1000000100101001001: color_data = Z;
		19'b1000000100101001010: color_data = Z;
		19'b1000000100101001011: color_data = Z;
		19'b1000000100101001100: color_data = Z;
		19'b1000000100101001101: color_data = Z;
		19'b1000000100101001110: color_data = Z;
		19'b1000000100101001111: color_data = Z;
		19'b1000000100101010000: color_data = Z;
		19'b1000000100101010001: color_data = Z;
		19'b1000000100101010010: color_data = Z;
		19'b1000000100101010011: color_data = Z;
		19'b1000000100101010100: color_data = Z;
		19'b1000000100101010101: color_data = Z;
		19'b1000000100101010110: color_data = Z;
		19'b1000000100101010111: color_data = Z;
		19'b1000000100101011110: color_data = Z;
		19'b1000000100101011111: color_data = Z;
		19'b1000000100101100000: color_data = Z;
		19'b1000000100101100001: color_data = Z;
		19'b1000000100101100010: color_data = Z;
		19'b1000000100101100011: color_data = Z;
		19'b1000000100101100100: color_data = Z;
		19'b1000000100101100101: color_data = Z;
		19'b1000000100101101010: color_data = Z;
		19'b1000000100101101011: color_data = Z;
		19'b1000000100101101100: color_data = Z;
		19'b1000000100101101101: color_data = Z;
		19'b1000000100101101110: color_data = Z;
		19'b1000000100101101111: color_data = Z;
		19'b1000000100101110000: color_data = Z;
		19'b1000000100101110001: color_data = Z;
		19'b1000000100101110010: color_data = Z;
		19'b1000000100101110011: color_data = Z;
		19'b1000000100101110100: color_data = Z;
		19'b1000000100101110101: color_data = Z;
		19'b1000000100101110110: color_data = Z;
		19'b1000000100101110111: color_data = Z;
		19'b1000000100101111000: color_data = Z;
		19'b1000000100101111001: color_data = Z;
		19'b1000000100101111010: color_data = Z;
		19'b1000000100101111011: color_data = Z;
		19'b1000000100101111100: color_data = Z;
		19'b1000000100101111101: color_data = Z;
		19'b1000000100101111110: color_data = Z;
		19'b1000000100101111111: color_data = Z;
		19'b1000000100110000000: color_data = Z;
		19'b1000000100110000001: color_data = Z;
		19'b1000000100110000010: color_data = Z;
		19'b1000000100110000011: color_data = Z;
		19'b1000000100110000100: color_data = Z;
		19'b1000000100110000101: color_data = Z;
		19'b1000000100110000110: color_data = Z;
		19'b1000000100110000111: color_data = Z;
		19'b1000000100110001000: color_data = Z;
		19'b1000000100110001001: color_data = Z;
		19'b1000000100110001010: color_data = Z;
		19'b1000000100110001011: color_data = Z;
		19'b1000000100110001100: color_data = Z;
		19'b1000000100110001101: color_data = Z;
		19'b1000000100110001110: color_data = Z;
		19'b1000000100110001111: color_data = Z;
		19'b1000000100110010000: color_data = Z;
		19'b1000000100110010100: color_data = Z;
		19'b1000000100110010101: color_data = Z;
		19'b1000000100110010110: color_data = Z;
		19'b1000000100110010111: color_data = Z;
		19'b1000000100110011000: color_data = Z;
		19'b1000000100110011001: color_data = Z;
		19'b1000000100110011010: color_data = Z;
		19'b1000000100110011011: color_data = Z;
		19'b1000000100110011100: color_data = Z;
		19'b1000000100110011101: color_data = Z;
		19'b1000000100110011110: color_data = Z;
		19'b1000000100110011111: color_data = Z;
		19'b1000000100110100000: color_data = Z;
		19'b1000000100110100001: color_data = Z;
		19'b1000000100110100010: color_data = Z;
		19'b1000000100110100011: color_data = Z;
		19'b1000000100110100100: color_data = Z;
		19'b1000000100110100101: color_data = Z;
		19'b1000000100110100110: color_data = Z;
		19'b1000000100110100111: color_data = Z;
		19'b1000000100110101000: color_data = Z;
		19'b1000000100110101001: color_data = Z;
		19'b1000000100110101010: color_data = Z;
		19'b1000000100110101011: color_data = Z;
		19'b1000000100110101100: color_data = Z;
		19'b1000000100110101101: color_data = Z;
		19'b1000000100110101110: color_data = Z;
		19'b1000000100110101111: color_data = Z;
		19'b1000000100110110000: color_data = Z;
		19'b1000000100110110001: color_data = Z;
		19'b1000000100110110010: color_data = Z;
		19'b1000000100110110011: color_data = Z;
		19'b1000000100110110100: color_data = Z;
		19'b1000000100110110101: color_data = Z;
		19'b1000000100110110110: color_data = Z;
		19'b1000000100110110111: color_data = Z;
		19'b1000000100110111000: color_data = Z;
		19'b1000000100110111001: color_data = Z;
		19'b1000000100110111010: color_data = Z;
		19'b1000000100110111011: color_data = Z;
		19'b1000000100110111100: color_data = Z;
		19'b1000000100111000001: color_data = Z;
		19'b1000000100111000010: color_data = Z;
		19'b1000000100111000011: color_data = Z;
		19'b1000000100111000100: color_data = Z;
		19'b1000000100111000101: color_data = Z;
		19'b1000000100111000110: color_data = Z;
		19'b1000000100111000111: color_data = Z;
		19'b1000000100111001000: color_data = Z;
		19'b1000000100111001001: color_data = Z;
		19'b1000000110010110110: color_data = Z;
		19'b1000000110010110111: color_data = Z;
		19'b1000000110010111000: color_data = Z;
		19'b1000000110010111001: color_data = Z;
		19'b1000000110010111010: color_data = Z;
		19'b1000000110010111011: color_data = Z;
		19'b1000000110010111100: color_data = Z;
		19'b1000000110010111101: color_data = Z;
		19'b1000000110010111110: color_data = Z;
		19'b1000000110010111111: color_data = Z;
		19'b1000000110011000000: color_data = Z;
		19'b1000000110011000001: color_data = Z;
		19'b1000000110011000010: color_data = Z;
		19'b1000000110011000011: color_data = Z;
		19'b1000000110011000100: color_data = Z;
		19'b1000000110011000101: color_data = Z;
		19'b1000000110011000110: color_data = Z;
		19'b1000000110011000111: color_data = Z;
		19'b1000000110011001000: color_data = Z;
		19'b1000000110011001001: color_data = Z;
		19'b1000000110011010001: color_data = Z;
		19'b1000000110011010010: color_data = Z;
		19'b1000000110011010011: color_data = Z;
		19'b1000000110011010100: color_data = Z;
		19'b1000000110011010101: color_data = Z;
		19'b1000000110011010110: color_data = Z;
		19'b1000000110011010111: color_data = Z;
		19'b1000000110011011000: color_data = Z;
		19'b1000000110011011001: color_data = Z;
		19'b1000000110011011010: color_data = Z;
		19'b1000000110011011011: color_data = Z;
		19'b1000000110011011100: color_data = Z;
		19'b1000000110011011101: color_data = Z;
		19'b1000000110011011110: color_data = Z;
		19'b1000000110011011111: color_data = Z;
		19'b1000000110011100000: color_data = Z;
		19'b1000000110011101011: color_data = Z;
		19'b1000000110011101100: color_data = Z;
		19'b1000000110011101101: color_data = Z;
		19'b1000000110011101110: color_data = Z;
		19'b1000000110011101111: color_data = Z;
		19'b1000000110011110000: color_data = Z;
		19'b1000000110011110001: color_data = Z;
		19'b1000000110011110010: color_data = Z;
		19'b1000000110011110011: color_data = Z;
		19'b1000000110011110100: color_data = Z;
		19'b1000000110011110101: color_data = Z;
		19'b1000000110011110110: color_data = Z;
		19'b1000000110011110111: color_data = Z;
		19'b1000000110011111000: color_data = Z;
		19'b1000000110100000101: color_data = Z;
		19'b1000000110100000110: color_data = Z;
		19'b1000000110100000111: color_data = Z;
		19'b1000000110100001000: color_data = Z;
		19'b1000000110100001001: color_data = Z;
		19'b1000000110100001010: color_data = Z;
		19'b1000000110100001011: color_data = Z;
		19'b1000000110100001100: color_data = Z;
		19'b1000000110100001101: color_data = Z;
		19'b1000000110100001110: color_data = Z;
		19'b1000000110100001111: color_data = Z;
		19'b1000000110100010000: color_data = Z;
		19'b1000000110100010001: color_data = Z;
		19'b1000000110100010010: color_data = Z;
		19'b1000000110100010011: color_data = Z;
		19'b1000000110100010100: color_data = Z;
		19'b1000000110100010101: color_data = Z;
		19'b1000000110100010110: color_data = Z;
		19'b1000000110100010111: color_data = Z;
		19'b1000000110100011000: color_data = Z;
		19'b1000000110100011001: color_data = Z;
		19'b1000000110100011010: color_data = Z;
		19'b1000000110100011011: color_data = Z;
		19'b1000000110100011100: color_data = Z;
		19'b1000000110100011101: color_data = Z;
		19'b1000000110100011110: color_data = Z;
		19'b1000000110100011111: color_data = Z;
		19'b1000000110100100000: color_data = Z;
		19'b1000000110100100001: color_data = Z;
		19'b1000000110100100010: color_data = Z;
		19'b1000000110100100011: color_data = Z;
		19'b1000000110100100100: color_data = Z;
		19'b1000000110100100101: color_data = Z;
		19'b1000000110100100110: color_data = Z;
		19'b1000000110100100111: color_data = Z;
		19'b1000000110100101000: color_data = Z;
		19'b1000000110100101001: color_data = Z;
		19'b1000000110100101010: color_data = Z;
		19'b1000000110100101011: color_data = Z;
		19'b1000000110100101100: color_data = Z;
		19'b1000000110100101101: color_data = Z;
		19'b1000000110100101110: color_data = Z;
		19'b1000000110100110111: color_data = Z;
		19'b1000000110100111000: color_data = Z;
		19'b1000000110100111001: color_data = Z;
		19'b1000000110100111010: color_data = Z;
		19'b1000000110100111011: color_data = Z;
		19'b1000000110100111100: color_data = Z;
		19'b1000000110100111101: color_data = Z;
		19'b1000000110101001001: color_data = Z;
		19'b1000000110101001010: color_data = Z;
		19'b1000000110101001011: color_data = Z;
		19'b1000000110101001100: color_data = Z;
		19'b1000000110101001101: color_data = Z;
		19'b1000000110101001110: color_data = Z;
		19'b1000000110101001111: color_data = Z;
		19'b1000000110101010000: color_data = Z;
		19'b1000000110101010001: color_data = Z;
		19'b1000000110101010010: color_data = Z;
		19'b1000000110101010011: color_data = Z;
		19'b1000000110101010100: color_data = Z;
		19'b1000000110101010101: color_data = Z;
		19'b1000000110101010110: color_data = Z;
		19'b1000000110101010111: color_data = Z;
		19'b1000000110101100000: color_data = Z;
		19'b1000000110101100001: color_data = Z;
		19'b1000000110101100010: color_data = Z;
		19'b1000000110101100011: color_data = Z;
		19'b1000000110101100100: color_data = Z;
		19'b1000000110101100101: color_data = Z;
		19'b1000000110101101010: color_data = Z;
		19'b1000000110101101011: color_data = Z;
		19'b1000000110101101100: color_data = Z;
		19'b1000000110101101101: color_data = Z;
		19'b1000000110101101110: color_data = Z;
		19'b1000000110101101111: color_data = Z;
		19'b1000000110101110000: color_data = Z;
		19'b1000000110101110001: color_data = Z;
		19'b1000000110101110010: color_data = Z;
		19'b1000000110101110011: color_data = Z;
		19'b1000000110101110100: color_data = Z;
		19'b1000000110101110101: color_data = Z;
		19'b1000000110101110110: color_data = Z;
		19'b1000000110101110111: color_data = Z;
		19'b1000000110101111000: color_data = Z;
		19'b1000000110101111001: color_data = Z;
		19'b1000000110101111010: color_data = Z;
		19'b1000000110101111011: color_data = Z;
		19'b1000000110101111100: color_data = Z;
		19'b1000000110101111101: color_data = Z;
		19'b1000000110101111110: color_data = Z;
		19'b1000000110101111111: color_data = Z;
		19'b1000000110110000000: color_data = Z;
		19'b1000000110110000001: color_data = Z;
		19'b1000000110110000010: color_data = Z;
		19'b1000000110110000011: color_data = Z;
		19'b1000000110110000100: color_data = Z;
		19'b1000000110110000101: color_data = Z;
		19'b1000000110110000110: color_data = Z;
		19'b1000000110110000111: color_data = Z;
		19'b1000000110110001000: color_data = Z;
		19'b1000000110110001001: color_data = Z;
		19'b1000000110110001010: color_data = Z;
		19'b1000000110110001011: color_data = Z;
		19'b1000000110110001100: color_data = Z;
		19'b1000000110110001101: color_data = Z;
		19'b1000000110110001110: color_data = Z;
		19'b1000000110110001111: color_data = Z;
		19'b1000000110110010000: color_data = Z;
		19'b1000000110110010001: color_data = Z;
		19'b1000000110110010010: color_data = Z;
		19'b1000000110110010110: color_data = Z;
		19'b1000000110110010111: color_data = Z;
		19'b1000000110110011000: color_data = Z;
		19'b1000000110110011001: color_data = Z;
		19'b1000000110110011010: color_data = Z;
		19'b1000000110110011011: color_data = Z;
		19'b1000000110110011100: color_data = Z;
		19'b1000000110110011101: color_data = Z;
		19'b1000000110110011110: color_data = Z;
		19'b1000000110110011111: color_data = Z;
		19'b1000000110110100000: color_data = Z;
		19'b1000000110110100001: color_data = Z;
		19'b1000000110110100010: color_data = Z;
		19'b1000000110110100011: color_data = Z;
		19'b1000000110110100100: color_data = Z;
		19'b1000000110110100101: color_data = Z;
		19'b1000000110110100110: color_data = Z;
		19'b1000000110110100111: color_data = Z;
		19'b1000000110110101000: color_data = Z;
		19'b1000000110110101001: color_data = Z;
		19'b1000000110110101010: color_data = Z;
		19'b1000000110110101011: color_data = Z;
		19'b1000000110110101100: color_data = Z;
		19'b1000000110110101101: color_data = Z;
		19'b1000000110110101110: color_data = Z;
		19'b1000000110110101111: color_data = Z;
		19'b1000000110110110000: color_data = Z;
		19'b1000000110110110001: color_data = Z;
		19'b1000000110110110010: color_data = Z;
		19'b1000000110110110011: color_data = Z;
		19'b1000000110110110100: color_data = Z;
		19'b1000000110110110101: color_data = Z;
		19'b1000000110110110110: color_data = Z;
		19'b1000000110110110111: color_data = Z;
		19'b1000000110110111000: color_data = Z;
		19'b1000000110110111001: color_data = Z;
		19'b1000000110110111010: color_data = Z;
		19'b1000000110110111011: color_data = Z;
		19'b1000000110110111100: color_data = Z;
		19'b1000000110111000001: color_data = Z;
		19'b1000000110111000010: color_data = Z;
		19'b1000000110111000011: color_data = Z;
		19'b1000000110111000100: color_data = Z;
		19'b1000000110111000101: color_data = Z;
		19'b1000000110111000110: color_data = Z;
		19'b1000000110111000111: color_data = Z;
		19'b1000000110111001000: color_data = Z;
		19'b1000000110111001001: color_data = Z;
		19'b1000000110111001010: color_data = Z;
		19'b1000001000010110111: color_data = Z;
		19'b1000001000010111000: color_data = Z;
		19'b1000001000010111001: color_data = Z;
		19'b1000001000010111010: color_data = Z;
		19'b1000001000010111011: color_data = Z;
		19'b1000001000010111100: color_data = Z;
		19'b1000001000010111101: color_data = Z;
		19'b1000001000010111110: color_data = Z;
		19'b1000001000010111111: color_data = Z;
		19'b1000001000011000000: color_data = Z;
		19'b1000001000011000001: color_data = Z;
		19'b1000001000011000010: color_data = Z;
		19'b1000001000011000011: color_data = Z;
		19'b1000001000011000100: color_data = Z;
		19'b1000001000011000101: color_data = Z;
		19'b1000001000011000110: color_data = Z;
		19'b1000001000011000111: color_data = Z;
		19'b1000001000011001000: color_data = Z;
		19'b1000001000011001001: color_data = Z;
		19'b1000001000011001010: color_data = Z;
		19'b1000001000011010001: color_data = Z;
		19'b1000001000011010010: color_data = Z;
		19'b1000001000011010011: color_data = Z;
		19'b1000001000011010100: color_data = Z;
		19'b1000001000011010101: color_data = Z;
		19'b1000001000011010110: color_data = Z;
		19'b1000001000011010111: color_data = Z;
		19'b1000001000011011000: color_data = Z;
		19'b1000001000011011001: color_data = Z;
		19'b1000001000011011010: color_data = Z;
		19'b1000001000011011011: color_data = Z;
		19'b1000001000011011100: color_data = Z;
		19'b1000001000011011101: color_data = Z;
		19'b1000001000011011110: color_data = Z;
		19'b1000001000011011111: color_data = Z;
		19'b1000001000011100000: color_data = Z;
		19'b1000001000011101100: color_data = Z;
		19'b1000001000011101101: color_data = Z;
		19'b1000001000011101110: color_data = Z;
		19'b1000001000011101111: color_data = Z;
		19'b1000001000011110000: color_data = Z;
		19'b1000001000011110001: color_data = Z;
		19'b1000001000011110010: color_data = Z;
		19'b1000001000011110011: color_data = Z;
		19'b1000001000011110100: color_data = Z;
		19'b1000001000011110101: color_data = Z;
		19'b1000001000011110110: color_data = Z;
		19'b1000001000100000011: color_data = Z;
		19'b1000001000100000100: color_data = Z;
		19'b1000001000100000101: color_data = Z;
		19'b1000001000100000110: color_data = Z;
		19'b1000001000100000111: color_data = Z;
		19'b1000001000100001000: color_data = Z;
		19'b1000001000100001001: color_data = Z;
		19'b1000001000100001010: color_data = Z;
		19'b1000001000100001011: color_data = Z;
		19'b1000001000100001100: color_data = Z;
		19'b1000001000100001101: color_data = Z;
		19'b1000001000100001110: color_data = Z;
		19'b1000001000100001111: color_data = Z;
		19'b1000001000100010000: color_data = Z;
		19'b1000001000100010001: color_data = Z;
		19'b1000001000100010010: color_data = Z;
		19'b1000001000100010011: color_data = Z;
		19'b1000001000100010100: color_data = Z;
		19'b1000001000100010101: color_data = Z;
		19'b1000001000100010110: color_data = Z;
		19'b1000001000100010111: color_data = Z;
		19'b1000001000100011000: color_data = Z;
		19'b1000001000100011001: color_data = Z;
		19'b1000001000100011010: color_data = Z;
		19'b1000001000100011011: color_data = Z;
		19'b1000001000100011100: color_data = Z;
		19'b1000001000100011101: color_data = Z;
		19'b1000001000100011110: color_data = Z;
		19'b1000001000100011111: color_data = Z;
		19'b1000001000100100000: color_data = Z;
		19'b1000001000100100001: color_data = Z;
		19'b1000001000100100010: color_data = Z;
		19'b1000001000100100011: color_data = Z;
		19'b1000001000100100100: color_data = Z;
		19'b1000001000100100101: color_data = Z;
		19'b1000001000100100110: color_data = Z;
		19'b1000001000100100111: color_data = Z;
		19'b1000001000100101000: color_data = Z;
		19'b1000001000100101001: color_data = Z;
		19'b1000001000100101010: color_data = Z;
		19'b1000001000100101011: color_data = Z;
		19'b1000001000100101100: color_data = Z;
		19'b1000001000100101101: color_data = Z;
		19'b1000001000100101110: color_data = Z;
		19'b1000001000100101111: color_data = Z;
		19'b1000001000100110111: color_data = Z;
		19'b1000001000100111000: color_data = Z;
		19'b1000001000100111001: color_data = Z;
		19'b1000001000100111010: color_data = Z;
		19'b1000001000100111011: color_data = Z;
		19'b1000001000101001011: color_data = Z;
		19'b1000001000101001100: color_data = Z;
		19'b1000001000101001101: color_data = Z;
		19'b1000001000101001110: color_data = Z;
		19'b1000001000101001111: color_data = Z;
		19'b1000001000101010000: color_data = Z;
		19'b1000001000101010001: color_data = Z;
		19'b1000001000101010010: color_data = Z;
		19'b1000001000101010011: color_data = Z;
		19'b1000001000101010100: color_data = Z;
		19'b1000001000101010101: color_data = Z;
		19'b1000001000101010110: color_data = Z;
		19'b1000001000101010111: color_data = Z;
		19'b1000001000101100011: color_data = Z;
		19'b1000001000101100100: color_data = Z;
		19'b1000001000101101010: color_data = Z;
		19'b1000001000101101011: color_data = Z;
		19'b1000001000101101100: color_data = Z;
		19'b1000001000101101101: color_data = Z;
		19'b1000001000101101110: color_data = Z;
		19'b1000001000101101111: color_data = Z;
		19'b1000001000101110000: color_data = Z;
		19'b1000001000101110001: color_data = Z;
		19'b1000001000101110010: color_data = Z;
		19'b1000001000101110011: color_data = Z;
		19'b1000001000101110100: color_data = Z;
		19'b1000001000101110101: color_data = Z;
		19'b1000001000101110110: color_data = Z;
		19'b1000001000101110111: color_data = Z;
		19'b1000001000101111000: color_data = Z;
		19'b1000001000101111001: color_data = Z;
		19'b1000001000101111010: color_data = Z;
		19'b1000001000101111011: color_data = Z;
		19'b1000001000101111100: color_data = Z;
		19'b1000001000101111101: color_data = Z;
		19'b1000001000101111110: color_data = Z;
		19'b1000001000101111111: color_data = Z;
		19'b1000001000110000000: color_data = Z;
		19'b1000001000110000001: color_data = Z;
		19'b1000001000110000010: color_data = Z;
		19'b1000001000110000011: color_data = Z;
		19'b1000001000110000100: color_data = Z;
		19'b1000001000110000101: color_data = Z;
		19'b1000001000110000110: color_data = Z;
		19'b1000001000110000111: color_data = Z;
		19'b1000001000110001000: color_data = Z;
		19'b1000001000110001001: color_data = Z;
		19'b1000001000110001010: color_data = Z;
		19'b1000001000110001011: color_data = Z;
		19'b1000001000110001100: color_data = Z;
		19'b1000001000110001101: color_data = Z;
		19'b1000001000110001110: color_data = Z;
		19'b1000001000110001111: color_data = Z;
		19'b1000001000110010000: color_data = Z;
		19'b1000001000110010001: color_data = Z;
		19'b1000001000110010010: color_data = Z;
		19'b1000001000110010011: color_data = Z;
		19'b1000001000110010100: color_data = Z;
		19'b1000001000110010101: color_data = Z;
		19'b1000001000110010111: color_data = Z;
		19'b1000001000110011001: color_data = Z;
		19'b1000001000110011010: color_data = Z;
		19'b1000001000110011011: color_data = Z;
		19'b1000001000110011101: color_data = Z;
		19'b1000001000110011110: color_data = Z;
		19'b1000001000110011111: color_data = Z;
		19'b1000001000110100000: color_data = Z;
		19'b1000001000110100001: color_data = Z;
		19'b1000001000110100010: color_data = Z;
		19'b1000001000110100011: color_data = Z;
		19'b1000001000110100100: color_data = Z;
		19'b1000001000110100101: color_data = Z;
		19'b1000001000110100110: color_data = Z;
		19'b1000001000110100111: color_data = Z;
		19'b1000001000110101000: color_data = Z;
		19'b1000001000110101001: color_data = Z;
		19'b1000001000110101010: color_data = Z;
		19'b1000001000110101011: color_data = Z;
		19'b1000001000110101100: color_data = Z;
		19'b1000001000110101101: color_data = Z;
		19'b1000001000110101110: color_data = Z;
		19'b1000001000110101111: color_data = Z;
		19'b1000001000110110000: color_data = Z;
		19'b1000001000110110001: color_data = Z;
		19'b1000001000110110010: color_data = Z;
		19'b1000001000110110011: color_data = Z;
		19'b1000001000110110100: color_data = Z;
		19'b1000001000110110101: color_data = Z;
		19'b1000001000110110110: color_data = Z;
		19'b1000001000110110111: color_data = Z;
		19'b1000001000110111000: color_data = Z;
		19'b1000001000110111001: color_data = Z;
		19'b1000001000110111010: color_data = Z;
		19'b1000001000110111011: color_data = Z;
		19'b1000001000110111100: color_data = Z;
		19'b1000001000111000001: color_data = Z;
		19'b1000001000111000010: color_data = Z;
		19'b1000001000111000011: color_data = Z;
		19'b1000001000111000100: color_data = Z;
		19'b1000001000111000101: color_data = Z;
		19'b1000001000111000110: color_data = Z;
		19'b1000001000111000111: color_data = Z;
		19'b1000001000111001000: color_data = Z;
		19'b1000001000111001001: color_data = Z;
		19'b1000001000111001010: color_data = Z;
		19'b1000001010010110111: color_data = Z;
		19'b1000001010010111000: color_data = Z;
		19'b1000001010010111001: color_data = Z;
		19'b1000001010010111010: color_data = Z;
		19'b1000001010010111011: color_data = Z;
		19'b1000001010010111100: color_data = Z;
		19'b1000001010010111101: color_data = Z;
		19'b1000001010010111110: color_data = Z;
		19'b1000001010010111111: color_data = Z;
		19'b1000001010011000000: color_data = Z;
		19'b1000001010011000001: color_data = Z;
		19'b1000001010011000010: color_data = Z;
		19'b1000001010011000011: color_data = Z;
		19'b1000001010011000100: color_data = Z;
		19'b1000001010011000101: color_data = Z;
		19'b1000001010011000110: color_data = Z;
		19'b1000001010011000111: color_data = Z;
		19'b1000001010011001000: color_data = Z;
		19'b1000001010011001001: color_data = Z;
		19'b1000001010011001010: color_data = Z;
		19'b1000001010011001011: color_data = Z;
		19'b1000001010011010011: color_data = Z;
		19'b1000001010011010100: color_data = Z;
		19'b1000001010011010101: color_data = Z;
		19'b1000001010011010110: color_data = Z;
		19'b1000001010011010111: color_data = Z;
		19'b1000001010011011000: color_data = Z;
		19'b1000001010011011001: color_data = Z;
		19'b1000001010011011010: color_data = Z;
		19'b1000001010011011011: color_data = Z;
		19'b1000001010011011100: color_data = Z;
		19'b1000001010011011101: color_data = Z;
		19'b1000001010011011110: color_data = Z;
		19'b1000001010011011111: color_data = Z;
		19'b1000001010011101101: color_data = Z;
		19'b1000001010011101110: color_data = Z;
		19'b1000001010011101111: color_data = Z;
		19'b1000001010011110000: color_data = Z;
		19'b1000001010011110001: color_data = Z;
		19'b1000001010011110010: color_data = Z;
		19'b1000001010011110011: color_data = Z;
		19'b1000001010011110100: color_data = Z;
		19'b1000001010100000010: color_data = Z;
		19'b1000001010100000011: color_data = Z;
		19'b1000001010100000100: color_data = Z;
		19'b1000001010100000101: color_data = Z;
		19'b1000001010100000110: color_data = Z;
		19'b1000001010100000111: color_data = Z;
		19'b1000001010100001000: color_data = Z;
		19'b1000001010100001001: color_data = Z;
		19'b1000001010100001010: color_data = Z;
		19'b1000001010100001011: color_data = Z;
		19'b1000001010100001100: color_data = Z;
		19'b1000001010100001101: color_data = Z;
		19'b1000001010100001110: color_data = Z;
		19'b1000001010100001111: color_data = Z;
		19'b1000001010100010000: color_data = Z;
		19'b1000001010100010001: color_data = Z;
		19'b1000001010100010010: color_data = Z;
		19'b1000001010100010011: color_data = Z;
		19'b1000001010100010100: color_data = Z;
		19'b1000001010100010101: color_data = Z;
		19'b1000001010100010110: color_data = Z;
		19'b1000001010100010111: color_data = Z;
		19'b1000001010100011000: color_data = Z;
		19'b1000001010100011001: color_data = Z;
		19'b1000001010100011010: color_data = Z;
		19'b1000001010100011011: color_data = Z;
		19'b1000001010100011100: color_data = Z;
		19'b1000001010100011101: color_data = Z;
		19'b1000001010100011110: color_data = Z;
		19'b1000001010100011111: color_data = Z;
		19'b1000001010100100000: color_data = Z;
		19'b1000001010100100001: color_data = Z;
		19'b1000001010100100010: color_data = Z;
		19'b1000001010100100011: color_data = Z;
		19'b1000001010100100100: color_data = Z;
		19'b1000001010100100101: color_data = Z;
		19'b1000001010100100110: color_data = Z;
		19'b1000001010100100111: color_data = Z;
		19'b1000001010100101000: color_data = Z;
		19'b1000001010100101001: color_data = Z;
		19'b1000001010100101010: color_data = Z;
		19'b1000001010100101011: color_data = Z;
		19'b1000001010100101100: color_data = Z;
		19'b1000001010100101101: color_data = Z;
		19'b1000001010100101110: color_data = Z;
		19'b1000001010100101111: color_data = Z;
		19'b1000001010100111000: color_data = Z;
		19'b1000001010100111001: color_data = Z;
		19'b1000001010100111010: color_data = Z;
		19'b1000001010101001110: color_data = Z;
		19'b1000001010101001111: color_data = Z;
		19'b1000001010101010000: color_data = Z;
		19'b1000001010101010001: color_data = Z;
		19'b1000001010101010010: color_data = Z;
		19'b1000001010101010011: color_data = Z;
		19'b1000001010101010100: color_data = Z;
		19'b1000001010101010101: color_data = Z;
		19'b1000001010101010110: color_data = Z;
		19'b1000001010101010111: color_data = Z;
		19'b1000001010101101010: color_data = Z;
		19'b1000001010101101011: color_data = Z;
		19'b1000001010101101100: color_data = Z;
		19'b1000001010101101101: color_data = Z;
		19'b1000001010101101110: color_data = Z;
		19'b1000001010101101111: color_data = Z;
		19'b1000001010101110000: color_data = Z;
		19'b1000001010101110001: color_data = Z;
		19'b1000001010101110010: color_data = Z;
		19'b1000001010101110011: color_data = Z;
		19'b1000001010101110100: color_data = Z;
		19'b1000001010101110101: color_data = Z;
		19'b1000001010101110110: color_data = Z;
		19'b1000001010101110111: color_data = Z;
		19'b1000001010101111000: color_data = Z;
		19'b1000001010101111001: color_data = Z;
		19'b1000001010101111010: color_data = Z;
		19'b1000001010101111011: color_data = Z;
		19'b1000001010101111100: color_data = Z;
		19'b1000001010101111101: color_data = Z;
		19'b1000001010101111110: color_data = Z;
		19'b1000001010101111111: color_data = Z;
		19'b1000001010110000000: color_data = Z;
		19'b1000001010110000001: color_data = Z;
		19'b1000001010110000010: color_data = Z;
		19'b1000001010110000011: color_data = Z;
		19'b1000001010110000100: color_data = Z;
		19'b1000001010110000101: color_data = Z;
		19'b1000001010110000110: color_data = Z;
		19'b1000001010110000111: color_data = Z;
		19'b1000001010110001000: color_data = Z;
		19'b1000001010110001001: color_data = Z;
		19'b1000001010110001010: color_data = Z;
		19'b1000001010110001011: color_data = Z;
		19'b1000001010110001100: color_data = Z;
		19'b1000001010110001101: color_data = Z;
		19'b1000001010110001110: color_data = Z;
		19'b1000001010110001111: color_data = Z;
		19'b1000001010110010000: color_data = Z;
		19'b1000001010110010001: color_data = Z;
		19'b1000001010110010010: color_data = Z;
		19'b1000001010110010011: color_data = Z;
		19'b1000001010110010100: color_data = Z;
		19'b1000001010110010101: color_data = Z;
		19'b1000001010110010110: color_data = Z;
		19'b1000001010110010111: color_data = Z;
		19'b1000001010110011000: color_data = Z;
		19'b1000001010110011001: color_data = Z;
		19'b1000001010110011010: color_data = Z;
		19'b1000001010110011011: color_data = Z;
		19'b1000001010110011101: color_data = Z;
		19'b1000001010110011110: color_data = Z;
		19'b1000001010110011111: color_data = Z;
		19'b1000001010110100000: color_data = Z;
		19'b1000001010110100001: color_data = Z;
		19'b1000001010110100010: color_data = Z;
		19'b1000001010110100011: color_data = Z;
		19'b1000001010110100100: color_data = Z;
		19'b1000001010110100101: color_data = Z;
		19'b1000001010110100110: color_data = Z;
		19'b1000001010110100111: color_data = Z;
		19'b1000001010110101000: color_data = Z;
		19'b1000001010110101001: color_data = Z;
		19'b1000001010110101010: color_data = Z;
		19'b1000001010110101011: color_data = Z;
		19'b1000001010110101100: color_data = Z;
		19'b1000001010110101101: color_data = Z;
		19'b1000001010110101110: color_data = Z;
		19'b1000001010110101111: color_data = Z;
		19'b1000001010110110000: color_data = Z;
		19'b1000001010110110001: color_data = Z;
		19'b1000001010110110010: color_data = Z;
		19'b1000001010110110011: color_data = Z;
		19'b1000001010110110100: color_data = Z;
		19'b1000001010110110101: color_data = Z;
		19'b1000001010110110110: color_data = Z;
		19'b1000001010110110111: color_data = Z;
		19'b1000001010110111000: color_data = Z;
		19'b1000001010110111001: color_data = Z;
		19'b1000001010110111010: color_data = Z;
		19'b1000001010110111011: color_data = Z;
		19'b1000001010110111100: color_data = Z;
		19'b1000001010111000001: color_data = Z;
		19'b1000001010111000010: color_data = Z;
		19'b1000001010111000011: color_data = Z;
		19'b1000001010111000100: color_data = Z;
		19'b1000001010111000101: color_data = Z;
		19'b1000001010111000110: color_data = Z;
		19'b1000001010111000111: color_data = Z;
		19'b1000001010111001000: color_data = Z;
		19'b1000001010111001001: color_data = Z;
		19'b1000001010111001010: color_data = Z;
		19'b1000001010111001011: color_data = Z;
		19'b1000001100010111000: color_data = Z;
		19'b1000001100010111001: color_data = Z;
		19'b1000001100010111010: color_data = Z;
		19'b1000001100010111011: color_data = Z;
		19'b1000001100010111100: color_data = Z;
		19'b1000001100010111101: color_data = Z;
		19'b1000001100010111110: color_data = Z;
		19'b1000001100010111111: color_data = Z;
		19'b1000001100011000000: color_data = Z;
		19'b1000001100011000001: color_data = Z;
		19'b1000001100011000010: color_data = Z;
		19'b1000001100011000011: color_data = Z;
		19'b1000001100011000100: color_data = Z;
		19'b1000001100011000101: color_data = Z;
		19'b1000001100011000110: color_data = Z;
		19'b1000001100011000111: color_data = Z;
		19'b1000001100011001000: color_data = Z;
		19'b1000001100011001001: color_data = Z;
		19'b1000001100011001010: color_data = Z;
		19'b1000001100011001011: color_data = Z;
		19'b1000001100011001100: color_data = Z;
		19'b1000001100011010100: color_data = Z;
		19'b1000001100011010101: color_data = Z;
		19'b1000001100011010110: color_data = Z;
		19'b1000001100011010111: color_data = Z;
		19'b1000001100011011000: color_data = Z;
		19'b1000001100011101110: color_data = Z;
		19'b1000001100011101111: color_data = Z;
		19'b1000001100011110000: color_data = Z;
		19'b1000001100011110001: color_data = Z;
		19'b1000001100011110010: color_data = Z;
		19'b1000001100011110011: color_data = Z;
		19'b1000001100100000001: color_data = Z;
		19'b1000001100100000010: color_data = Z;
		19'b1000001100100000011: color_data = Z;
		19'b1000001100100000100: color_data = Z;
		19'b1000001100100000101: color_data = Z;
		19'b1000001100100000110: color_data = Z;
		19'b1000001100100000111: color_data = Z;
		19'b1000001100100001000: color_data = Z;
		19'b1000001100100001001: color_data = Z;
		19'b1000001100100001010: color_data = Z;
		19'b1000001100100001011: color_data = Z;
		19'b1000001100100001100: color_data = Z;
		19'b1000001100100001101: color_data = Z;
		19'b1000001100100001110: color_data = Z;
		19'b1000001100100001111: color_data = Z;
		19'b1000001100100010000: color_data = Z;
		19'b1000001100100010001: color_data = Z;
		19'b1000001100100010010: color_data = Z;
		19'b1000001100100010011: color_data = Z;
		19'b1000001100100010100: color_data = Z;
		19'b1000001100100010101: color_data = Z;
		19'b1000001100100010110: color_data = Z;
		19'b1000001100100010111: color_data = Z;
		19'b1000001100100011000: color_data = Z;
		19'b1000001100100011001: color_data = Z;
		19'b1000001100100011010: color_data = Z;
		19'b1000001100100011011: color_data = Z;
		19'b1000001100100011100: color_data = Z;
		19'b1000001100100011101: color_data = Z;
		19'b1000001100100011110: color_data = Z;
		19'b1000001100100011111: color_data = Z;
		19'b1000001100100100000: color_data = Z;
		19'b1000001100100100001: color_data = Z;
		19'b1000001100100100010: color_data = Z;
		19'b1000001100100100011: color_data = Z;
		19'b1000001100100100100: color_data = Z;
		19'b1000001100100100101: color_data = Z;
		19'b1000001100100100110: color_data = Z;
		19'b1000001100100100111: color_data = Z;
		19'b1000001100100101000: color_data = Z;
		19'b1000001100100101001: color_data = Z;
		19'b1000001100100101010: color_data = Z;
		19'b1000001100100101011: color_data = Z;
		19'b1000001100100101100: color_data = Z;
		19'b1000001100100101101: color_data = Z;
		19'b1000001100100101110: color_data = Z;
		19'b1000001100100111000: color_data = Z;
		19'b1000001100100111001: color_data = Z;
		19'b1000001100101010000: color_data = Z;
		19'b1000001100101010001: color_data = Z;
		19'b1000001100101010010: color_data = Z;
		19'b1000001100101010011: color_data = Z;
		19'b1000001100101010100: color_data = Z;
		19'b1000001100101010101: color_data = Z;
		19'b1000001100101010110: color_data = Z;
		19'b1000001100101010111: color_data = Z;
		19'b1000001100101101010: color_data = Z;
		19'b1000001100101101011: color_data = Z;
		19'b1000001100101101100: color_data = Z;
		19'b1000001100101101101: color_data = Z;
		19'b1000001100101101110: color_data = Z;
		19'b1000001100101101111: color_data = Z;
		19'b1000001100101110000: color_data = Z;
		19'b1000001100101110001: color_data = Z;
		19'b1000001100101110010: color_data = Z;
		19'b1000001100101110011: color_data = Z;
		19'b1000001100101110100: color_data = Z;
		19'b1000001100101110101: color_data = Z;
		19'b1000001100101110110: color_data = Z;
		19'b1000001100101110111: color_data = Z;
		19'b1000001100101111000: color_data = Z;
		19'b1000001100101111001: color_data = Z;
		19'b1000001100101111010: color_data = Z;
		19'b1000001100101111011: color_data = Z;
		19'b1000001100101111100: color_data = Z;
		19'b1000001100101111101: color_data = Z;
		19'b1000001100101111110: color_data = Z;
		19'b1000001100101111111: color_data = Z;
		19'b1000001100110000000: color_data = Z;
		19'b1000001100110000001: color_data = Z;
		19'b1000001100110000010: color_data = Z;
		19'b1000001100110000011: color_data = Z;
		19'b1000001100110000100: color_data = Z;
		19'b1000001100110000101: color_data = Z;
		19'b1000001100110000110: color_data = Z;
		19'b1000001100110000111: color_data = Z;
		19'b1000001100110001000: color_data = Z;
		19'b1000001100110001001: color_data = Z;
		19'b1000001100110001010: color_data = Z;
		19'b1000001100110001011: color_data = Z;
		19'b1000001100110001100: color_data = Z;
		19'b1000001100110001101: color_data = Z;
		19'b1000001100110001110: color_data = Z;
		19'b1000001100110001111: color_data = Z;
		19'b1000001100110010000: color_data = Z;
		19'b1000001100110010001: color_data = Z;
		19'b1000001100110010010: color_data = Z;
		19'b1000001100110010011: color_data = Z;
		19'b1000001100110010100: color_data = Z;
		19'b1000001100110010101: color_data = Z;
		19'b1000001100110010110: color_data = Z;
		19'b1000001100110010111: color_data = Z;
		19'b1000001100110011000: color_data = Z;
		19'b1000001100110011001: color_data = Z;
		19'b1000001100110011010: color_data = Z;
		19'b1000001100110011011: color_data = Z;
		19'b1000001100110011100: color_data = Z;
		19'b1000001100110011101: color_data = Z;
		19'b1000001100110011110: color_data = Z;
		19'b1000001100110011111: color_data = Z;
		19'b1000001100110100000: color_data = Z;
		19'b1000001100110100001: color_data = Z;
		19'b1000001100110100010: color_data = Z;
		19'b1000001100110100011: color_data = Z;
		19'b1000001100110100100: color_data = Z;
		19'b1000001100110100101: color_data = Z;
		19'b1000001100110100110: color_data = Z;
		19'b1000001100110100111: color_data = Z;
		19'b1000001100110101000: color_data = Z;
		19'b1000001100110101001: color_data = Z;
		19'b1000001100110101010: color_data = Z;
		19'b1000001100110101011: color_data = Z;
		19'b1000001100110101100: color_data = Z;
		19'b1000001100110101101: color_data = Z;
		19'b1000001100110101110: color_data = Z;
		19'b1000001100110101111: color_data = Z;
		19'b1000001100110110000: color_data = Z;
		19'b1000001100110110001: color_data = Z;
		19'b1000001100110110010: color_data = Z;
		19'b1000001100110110011: color_data = Z;
		19'b1000001100110110100: color_data = Z;
		19'b1000001100110110101: color_data = Z;
		19'b1000001100110110110: color_data = Z;
		19'b1000001100110110111: color_data = Z;
		19'b1000001100110111000: color_data = Z;
		19'b1000001100110111001: color_data = Z;
		19'b1000001100110111010: color_data = Z;
		19'b1000001100110111011: color_data = Z;
		19'b1000001100110111100: color_data = Z;
		19'b1000001100110111101: color_data = Z;
		19'b1000001100111000010: color_data = Z;
		19'b1000001100111000011: color_data = Z;
		19'b1000001100111000100: color_data = Z;
		19'b1000001100111000101: color_data = Z;
		19'b1000001100111000110: color_data = Z;
		19'b1000001100111000111: color_data = Z;
		19'b1000001100111001000: color_data = Z;
		19'b1000001100111001001: color_data = Z;
		19'b1000001100111001010: color_data = Z;
		19'b1000001100111001011: color_data = Z;
		19'b1000001110010111001: color_data = Z;
		19'b1000001110010111010: color_data = Z;
		19'b1000001110010111011: color_data = Z;
		19'b1000001110010111100: color_data = Z;
		19'b1000001110010111101: color_data = Z;
		19'b1000001110010111110: color_data = Z;
		19'b1000001110010111111: color_data = Z;
		19'b1000001110011000000: color_data = Z;
		19'b1000001110011000001: color_data = Z;
		19'b1000001110011000010: color_data = Z;
		19'b1000001110011000011: color_data = Z;
		19'b1000001110011000100: color_data = Z;
		19'b1000001110011000101: color_data = Z;
		19'b1000001110011000110: color_data = Z;
		19'b1000001110011000111: color_data = Z;
		19'b1000001110011001000: color_data = Z;
		19'b1000001110011001001: color_data = Z;
		19'b1000001110011001010: color_data = Z;
		19'b1000001110011001011: color_data = Z;
		19'b1000001110011001100: color_data = Z;
		19'b1000001110011001101: color_data = Z;
		19'b1000001110011101111: color_data = Z;
		19'b1000001110100000000: color_data = Z;
		19'b1000001110100000001: color_data = Z;
		19'b1000001110100000010: color_data = Z;
		19'b1000001110100000011: color_data = Z;
		19'b1000001110100000100: color_data = Z;
		19'b1000001110100000101: color_data = Z;
		19'b1000001110100000110: color_data = Z;
		19'b1000001110100000111: color_data = Z;
		19'b1000001110100001000: color_data = Z;
		19'b1000001110100001001: color_data = Z;
		19'b1000001110100001010: color_data = Z;
		19'b1000001110100001011: color_data = Z;
		19'b1000001110100001100: color_data = Z;
		19'b1000001110100001101: color_data = Z;
		19'b1000001110100001110: color_data = Z;
		19'b1000001110100001111: color_data = Z;
		19'b1000001110100010000: color_data = Z;
		19'b1000001110100010001: color_data = Z;
		19'b1000001110100010010: color_data = Z;
		19'b1000001110100010011: color_data = Z;
		19'b1000001110100010100: color_data = Z;
		19'b1000001110100010101: color_data = Z;
		19'b1000001110100010110: color_data = Z;
		19'b1000001110100010111: color_data = Z;
		19'b1000001110100011000: color_data = Z;
		19'b1000001110100011001: color_data = Z;
		19'b1000001110100011010: color_data = Z;
		19'b1000001110100011011: color_data = Z;
		19'b1000001110100011100: color_data = Z;
		19'b1000001110100011101: color_data = Z;
		19'b1000001110100011110: color_data = Z;
		19'b1000001110100011111: color_data = Z;
		19'b1000001110100100000: color_data = Z;
		19'b1000001110100100001: color_data = Z;
		19'b1000001110100100010: color_data = Z;
		19'b1000001110100100011: color_data = Z;
		19'b1000001110100100100: color_data = Z;
		19'b1000001110100100101: color_data = Z;
		19'b1000001110100100110: color_data = Z;
		19'b1000001110100100111: color_data = Z;
		19'b1000001110100101000: color_data = Z;
		19'b1000001110100101001: color_data = Z;
		19'b1000001110100101010: color_data = Z;
		19'b1000001110100101011: color_data = Z;
		19'b1000001110100101100: color_data = Z;
		19'b1000001110100101101: color_data = Z;
		19'b1000001110100101110: color_data = Z;
		19'b1000001110100111000: color_data = Z;
		19'b1000001110100111001: color_data = Z;
		19'b1000001110101001110: color_data = Z;
		19'b1000001110101001111: color_data = Z;
		19'b1000001110101010000: color_data = Z;
		19'b1000001110101010001: color_data = Z;
		19'b1000001110101010010: color_data = Z;
		19'b1000001110101010011: color_data = Z;
		19'b1000001110101010100: color_data = Z;
		19'b1000001110101010101: color_data = Z;
		19'b1000001110101010110: color_data = Z;
		19'b1000001110101010111: color_data = Z;
		19'b1000001110101101010: color_data = Z;
		19'b1000001110101101011: color_data = Z;
		19'b1000001110101101100: color_data = Z;
		19'b1000001110101101101: color_data = Z;
		19'b1000001110101101110: color_data = Z;
		19'b1000001110101101111: color_data = Z;
		19'b1000001110101110000: color_data = Z;
		19'b1000001110101110001: color_data = Z;
		19'b1000001110101110010: color_data = Z;
		19'b1000001110101110011: color_data = Z;
		19'b1000001110101110100: color_data = Z;
		19'b1000001110101110101: color_data = Z;
		19'b1000001110101110110: color_data = Z;
		19'b1000001110101110111: color_data = Z;
		19'b1000001110101111000: color_data = Z;
		19'b1000001110101111001: color_data = Z;
		19'b1000001110101111010: color_data = Z;
		19'b1000001110101111011: color_data = Z;
		19'b1000001110101111100: color_data = Z;
		19'b1000001110101111101: color_data = Z;
		19'b1000001110101111110: color_data = Z;
		19'b1000001110101111111: color_data = Z;
		19'b1000001110110000000: color_data = Z;
		19'b1000001110110000001: color_data = Z;
		19'b1000001110110000010: color_data = Z;
		19'b1000001110110000011: color_data = Z;
		19'b1000001110110000100: color_data = Z;
		19'b1000001110110000101: color_data = Z;
		19'b1000001110110000110: color_data = Z;
		19'b1000001110110000111: color_data = Z;
		19'b1000001110110001000: color_data = Z;
		19'b1000001110110001001: color_data = Z;
		19'b1000001110110001010: color_data = Z;
		19'b1000001110110001011: color_data = Z;
		19'b1000001110110001100: color_data = Z;
		19'b1000001110110001101: color_data = Z;
		19'b1000001110110001110: color_data = Z;
		19'b1000001110110001111: color_data = Z;
		19'b1000001110110010000: color_data = Z;
		19'b1000001110110010001: color_data = Z;
		19'b1000001110110010010: color_data = Z;
		19'b1000001110110010011: color_data = Z;
		19'b1000001110110010100: color_data = Z;
		19'b1000001110110010101: color_data = Z;
		19'b1000001110110010110: color_data = Z;
		19'b1000001110110010111: color_data = Z;
		19'b1000001110110011000: color_data = Z;
		19'b1000001110110011001: color_data = Z;
		19'b1000001110110011010: color_data = Z;
		19'b1000001110110011011: color_data = Z;
		19'b1000001110110011100: color_data = Z;
		19'b1000001110110011101: color_data = Z;
		19'b1000001110110011110: color_data = Z;
		19'b1000001110110011111: color_data = Z;
		19'b1000001110110100000: color_data = Z;
		19'b1000001110110100001: color_data = Z;
		19'b1000001110110100010: color_data = Z;
		19'b1000001110110100011: color_data = Z;
		19'b1000001110110100100: color_data = Z;
		19'b1000001110110100101: color_data = Z;
		19'b1000001110110100110: color_data = Z;
		19'b1000001110110100111: color_data = Z;
		19'b1000001110110101000: color_data = Z;
		19'b1000001110110101001: color_data = Z;
		19'b1000001110110101010: color_data = Z;
		19'b1000001110110101011: color_data = Z;
		19'b1000001110110101100: color_data = Z;
		19'b1000001110110101101: color_data = Z;
		19'b1000001110110101110: color_data = Z;
		19'b1000001110110101111: color_data = Z;
		19'b1000001110110110000: color_data = Z;
		19'b1000001110110110001: color_data = Z;
		19'b1000001110110110010: color_data = Z;
		19'b1000001110110110011: color_data = Z;
		19'b1000001110110110100: color_data = Z;
		19'b1000001110110110101: color_data = Z;
		19'b1000001110110110110: color_data = Z;
		19'b1000001110110110111: color_data = Z;
		19'b1000001110110111000: color_data = Z;
		19'b1000001110110111001: color_data = Z;
		19'b1000001110110111010: color_data = Z;
		19'b1000001110110111011: color_data = Z;
		19'b1000001110110111100: color_data = Z;
		19'b1000001110110111101: color_data = Z;
		19'b1000001110111000010: color_data = Z;
		19'b1000001110111000011: color_data = Z;
		19'b1000001110111000100: color_data = Z;
		19'b1000001110111000101: color_data = Z;
		19'b1000001110111000110: color_data = Z;
		19'b1000001110111000111: color_data = Z;
		19'b1000001110111001000: color_data = Z;
		19'b1000001110111001001: color_data = Z;
		19'b1000001110111001010: color_data = Z;
		19'b1000001110111001011: color_data = Z;
		19'b1000001110111001100: color_data = Z;
		19'b1000010000010111001: color_data = Z;
		19'b1000010000010111010: color_data = Z;
		19'b1000010000010111011: color_data = Z;
		19'b1000010000010111100: color_data = Z;
		19'b1000010000010111101: color_data = Z;
		19'b1000010000010111110: color_data = Z;
		19'b1000010000010111111: color_data = Z;
		19'b1000010000011000000: color_data = Z;
		19'b1000010000011000001: color_data = Z;
		19'b1000010000011000010: color_data = Z;
		19'b1000010000011000011: color_data = Z;
		19'b1000010000011000100: color_data = Z;
		19'b1000010000011000101: color_data = Z;
		19'b1000010000011000110: color_data = Z;
		19'b1000010000011000111: color_data = Z;
		19'b1000010000011001000: color_data = Z;
		19'b1000010000011001001: color_data = Z;
		19'b1000010000011001010: color_data = Z;
		19'b1000010000011001011: color_data = Z;
		19'b1000010000011001100: color_data = Z;
		19'b1000010000011001101: color_data = Z;
		19'b1000010000011001110: color_data = Z;
		19'b1000010000011111110: color_data = Z;
		19'b1000010000011111111: color_data = Z;
		19'b1000010000100000000: color_data = Z;
		19'b1000010000100000001: color_data = Z;
		19'b1000010000100000010: color_data = Z;
		19'b1000010000100000011: color_data = Z;
		19'b1000010000100000100: color_data = Z;
		19'b1000010000100000101: color_data = Z;
		19'b1000010000100000110: color_data = Z;
		19'b1000010000100000111: color_data = Z;
		19'b1000010000100001000: color_data = Z;
		19'b1000010000100001001: color_data = Z;
		19'b1000010000100001010: color_data = Z;
		19'b1000010000100001011: color_data = Z;
		19'b1000010000100001100: color_data = Z;
		19'b1000010000100001101: color_data = Z;
		19'b1000010000100001110: color_data = Z;
		19'b1000010000100001111: color_data = Z;
		19'b1000010000100010000: color_data = Z;
		19'b1000010000100010001: color_data = Z;
		19'b1000010000100010010: color_data = Z;
		19'b1000010000100010011: color_data = Z;
		19'b1000010000100010100: color_data = Z;
		19'b1000010000100010101: color_data = Z;
		19'b1000010000100010110: color_data = Z;
		19'b1000010000100010111: color_data = Z;
		19'b1000010000100011000: color_data = Z;
		19'b1000010000100011001: color_data = Z;
		19'b1000010000100011010: color_data = Z;
		19'b1000010000100011011: color_data = Z;
		19'b1000010000100011100: color_data = Z;
		19'b1000010000100011101: color_data = Z;
		19'b1000010000100011110: color_data = Z;
		19'b1000010000100011111: color_data = Z;
		19'b1000010000100100000: color_data = Z;
		19'b1000010000100100001: color_data = Z;
		19'b1000010000100100010: color_data = Z;
		19'b1000010000100100011: color_data = Z;
		19'b1000010000100100100: color_data = Z;
		19'b1000010000100100101: color_data = Z;
		19'b1000010000100100110: color_data = Z;
		19'b1000010000100100111: color_data = Z;
		19'b1000010000100101000: color_data = Z;
		19'b1000010000100101001: color_data = Z;
		19'b1000010000100101010: color_data = Z;
		19'b1000010000100101011: color_data = Z;
		19'b1000010000100101100: color_data = Z;
		19'b1000010000100101101: color_data = Z;
		19'b1000010000100101110: color_data = Z;
		19'b1000010000100111001: color_data = Z;
		19'b1000010000101001110: color_data = Z;
		19'b1000010000101001111: color_data = Z;
		19'b1000010000101010000: color_data = Z;
		19'b1000010000101010001: color_data = Z;
		19'b1000010000101010010: color_data = Z;
		19'b1000010000101010011: color_data = Z;
		19'b1000010000101010100: color_data = Z;
		19'b1000010000101010101: color_data = Z;
		19'b1000010000101010110: color_data = Z;
		19'b1000010000101010111: color_data = Z;
		19'b1000010000101101010: color_data = Z;
		19'b1000010000101101011: color_data = Z;
		19'b1000010000101101100: color_data = Z;
		19'b1000010000101101101: color_data = Z;
		19'b1000010000101101110: color_data = Z;
		19'b1000010000101101111: color_data = Z;
		19'b1000010000101110000: color_data = Z;
		19'b1000010000101110001: color_data = Z;
		19'b1000010000101110010: color_data = Z;
		19'b1000010000101110011: color_data = Z;
		19'b1000010000101110100: color_data = Z;
		19'b1000010000101110101: color_data = Z;
		19'b1000010000101110110: color_data = Z;
		19'b1000010000101110111: color_data = Z;
		19'b1000010000101111000: color_data = Z;
		19'b1000010000101111001: color_data = Z;
		19'b1000010000101111010: color_data = Z;
		19'b1000010000101111011: color_data = Z;
		19'b1000010000101111100: color_data = Z;
		19'b1000010000101111101: color_data = Z;
		19'b1000010000101111110: color_data = Z;
		19'b1000010000101111111: color_data = Z;
		19'b1000010000110000000: color_data = Z;
		19'b1000010000110000001: color_data = Z;
		19'b1000010000110000010: color_data = Z;
		19'b1000010000110000011: color_data = Z;
		19'b1000010000110000100: color_data = Z;
		19'b1000010000110000101: color_data = Z;
		19'b1000010000110000110: color_data = Z;
		19'b1000010000110000111: color_data = Z;
		19'b1000010000110001000: color_data = Z;
		19'b1000010000110001001: color_data = Z;
		19'b1000010000110001010: color_data = Z;
		19'b1000010000110001011: color_data = Z;
		19'b1000010000110001100: color_data = Z;
		19'b1000010000110001101: color_data = Z;
		19'b1000010000110001110: color_data = Z;
		19'b1000010000110001111: color_data = Z;
		19'b1000010000110010000: color_data = Z;
		19'b1000010000110010001: color_data = Z;
		19'b1000010000110010010: color_data = Z;
		19'b1000010000110010011: color_data = Z;
		19'b1000010000110010100: color_data = Z;
		19'b1000010000110010101: color_data = Z;
		19'b1000010000110010110: color_data = Z;
		19'b1000010000110010111: color_data = Z;
		19'b1000010000110011000: color_data = Z;
		19'b1000010000110011001: color_data = Z;
		19'b1000010000110011010: color_data = Z;
		19'b1000010000110011011: color_data = Z;
		19'b1000010000110011100: color_data = Z;
		19'b1000010000110011101: color_data = Z;
		19'b1000010000110011110: color_data = Z;
		19'b1000010000110011111: color_data = Z;
		19'b1000010000110100000: color_data = Z;
		19'b1000010000110100001: color_data = Z;
		19'b1000010000110100010: color_data = Z;
		19'b1000010000110100011: color_data = Z;
		19'b1000010000110100100: color_data = Z;
		19'b1000010000110100101: color_data = Z;
		19'b1000010000110100110: color_data = Z;
		19'b1000010000110100111: color_data = Z;
		19'b1000010000110101000: color_data = Z;
		19'b1000010000110101001: color_data = Z;
		19'b1000010000110101010: color_data = Z;
		19'b1000010000110101011: color_data = Z;
		19'b1000010000110101100: color_data = Z;
		19'b1000010000110101101: color_data = Z;
		19'b1000010000110101110: color_data = Z;
		19'b1000010000110101111: color_data = Z;
		19'b1000010000110110000: color_data = Z;
		19'b1000010000110110001: color_data = Z;
		19'b1000010000110110010: color_data = Z;
		19'b1000010000110110011: color_data = Z;
		19'b1000010000110110100: color_data = Z;
		19'b1000010000110110101: color_data = Z;
		19'b1000010000110110110: color_data = Z;
		19'b1000010000110110111: color_data = Z;
		19'b1000010000110111000: color_data = Z;
		19'b1000010000110111001: color_data = Z;
		19'b1000010000110111010: color_data = Z;
		19'b1000010000110111011: color_data = Z;
		19'b1000010000110111100: color_data = Z;
		19'b1000010000110111101: color_data = Z;
		19'b1000010000111000010: color_data = Z;
		19'b1000010000111000011: color_data = Z;
		19'b1000010000111000100: color_data = Z;
		19'b1000010000111000101: color_data = Z;
		19'b1000010000111000110: color_data = Z;
		19'b1000010000111000111: color_data = Z;
		19'b1000010000111001000: color_data = Z;
		19'b1000010000111001001: color_data = Z;
		19'b1000010000111001010: color_data = Z;
		19'b1000010000111001011: color_data = Z;
		19'b1000010000111001100: color_data = Z;
		19'b1000010010010111010: color_data = Z;
		19'b1000010010010111011: color_data = Z;
		19'b1000010010010111100: color_data = Z;
		19'b1000010010010111101: color_data = Z;
		19'b1000010010010111110: color_data = Z;
		19'b1000010010010111111: color_data = Z;
		19'b1000010010011000000: color_data = Z;
		19'b1000010010011000001: color_data = Z;
		19'b1000010010011000010: color_data = Z;
		19'b1000010010011000011: color_data = Z;
		19'b1000010010011000100: color_data = Z;
		19'b1000010010011000101: color_data = Z;
		19'b1000010010011000110: color_data = Z;
		19'b1000010010011000111: color_data = Z;
		19'b1000010010011001000: color_data = Z;
		19'b1000010010011001001: color_data = Z;
		19'b1000010010011001010: color_data = Z;
		19'b1000010010011001011: color_data = Z;
		19'b1000010010011001100: color_data = Z;
		19'b1000010010011001101: color_data = Z;
		19'b1000010010011001110: color_data = Z;
		19'b1000010010011001111: color_data = Z;
		19'b1000010010011111100: color_data = Z;
		19'b1000010010011111101: color_data = Z;
		19'b1000010010011111110: color_data = Z;
		19'b1000010010011111111: color_data = Z;
		19'b1000010010100000000: color_data = Z;
		19'b1000010010100000001: color_data = Z;
		19'b1000010010100000010: color_data = Z;
		19'b1000010010100000011: color_data = Z;
		19'b1000010010100000100: color_data = Z;
		19'b1000010010100000101: color_data = Z;
		19'b1000010010100000110: color_data = Z;
		19'b1000010010100000111: color_data = Z;
		19'b1000010010100001000: color_data = Z;
		19'b1000010010100001001: color_data = Z;
		19'b1000010010100001010: color_data = Z;
		19'b1000010010100001011: color_data = Z;
		19'b1000010010100001100: color_data = Z;
		19'b1000010010100001101: color_data = Z;
		19'b1000010010100001110: color_data = Z;
		19'b1000010010100001111: color_data = Z;
		19'b1000010010100010000: color_data = Z;
		19'b1000010010100010001: color_data = Z;
		19'b1000010010100010010: color_data = Z;
		19'b1000010010100010011: color_data = Z;
		19'b1000010010100010100: color_data = Z;
		19'b1000010010100010101: color_data = Z;
		19'b1000010010100010110: color_data = Z;
		19'b1000010010100010111: color_data = Z;
		19'b1000010010100011000: color_data = Z;
		19'b1000010010100011001: color_data = Z;
		19'b1000010010100011010: color_data = Z;
		19'b1000010010100011011: color_data = Z;
		19'b1000010010100011100: color_data = Z;
		19'b1000010010100011101: color_data = Z;
		19'b1000010010100011110: color_data = Z;
		19'b1000010010100011111: color_data = Z;
		19'b1000010010100100000: color_data = Z;
		19'b1000010010100100001: color_data = Z;
		19'b1000010010100100010: color_data = Z;
		19'b1000010010100100011: color_data = Z;
		19'b1000010010100100100: color_data = Z;
		19'b1000010010100100101: color_data = Z;
		19'b1000010010100100110: color_data = Z;
		19'b1000010010100100111: color_data = Z;
		19'b1000010010100101000: color_data = Z;
		19'b1000010010100101001: color_data = Z;
		19'b1000010010100101010: color_data = Z;
		19'b1000010010100101011: color_data = Z;
		19'b1000010010100101100: color_data = Z;
		19'b1000010010100101101: color_data = Z;
		19'b1000010010100101110: color_data = Z;
		19'b1000010010100111001: color_data = Z;
		19'b1000010010101001111: color_data = Z;
		19'b1000010010101010000: color_data = Z;
		19'b1000010010101010001: color_data = Z;
		19'b1000010010101010010: color_data = Z;
		19'b1000010010101010011: color_data = Z;
		19'b1000010010101010100: color_data = Z;
		19'b1000010010101010101: color_data = Z;
		19'b1000010010101010110: color_data = Z;
		19'b1000010010101010111: color_data = Z;
		19'b1000010010101101010: color_data = Z;
		19'b1000010010101101011: color_data = Z;
		19'b1000010010101101100: color_data = Z;
		19'b1000010010101101101: color_data = Z;
		19'b1000010010101101110: color_data = Z;
		19'b1000010010101101111: color_data = Z;
		19'b1000010010101110000: color_data = Z;
		19'b1000010010101110001: color_data = Z;
		19'b1000010010101110010: color_data = Z;
		19'b1000010010101110011: color_data = Z;
		19'b1000010010101110100: color_data = Z;
		19'b1000010010101110101: color_data = Z;
		19'b1000010010101110110: color_data = Z;
		19'b1000010010101110111: color_data = Z;
		19'b1000010010101111000: color_data = Z;
		19'b1000010010101111001: color_data = Z;
		19'b1000010010101111010: color_data = Z;
		19'b1000010010101111011: color_data = Z;
		19'b1000010010101111100: color_data = Z;
		19'b1000010010101111101: color_data = Z;
		19'b1000010010101111110: color_data = Z;
		19'b1000010010101111111: color_data = Z;
		19'b1000010010110000000: color_data = Z;
		19'b1000010010110000001: color_data = Z;
		19'b1000010010110000010: color_data = Z;
		19'b1000010010110000011: color_data = Z;
		19'b1000010010110000100: color_data = Z;
		19'b1000010010110000101: color_data = Z;
		19'b1000010010110000110: color_data = Z;
		19'b1000010010110000111: color_data = Z;
		19'b1000010010110001000: color_data = Z;
		19'b1000010010110001001: color_data = Z;
		19'b1000010010110001010: color_data = Z;
		19'b1000010010110001011: color_data = Z;
		19'b1000010010110001100: color_data = Z;
		19'b1000010010110001101: color_data = Z;
		19'b1000010010110001110: color_data = Z;
		19'b1000010010110001111: color_data = Z;
		19'b1000010010110010000: color_data = Z;
		19'b1000010010110010001: color_data = Z;
		19'b1000010010110010010: color_data = Z;
		19'b1000010010110010011: color_data = Z;
		19'b1000010010110010100: color_data = Z;
		19'b1000010010110010101: color_data = Z;
		19'b1000010010110010110: color_data = Z;
		19'b1000010010110010111: color_data = Z;
		19'b1000010010110011000: color_data = Z;
		19'b1000010010110011001: color_data = Z;
		19'b1000010010110011010: color_data = Z;
		19'b1000010010110011011: color_data = Z;
		19'b1000010010110011100: color_data = Z;
		19'b1000010010110011101: color_data = Z;
		19'b1000010010110011110: color_data = Z;
		19'b1000010010110011111: color_data = Z;
		19'b1000010010110100000: color_data = Z;
		19'b1000010010110100001: color_data = Z;
		19'b1000010010110100010: color_data = Z;
		19'b1000010010110100011: color_data = Z;
		19'b1000010010110100100: color_data = Z;
		19'b1000010010110100101: color_data = Z;
		19'b1000010010110100110: color_data = Z;
		19'b1000010010110100111: color_data = Z;
		19'b1000010010110101000: color_data = Z;
		19'b1000010010110101001: color_data = Z;
		19'b1000010010110101010: color_data = Z;
		19'b1000010010110101011: color_data = Z;
		19'b1000010010110101100: color_data = Z;
		19'b1000010010110101101: color_data = Z;
		19'b1000010010110101110: color_data = Z;
		19'b1000010010110101111: color_data = Z;
		19'b1000010010110110000: color_data = Z;
		19'b1000010010110110001: color_data = Z;
		19'b1000010010110110010: color_data = Z;
		19'b1000010010110110011: color_data = Z;
		19'b1000010010110110100: color_data = Z;
		19'b1000010010110110101: color_data = Z;
		19'b1000010010110110110: color_data = Z;
		19'b1000010010110110111: color_data = Z;
		19'b1000010010110111000: color_data = Z;
		19'b1000010010110111001: color_data = Z;
		19'b1000010010110111010: color_data = Z;
		19'b1000010010110111011: color_data = Z;
		19'b1000010010110111100: color_data = Z;
		19'b1000010010110111101: color_data = Z;
		19'b1000010010111000011: color_data = Z;
		19'b1000010010111000100: color_data = Z;
		19'b1000010010111000101: color_data = Z;
		19'b1000010010111000110: color_data = Z;
		19'b1000010010111000111: color_data = Z;
		19'b1000010010111001000: color_data = Z;
		19'b1000010010111001001: color_data = Z;
		19'b1000010010111001010: color_data = Z;
		19'b1000010010111001011: color_data = Z;
		19'b1000010010111001100: color_data = Z;
		19'b1000010100010111011: color_data = Z;
		19'b1000010100010111100: color_data = Z;
		19'b1000010100010111101: color_data = Z;
		19'b1000010100010111110: color_data = Z;
		19'b1000010100010111111: color_data = Z;
		19'b1000010100011000000: color_data = Z;
		19'b1000010100011000001: color_data = Z;
		19'b1000010100011000010: color_data = Z;
		19'b1000010100011000011: color_data = Z;
		19'b1000010100011000100: color_data = Z;
		19'b1000010100011000101: color_data = Z;
		19'b1000010100011000110: color_data = Z;
		19'b1000010100011000111: color_data = Z;
		19'b1000010100011001000: color_data = Z;
		19'b1000010100011001001: color_data = Z;
		19'b1000010100011001010: color_data = Z;
		19'b1000010100011001011: color_data = Z;
		19'b1000010100011001100: color_data = Z;
		19'b1000010100011001101: color_data = Z;
		19'b1000010100011001110: color_data = Z;
		19'b1000010100011001111: color_data = Z;
		19'b1000010100011010000: color_data = Z;
		19'b1000010100011111010: color_data = Z;
		19'b1000010100011111011: color_data = Z;
		19'b1000010100011111100: color_data = Z;
		19'b1000010100011111101: color_data = Z;
		19'b1000010100011111110: color_data = Z;
		19'b1000010100011111111: color_data = Z;
		19'b1000010100100000000: color_data = Z;
		19'b1000010100100000001: color_data = Z;
		19'b1000010100100000010: color_data = Z;
		19'b1000010100100000011: color_data = Z;
		19'b1000010100100000100: color_data = Z;
		19'b1000010100100000101: color_data = Z;
		19'b1000010100100000110: color_data = Z;
		19'b1000010100100000111: color_data = Z;
		19'b1000010100100001000: color_data = Z;
		19'b1000010100100001001: color_data = Z;
		19'b1000010100100001010: color_data = Z;
		19'b1000010100100001011: color_data = Z;
		19'b1000010100100001100: color_data = Z;
		19'b1000010100100001101: color_data = Z;
		19'b1000010100100001110: color_data = Z;
		19'b1000010100100001111: color_data = Z;
		19'b1000010100100010000: color_data = Z;
		19'b1000010100100010001: color_data = Z;
		19'b1000010100100010010: color_data = Z;
		19'b1000010100100010011: color_data = Z;
		19'b1000010100100010100: color_data = Z;
		19'b1000010100100010101: color_data = Z;
		19'b1000010100100010110: color_data = Z;
		19'b1000010100100010111: color_data = Z;
		19'b1000010100100011000: color_data = Z;
		19'b1000010100100011001: color_data = Z;
		19'b1000010100100011010: color_data = Z;
		19'b1000010100100011011: color_data = Z;
		19'b1000010100100011100: color_data = Z;
		19'b1000010100100011101: color_data = Z;
		19'b1000010100100011110: color_data = Z;
		19'b1000010100100011111: color_data = Z;
		19'b1000010100100100000: color_data = Z;
		19'b1000010100100100001: color_data = Z;
		19'b1000010100100100010: color_data = Z;
		19'b1000010100100100011: color_data = Z;
		19'b1000010100100100100: color_data = Z;
		19'b1000010100100100101: color_data = Z;
		19'b1000010100100100110: color_data = Z;
		19'b1000010100100100111: color_data = Z;
		19'b1000010100100101000: color_data = Z;
		19'b1000010100100101001: color_data = Z;
		19'b1000010100100101010: color_data = Z;
		19'b1000010100100101011: color_data = Z;
		19'b1000010100100101100: color_data = Z;
		19'b1000010100100101101: color_data = Z;
		19'b1000010100100101110: color_data = Z;
		19'b1000010100100101111: color_data = Z;
		19'b1000010100100111001: color_data = Z;
		19'b1000010100101010011: color_data = Z;
		19'b1000010100101010100: color_data = Z;
		19'b1000010100101010101: color_data = Z;
		19'b1000010100101010110: color_data = Z;
		19'b1000010100101010111: color_data = Z;
		19'b1000010100101101001: color_data = Z;
		19'b1000010100101101010: color_data = Z;
		19'b1000010100101101011: color_data = Z;
		19'b1000010100101101100: color_data = Z;
		19'b1000010100101101101: color_data = Z;
		19'b1000010100101101110: color_data = Z;
		19'b1000010100101101111: color_data = Z;
		19'b1000010100101110000: color_data = Z;
		19'b1000010100101110001: color_data = Z;
		19'b1000010100101110010: color_data = Z;
		19'b1000010100101110011: color_data = Z;
		19'b1000010100101110100: color_data = Z;
		19'b1000010100101110101: color_data = Z;
		19'b1000010100101110110: color_data = Z;
		19'b1000010100101110111: color_data = Z;
		19'b1000010100101111000: color_data = Z;
		19'b1000010100101111001: color_data = Z;
		19'b1000010100101111010: color_data = Z;
		19'b1000010100101111011: color_data = Z;
		19'b1000010100101111100: color_data = Z;
		19'b1000010100101111101: color_data = Z;
		19'b1000010100101111110: color_data = Z;
		19'b1000010100101111111: color_data = Z;
		19'b1000010100110000000: color_data = Z;
		19'b1000010100110000001: color_data = Z;
		19'b1000010100110000010: color_data = Z;
		19'b1000010100110000011: color_data = Z;
		19'b1000010100110000100: color_data = Z;
		19'b1000010100110000101: color_data = Z;
		19'b1000010100110000110: color_data = Z;
		19'b1000010100110000111: color_data = Z;
		19'b1000010100110001000: color_data = Z;
		19'b1000010100110001001: color_data = Z;
		19'b1000010100110001010: color_data = Z;
		19'b1000010100110001011: color_data = Z;
		19'b1000010100110001100: color_data = Z;
		19'b1000010100110001101: color_data = Z;
		19'b1000010100110001110: color_data = Z;
		19'b1000010100110001111: color_data = Z;
		19'b1000010100110010000: color_data = Z;
		19'b1000010100110010001: color_data = Z;
		19'b1000010100110010010: color_data = Z;
		19'b1000010100110010011: color_data = Z;
		19'b1000010100110010100: color_data = Z;
		19'b1000010100110010101: color_data = Z;
		19'b1000010100110010110: color_data = Z;
		19'b1000010100110010111: color_data = Z;
		19'b1000010100110011000: color_data = Z;
		19'b1000010100110011001: color_data = Z;
		19'b1000010100110011010: color_data = Z;
		19'b1000010100110011011: color_data = Z;
		19'b1000010100110011100: color_data = Z;
		19'b1000010100110011101: color_data = Z;
		19'b1000010100110011110: color_data = Z;
		19'b1000010100110011111: color_data = Z;
		19'b1000010100110100000: color_data = Z;
		19'b1000010100110100001: color_data = Z;
		19'b1000010100110100010: color_data = Z;
		19'b1000010100110100011: color_data = Z;
		19'b1000010100110100100: color_data = Z;
		19'b1000010100110100101: color_data = Z;
		19'b1000010100110100110: color_data = Z;
		19'b1000010100110100111: color_data = Z;
		19'b1000010100110101000: color_data = Z;
		19'b1000010100110101001: color_data = Z;
		19'b1000010100110101010: color_data = Z;
		19'b1000010100110101011: color_data = Z;
		19'b1000010100110101100: color_data = Z;
		19'b1000010100110101101: color_data = Z;
		19'b1000010100110101110: color_data = Z;
		19'b1000010100110101111: color_data = Z;
		19'b1000010100110110000: color_data = Z;
		19'b1000010100110110001: color_data = Z;
		19'b1000010100110110010: color_data = Z;
		19'b1000010100110110011: color_data = Z;
		19'b1000010100110110100: color_data = Z;
		19'b1000010100110110101: color_data = Z;
		19'b1000010100110110110: color_data = Z;
		19'b1000010100110110111: color_data = Z;
		19'b1000010100110111000: color_data = Z;
		19'b1000010100110111001: color_data = Z;
		19'b1000010100110111010: color_data = Z;
		19'b1000010100110111011: color_data = Z;
		19'b1000010100110111100: color_data = Z;
		19'b1000010100110111101: color_data = Z;
		19'b1000010100111000100: color_data = Z;
		19'b1000010100111000101: color_data = Z;
		19'b1000010100111000110: color_data = Z;
		19'b1000010100111000111: color_data = Z;
		19'b1000010100111001000: color_data = Z;
		19'b1000010100111001001: color_data = Z;
		19'b1000010100111001010: color_data = Z;
		19'b1000010100111001011: color_data = Z;
		19'b1000010100111001100: color_data = Z;
		19'b1000010110010111011: color_data = Z;
		19'b1000010110010111100: color_data = Z;
		19'b1000010110010111101: color_data = Z;
		19'b1000010110010111110: color_data = Z;
		19'b1000010110010111111: color_data = Z;
		19'b1000010110011000000: color_data = Z;
		19'b1000010110011000001: color_data = Z;
		19'b1000010110011000010: color_data = Z;
		19'b1000010110011000011: color_data = Z;
		19'b1000010110011000100: color_data = Z;
		19'b1000010110011000101: color_data = Z;
		19'b1000010110011000110: color_data = Z;
		19'b1000010110011000111: color_data = Z;
		19'b1000010110011001000: color_data = Z;
		19'b1000010110011001001: color_data = Z;
		19'b1000010110011001010: color_data = Z;
		19'b1000010110011001011: color_data = Z;
		19'b1000010110011001100: color_data = Z;
		19'b1000010110011001101: color_data = Z;
		19'b1000010110011001110: color_data = Z;
		19'b1000010110011001111: color_data = Z;
		19'b1000010110011010000: color_data = Z;
		19'b1000010110011010001: color_data = Z;
		19'b1000010110011010010: color_data = Z;
		19'b1000010110011111000: color_data = Z;
		19'b1000010110011111001: color_data = Z;
		19'b1000010110011111010: color_data = Z;
		19'b1000010110011111011: color_data = Z;
		19'b1000010110011111100: color_data = Z;
		19'b1000010110011111101: color_data = Z;
		19'b1000010110011111110: color_data = Z;
		19'b1000010110011111111: color_data = Z;
		19'b1000010110100000000: color_data = Z;
		19'b1000010110100000001: color_data = Z;
		19'b1000010110100000010: color_data = Z;
		19'b1000010110100000011: color_data = Z;
		19'b1000010110100000100: color_data = Z;
		19'b1000010110100000101: color_data = Z;
		19'b1000010110100000110: color_data = Z;
		19'b1000010110100000111: color_data = Z;
		19'b1000010110100001000: color_data = Z;
		19'b1000010110100001001: color_data = Z;
		19'b1000010110100001010: color_data = Z;
		19'b1000010110100001011: color_data = Z;
		19'b1000010110100001100: color_data = Z;
		19'b1000010110100001101: color_data = Z;
		19'b1000010110100001110: color_data = Z;
		19'b1000010110100001111: color_data = Z;
		19'b1000010110100010000: color_data = Z;
		19'b1000010110100010001: color_data = Z;
		19'b1000010110100010010: color_data = Z;
		19'b1000010110100010011: color_data = Z;
		19'b1000010110100010100: color_data = Z;
		19'b1000010110100010101: color_data = Z;
		19'b1000010110100010110: color_data = Z;
		19'b1000010110100010111: color_data = Z;
		19'b1000010110100011000: color_data = Z;
		19'b1000010110100011001: color_data = Z;
		19'b1000010110100011010: color_data = Z;
		19'b1000010110100011011: color_data = Z;
		19'b1000010110100011100: color_data = Z;
		19'b1000010110100011101: color_data = Z;
		19'b1000010110100011110: color_data = Z;
		19'b1000010110100011111: color_data = Z;
		19'b1000010110100100000: color_data = Z;
		19'b1000010110100100001: color_data = Z;
		19'b1000010110100100010: color_data = Z;
		19'b1000010110100100011: color_data = Z;
		19'b1000010110100100100: color_data = Z;
		19'b1000010110100100101: color_data = Z;
		19'b1000010110100100110: color_data = Z;
		19'b1000010110100100111: color_data = Z;
		19'b1000010110100101000: color_data = Z;
		19'b1000010110100101001: color_data = Z;
		19'b1000010110100101010: color_data = Z;
		19'b1000010110100101011: color_data = Z;
		19'b1000010110100101100: color_data = Z;
		19'b1000010110100101101: color_data = Z;
		19'b1000010110100101110: color_data = Z;
		19'b1000010110100101111: color_data = Z;
		19'b1000010110101010101: color_data = Z;
		19'b1000010110101010110: color_data = Z;
		19'b1000010110101010111: color_data = Z;
		19'b1000010110101101001: color_data = Z;
		19'b1000010110101101010: color_data = Z;
		19'b1000010110101101011: color_data = Z;
		19'b1000010110101101100: color_data = Z;
		19'b1000010110101101101: color_data = Z;
		19'b1000010110101101110: color_data = Z;
		19'b1000010110101101111: color_data = Z;
		19'b1000010110101110000: color_data = Z;
		19'b1000010110101110001: color_data = Z;
		19'b1000010110101110010: color_data = Z;
		19'b1000010110101110011: color_data = Z;
		19'b1000010110101110100: color_data = Z;
		19'b1000010110101110101: color_data = Z;
		19'b1000010110101110110: color_data = Z;
		19'b1000010110101110111: color_data = Z;
		19'b1000010110101111000: color_data = Z;
		19'b1000010110101111001: color_data = Z;
		19'b1000010110101111010: color_data = Z;
		19'b1000010110101111011: color_data = Z;
		19'b1000010110101111100: color_data = Z;
		19'b1000010110101111101: color_data = Z;
		19'b1000010110101111110: color_data = Z;
		19'b1000010110101111111: color_data = Z;
		19'b1000010110110000000: color_data = Z;
		19'b1000010110110000001: color_data = Z;
		19'b1000010110110000010: color_data = Z;
		19'b1000010110110000011: color_data = Z;
		19'b1000010110110000100: color_data = Z;
		19'b1000010110110000101: color_data = Z;
		19'b1000010110110000110: color_data = Z;
		19'b1000010110110000111: color_data = Z;
		19'b1000010110110001000: color_data = Z;
		19'b1000010110110001001: color_data = Z;
		19'b1000010110110001010: color_data = Z;
		19'b1000010110110001011: color_data = Z;
		19'b1000010110110001100: color_data = Z;
		19'b1000010110110001101: color_data = Z;
		19'b1000010110110001110: color_data = Z;
		19'b1000010110110001111: color_data = Z;
		19'b1000010110110010000: color_data = Z;
		19'b1000010110110010001: color_data = Z;
		19'b1000010110110010010: color_data = Z;
		19'b1000010110110010011: color_data = Z;
		19'b1000010110110010100: color_data = Z;
		19'b1000010110110010101: color_data = Z;
		19'b1000010110110010110: color_data = Z;
		19'b1000010110110010111: color_data = Z;
		19'b1000010110110011000: color_data = Z;
		19'b1000010110110011001: color_data = Z;
		19'b1000010110110011010: color_data = Z;
		19'b1000010110110011011: color_data = Z;
		19'b1000010110110011100: color_data = Z;
		19'b1000010110110011101: color_data = Z;
		19'b1000010110110011110: color_data = Z;
		19'b1000010110110011111: color_data = Z;
		19'b1000010110110100000: color_data = Z;
		19'b1000010110110100001: color_data = Z;
		19'b1000010110110100010: color_data = Z;
		19'b1000010110110100011: color_data = Z;
		19'b1000010110110100100: color_data = Z;
		19'b1000010110110100101: color_data = Z;
		19'b1000010110110100110: color_data = Z;
		19'b1000010110110100111: color_data = Z;
		19'b1000010110110101000: color_data = Z;
		19'b1000010110110101001: color_data = Z;
		19'b1000010110110101010: color_data = Z;
		19'b1000010110110101011: color_data = Z;
		19'b1000010110110101100: color_data = Z;
		19'b1000010110110101101: color_data = Z;
		19'b1000010110110101110: color_data = Z;
		19'b1000010110110101111: color_data = Z;
		19'b1000010110110110000: color_data = Z;
		19'b1000010110110110001: color_data = Z;
		19'b1000010110110110010: color_data = Z;
		19'b1000010110110110011: color_data = Z;
		19'b1000010110110110100: color_data = Z;
		19'b1000010110110110101: color_data = Z;
		19'b1000010110110110110: color_data = Z;
		19'b1000010110110110111: color_data = Z;
		19'b1000010110110111000: color_data = Z;
		19'b1000010110110111001: color_data = Z;
		19'b1000010110110111010: color_data = Z;
		19'b1000010110110111011: color_data = Z;
		19'b1000010110110111100: color_data = Z;
		19'b1000010110110111101: color_data = Z;
		19'b1000010110111000101: color_data = Z;
		19'b1000010110111000110: color_data = Z;
		19'b1000010110111000111: color_data = Z;
		19'b1000010110111001000: color_data = Z;
		19'b1000010110111001001: color_data = Z;
		19'b1000010110111001010: color_data = Z;
		19'b1000010110111001011: color_data = Z;
		19'b1000010110111001100: color_data = Z;
		19'b1000011000010111100: color_data = Z;
		19'b1000011000010111101: color_data = Z;
		19'b1000011000010111110: color_data = Z;
		19'b1000011000010111111: color_data = Z;
		19'b1000011000011000000: color_data = Z;
		19'b1000011000011000001: color_data = Z;
		19'b1000011000011000010: color_data = Z;
		19'b1000011000011000011: color_data = Z;
		19'b1000011000011000100: color_data = Z;
		19'b1000011000011000101: color_data = Z;
		19'b1000011000011000110: color_data = Z;
		19'b1000011000011000111: color_data = Z;
		19'b1000011000011001000: color_data = Z;
		19'b1000011000011001001: color_data = Z;
		19'b1000011000011001010: color_data = Z;
		19'b1000011000011001011: color_data = Z;
		19'b1000011000011001100: color_data = Z;
		19'b1000011000011001101: color_data = Z;
		19'b1000011000011001110: color_data = Z;
		19'b1000011000011001111: color_data = Z;
		19'b1000011000011010000: color_data = Z;
		19'b1000011000011010001: color_data = Z;
		19'b1000011000011010010: color_data = Z;
		19'b1000011000011010011: color_data = Z;
		19'b1000011000011010100: color_data = Z;
		19'b1000011000011010101: color_data = Z;
		19'b1000011000011011100: color_data = Z;
		19'b1000011000011011101: color_data = Z;
		19'b1000011000011110110: color_data = Z;
		19'b1000011000011110111: color_data = Z;
		19'b1000011000011111000: color_data = Z;
		19'b1000011000011111001: color_data = Z;
		19'b1000011000011111010: color_data = Z;
		19'b1000011000011111011: color_data = Z;
		19'b1000011000011111100: color_data = Z;
		19'b1000011000011111101: color_data = Z;
		19'b1000011000011111110: color_data = Z;
		19'b1000011000011111111: color_data = Z;
		19'b1000011000100000000: color_data = Z;
		19'b1000011000100000001: color_data = Z;
		19'b1000011000100000010: color_data = Z;
		19'b1000011000100000011: color_data = Z;
		19'b1000011000100000100: color_data = Z;
		19'b1000011000100000101: color_data = Z;
		19'b1000011000100000110: color_data = Z;
		19'b1000011000100000111: color_data = Z;
		19'b1000011000100001000: color_data = Z;
		19'b1000011000100001001: color_data = Z;
		19'b1000011000100001010: color_data = Z;
		19'b1000011000100001011: color_data = Z;
		19'b1000011000100001100: color_data = Z;
		19'b1000011000100001101: color_data = Z;
		19'b1000011000100001110: color_data = Z;
		19'b1000011000100001111: color_data = Z;
		19'b1000011000100010000: color_data = Z;
		19'b1000011000100010001: color_data = Z;
		19'b1000011000100010010: color_data = Z;
		19'b1000011000100010011: color_data = Z;
		19'b1000011000100010100: color_data = Z;
		19'b1000011000100010101: color_data = Z;
		19'b1000011000100010110: color_data = Z;
		19'b1000011000100010111: color_data = Z;
		19'b1000011000100011000: color_data = Z;
		19'b1000011000100011001: color_data = Z;
		19'b1000011000100011010: color_data = Z;
		19'b1000011000100011011: color_data = Z;
		19'b1000011000100011100: color_data = Z;
		19'b1000011000100011101: color_data = Z;
		19'b1000011000100011110: color_data = Z;
		19'b1000011000100011111: color_data = Z;
		19'b1000011000100100000: color_data = Z;
		19'b1000011000100100001: color_data = Z;
		19'b1000011000100100010: color_data = Z;
		19'b1000011000100100011: color_data = Z;
		19'b1000011000100100100: color_data = Z;
		19'b1000011000100100101: color_data = Z;
		19'b1000011000100100110: color_data = Z;
		19'b1000011000100100111: color_data = Z;
		19'b1000011000100101000: color_data = Z;
		19'b1000011000100101001: color_data = Z;
		19'b1000011000100101010: color_data = Z;
		19'b1000011000100101011: color_data = Z;
		19'b1000011000100101100: color_data = Z;
		19'b1000011000100101101: color_data = Z;
		19'b1000011000100101110: color_data = Z;
		19'b1000011000100101111: color_data = Z;
		19'b1000011000101010101: color_data = Z;
		19'b1000011000101010110: color_data = Z;
		19'b1000011000101010111: color_data = Z;
		19'b1000011000101101000: color_data = Z;
		19'b1000011000101101001: color_data = Z;
		19'b1000011000101101010: color_data = Z;
		19'b1000011000101101011: color_data = Z;
		19'b1000011000101101100: color_data = Z;
		19'b1000011000101101101: color_data = Z;
		19'b1000011000101101110: color_data = Z;
		19'b1000011000101101111: color_data = Z;
		19'b1000011000101110000: color_data = Z;
		19'b1000011000101110001: color_data = Z;
		19'b1000011000101110010: color_data = Z;
		19'b1000011000101110011: color_data = Z;
		19'b1000011000101110100: color_data = Z;
		19'b1000011000101110101: color_data = Z;
		19'b1000011000101110110: color_data = Z;
		19'b1000011000101110111: color_data = Z;
		19'b1000011000101111000: color_data = Z;
		19'b1000011000101111001: color_data = Z;
		19'b1000011000101111010: color_data = Z;
		19'b1000011000101111011: color_data = Z;
		19'b1000011000101111100: color_data = Z;
		19'b1000011000101111101: color_data = Z;
		19'b1000011000101111110: color_data = Z;
		19'b1000011000101111111: color_data = Z;
		19'b1000011000110000000: color_data = Z;
		19'b1000011000110000001: color_data = Z;
		19'b1000011000110000010: color_data = Z;
		19'b1000011000110000011: color_data = Z;
		19'b1000011000110000100: color_data = Z;
		19'b1000011000110000101: color_data = Z;
		19'b1000011000110000110: color_data = Z;
		19'b1000011000110000111: color_data = Z;
		19'b1000011000110001000: color_data = Z;
		19'b1000011000110001001: color_data = Z;
		19'b1000011000110001010: color_data = Z;
		19'b1000011000110001011: color_data = Z;
		19'b1000011000110001100: color_data = Z;
		19'b1000011000110001101: color_data = Z;
		19'b1000011000110001110: color_data = Z;
		19'b1000011000110001111: color_data = Z;
		19'b1000011000110010000: color_data = Z;
		19'b1000011000110010001: color_data = Z;
		19'b1000011000110010010: color_data = Z;
		19'b1000011000110010011: color_data = Z;
		19'b1000011000110010100: color_data = Z;
		19'b1000011000110010101: color_data = Z;
		19'b1000011000110010110: color_data = Z;
		19'b1000011000110010111: color_data = Z;
		19'b1000011000110011000: color_data = Z;
		19'b1000011000110011001: color_data = Z;
		19'b1000011000110011010: color_data = Z;
		19'b1000011000110011011: color_data = Z;
		19'b1000011000110011100: color_data = Z;
		19'b1000011000110011101: color_data = Z;
		19'b1000011000110011110: color_data = Z;
		19'b1000011000110011111: color_data = Z;
		19'b1000011000110100000: color_data = Z;
		19'b1000011000110100001: color_data = Z;
		19'b1000011000110100010: color_data = Z;
		19'b1000011000110100011: color_data = Z;
		19'b1000011000110100100: color_data = Z;
		19'b1000011000110100101: color_data = Z;
		19'b1000011000110100110: color_data = Z;
		19'b1000011000110100111: color_data = Z;
		19'b1000011000110101000: color_data = Z;
		19'b1000011000110101001: color_data = Z;
		19'b1000011000110101010: color_data = Z;
		19'b1000011000110101011: color_data = Z;
		19'b1000011000110101100: color_data = Z;
		19'b1000011000110101101: color_data = Z;
		19'b1000011000110101110: color_data = Z;
		19'b1000011000110101111: color_data = Z;
		19'b1000011000110110000: color_data = Z;
		19'b1000011000110110001: color_data = Z;
		19'b1000011000110110010: color_data = Z;
		19'b1000011000110110011: color_data = Z;
		19'b1000011000110110100: color_data = Z;
		19'b1000011000110110101: color_data = Z;
		19'b1000011000110110110: color_data = Z;
		19'b1000011000110110111: color_data = Z;
		19'b1000011000110111000: color_data = Z;
		19'b1000011000110111001: color_data = Z;
		19'b1000011000110111010: color_data = Z;
		19'b1000011000110111011: color_data = Z;
		19'b1000011000110111100: color_data = Z;
		19'b1000011000110111101: color_data = Z;
		19'b1000011000111000110: color_data = Z;
		19'b1000011000111000111: color_data = Z;
		19'b1000011000111001000: color_data = Z;
		19'b1000011000111001001: color_data = Z;
		19'b1000011000111001010: color_data = Z;
		19'b1000011000111001011: color_data = Z;
		19'b1000011000111001100: color_data = Z;
		19'b1000011010010111101: color_data = Z;
		19'b1000011010010111110: color_data = Z;
		19'b1000011010010111111: color_data = Z;
		19'b1000011010011000000: color_data = Z;
		19'b1000011010011000001: color_data = Z;
		19'b1000011010011000010: color_data = Z;
		19'b1000011010011000011: color_data = Z;
		19'b1000011010011000100: color_data = Z;
		19'b1000011010011000101: color_data = Z;
		19'b1000011010011000110: color_data = Z;
		19'b1000011010011000111: color_data = Z;
		19'b1000011010011001000: color_data = Z;
		19'b1000011010011001001: color_data = Z;
		19'b1000011010011001010: color_data = Z;
		19'b1000011010011001011: color_data = Z;
		19'b1000011010011001100: color_data = Z;
		19'b1000011010011001101: color_data = Z;
		19'b1000011010011001110: color_data = Z;
		19'b1000011010011001111: color_data = Z;
		19'b1000011010011010000: color_data = Z;
		19'b1000011010011010001: color_data = Z;
		19'b1000011010011010010: color_data = Z;
		19'b1000011010011010011: color_data = Z;
		19'b1000011010011010100: color_data = Z;
		19'b1000011010011010101: color_data = Z;
		19'b1000011010011010110: color_data = Z;
		19'b1000011010011010111: color_data = Z;
		19'b1000011010011011010: color_data = Z;
		19'b1000011010011011011: color_data = Z;
		19'b1000011010011011100: color_data = Z;
		19'b1000011010011011101: color_data = Z;
		19'b1000011010011011110: color_data = Z;
		19'b1000011010011011111: color_data = Z;
		19'b1000011010011100000: color_data = Z;
		19'b1000011010011110010: color_data = Z;
		19'b1000011010011110011: color_data = Z;
		19'b1000011010011110100: color_data = Z;
		19'b1000011010011110101: color_data = Z;
		19'b1000011010011110110: color_data = Z;
		19'b1000011010011110111: color_data = Z;
		19'b1000011010011111000: color_data = Z;
		19'b1000011010011111001: color_data = Z;
		19'b1000011010011111010: color_data = Z;
		19'b1000011010011111011: color_data = Z;
		19'b1000011010011111100: color_data = Z;
		19'b1000011010011111101: color_data = Z;
		19'b1000011010011111110: color_data = Z;
		19'b1000011010011111111: color_data = Z;
		19'b1000011010100000000: color_data = Z;
		19'b1000011010100000001: color_data = Z;
		19'b1000011010100000010: color_data = Z;
		19'b1000011010100000011: color_data = Z;
		19'b1000011010100000100: color_data = Z;
		19'b1000011010100000101: color_data = Z;
		19'b1000011010100000110: color_data = Z;
		19'b1000011010100000111: color_data = Z;
		19'b1000011010100001000: color_data = Z;
		19'b1000011010100001001: color_data = Z;
		19'b1000011010100001010: color_data = Z;
		19'b1000011010100001011: color_data = Z;
		19'b1000011010100001100: color_data = Z;
		19'b1000011010100001101: color_data = Z;
		19'b1000011010100001110: color_data = Z;
		19'b1000011010100001111: color_data = Z;
		19'b1000011010100010000: color_data = Z;
		19'b1000011010100010001: color_data = Z;
		19'b1000011010100010010: color_data = Z;
		19'b1000011010100010011: color_data = Z;
		19'b1000011010100010100: color_data = Z;
		19'b1000011010100010101: color_data = Z;
		19'b1000011010100010110: color_data = Z;
		19'b1000011010100010111: color_data = Z;
		19'b1000011010100011000: color_data = Z;
		19'b1000011010100011001: color_data = Z;
		19'b1000011010100011010: color_data = Z;
		19'b1000011010100011011: color_data = Z;
		19'b1000011010100011100: color_data = Z;
		19'b1000011010100011101: color_data = Z;
		19'b1000011010100011110: color_data = Z;
		19'b1000011010100011111: color_data = Z;
		19'b1000011010100100000: color_data = Z;
		19'b1000011010100100001: color_data = Z;
		19'b1000011010100100010: color_data = Z;
		19'b1000011010100100011: color_data = Z;
		19'b1000011010100100100: color_data = Z;
		19'b1000011010100100101: color_data = Z;
		19'b1000011010100100110: color_data = Z;
		19'b1000011010100100111: color_data = Z;
		19'b1000011010100101000: color_data = Z;
		19'b1000011010100101001: color_data = Z;
		19'b1000011010100101011: color_data = Z;
		19'b1000011010100101100: color_data = Z;
		19'b1000011010100101101: color_data = Z;
		19'b1000011010100101110: color_data = Z;
		19'b1000011010100101111: color_data = Z;
		19'b1000011010101010100: color_data = Z;
		19'b1000011010101010101: color_data = Z;
		19'b1000011010101010110: color_data = Z;
		19'b1000011010101010111: color_data = Z;
		19'b1000011010101101000: color_data = Z;
		19'b1000011010101101001: color_data = Z;
		19'b1000011010101101010: color_data = Z;
		19'b1000011010101101011: color_data = Z;
		19'b1000011010101101100: color_data = Z;
		19'b1000011010101101101: color_data = Z;
		19'b1000011010101101110: color_data = Z;
		19'b1000011010101101111: color_data = Z;
		19'b1000011010101110000: color_data = Z;
		19'b1000011010101110001: color_data = Z;
		19'b1000011010101110010: color_data = Z;
		19'b1000011010101110011: color_data = Z;
		19'b1000011010101110100: color_data = Z;
		19'b1000011010101110101: color_data = Z;
		19'b1000011010101110110: color_data = Z;
		19'b1000011010101110111: color_data = Z;
		19'b1000011010101111000: color_data = Z;
		19'b1000011010101111001: color_data = Z;
		19'b1000011010101111010: color_data = Z;
		19'b1000011010101111011: color_data = Z;
		19'b1000011010101111100: color_data = Z;
		19'b1000011010101111101: color_data = Z;
		19'b1000011010101111110: color_data = Z;
		19'b1000011010101111111: color_data = Z;
		19'b1000011010110000000: color_data = Z;
		19'b1000011010110000001: color_data = Z;
		19'b1000011010110000010: color_data = Z;
		19'b1000011010110000011: color_data = Z;
		19'b1000011010110000100: color_data = Z;
		19'b1000011010110000101: color_data = Z;
		19'b1000011010110000110: color_data = Z;
		19'b1000011010110000111: color_data = Z;
		19'b1000011010110001000: color_data = Z;
		19'b1000011010110001001: color_data = Z;
		19'b1000011010110001010: color_data = Z;
		19'b1000011010110001011: color_data = Z;
		19'b1000011010110001100: color_data = Z;
		19'b1000011010110001101: color_data = Z;
		19'b1000011010110001110: color_data = Z;
		19'b1000011010110001111: color_data = Z;
		19'b1000011010110010000: color_data = Z;
		19'b1000011010110010001: color_data = Z;
		19'b1000011010110010010: color_data = Z;
		19'b1000011010110010011: color_data = Z;
		19'b1000011010110010100: color_data = Z;
		19'b1000011010110010101: color_data = Z;
		19'b1000011010110010110: color_data = Z;
		19'b1000011010110010111: color_data = Z;
		19'b1000011010110011000: color_data = Z;
		19'b1000011010110011001: color_data = Z;
		19'b1000011010110011010: color_data = Z;
		19'b1000011010110011011: color_data = Z;
		19'b1000011010110011100: color_data = Z;
		19'b1000011010110011101: color_data = Z;
		19'b1000011010110011110: color_data = Z;
		19'b1000011010110011111: color_data = Z;
		19'b1000011010110100000: color_data = Z;
		19'b1000011010110100001: color_data = Z;
		19'b1000011010110100010: color_data = Z;
		19'b1000011010110100011: color_data = Z;
		19'b1000011010110100100: color_data = Z;
		19'b1000011010110100101: color_data = Z;
		19'b1000011010110100110: color_data = Z;
		19'b1000011010110100111: color_data = Z;
		19'b1000011010110101000: color_data = Z;
		19'b1000011010110101001: color_data = Z;
		19'b1000011010110101010: color_data = Z;
		19'b1000011010110101011: color_data = Z;
		19'b1000011010110101100: color_data = Z;
		19'b1000011010110101101: color_data = Z;
		19'b1000011010110101110: color_data = Z;
		19'b1000011010110101111: color_data = Z;
		19'b1000011010110110000: color_data = Z;
		19'b1000011010110110001: color_data = Z;
		19'b1000011010110110010: color_data = Z;
		19'b1000011010110110011: color_data = Z;
		19'b1000011010110110100: color_data = Z;
		19'b1000011010110110101: color_data = Z;
		19'b1000011010110110110: color_data = Z;
		19'b1000011010110110111: color_data = Z;
		19'b1000011010110111000: color_data = Z;
		19'b1000011010110111001: color_data = Z;
		19'b1000011010110111010: color_data = Z;
		19'b1000011010110111011: color_data = Z;
		19'b1000011010110111100: color_data = Z;
		19'b1000011010110111101: color_data = Z;
		19'b1000011010111000110: color_data = Z;
		19'b1000011010111000111: color_data = Z;
		19'b1000011010111001000: color_data = Z;
		19'b1000011010111001001: color_data = Z;
		19'b1000011010111001010: color_data = Z;
		19'b1000011010111001011: color_data = Z;
		19'b1000011010111001100: color_data = Z;
		19'b1000011100010111110: color_data = Z;
		19'b1000011100010111111: color_data = Z;
		19'b1000011100011000000: color_data = Z;
		19'b1000011100011000001: color_data = Z;
		19'b1000011100011000010: color_data = Z;
		19'b1000011100011000011: color_data = Z;
		19'b1000011100011000100: color_data = Z;
		19'b1000011100011000101: color_data = Z;
		19'b1000011100011000110: color_data = Z;
		19'b1000011100011000111: color_data = Z;
		19'b1000011100011001000: color_data = Z;
		19'b1000011100011001001: color_data = Z;
		19'b1000011100011001010: color_data = Z;
		19'b1000011100011001011: color_data = Z;
		19'b1000011100011001100: color_data = Z;
		19'b1000011100011001101: color_data = Z;
		19'b1000011100011001110: color_data = Z;
		19'b1000011100011001111: color_data = Z;
		19'b1000011100011010000: color_data = Z;
		19'b1000011100011010001: color_data = Z;
		19'b1000011100011010010: color_data = Z;
		19'b1000011100011010011: color_data = Z;
		19'b1000011100011010100: color_data = Z;
		19'b1000011100011010101: color_data = Z;
		19'b1000011100011010110: color_data = Z;
		19'b1000011100011010111: color_data = Z;
		19'b1000011100011011000: color_data = Z;
		19'b1000011100011011001: color_data = Z;
		19'b1000011100011011010: color_data = Z;
		19'b1000011100011011011: color_data = Z;
		19'b1000011100011011100: color_data = Z;
		19'b1000011100011011101: color_data = Z;
		19'b1000011100011011110: color_data = Z;
		19'b1000011100011011111: color_data = Z;
		19'b1000011100011100000: color_data = Z;
		19'b1000011100011100001: color_data = Z;
		19'b1000011100011100010: color_data = Z;
		19'b1000011100011100011: color_data = Z;
		19'b1000011100011110000: color_data = Z;
		19'b1000011100011110001: color_data = Z;
		19'b1000011100011110010: color_data = Z;
		19'b1000011100011110011: color_data = Z;
		19'b1000011100011110100: color_data = Z;
		19'b1000011100011110101: color_data = Z;
		19'b1000011100011110110: color_data = Z;
		19'b1000011100011110111: color_data = Z;
		19'b1000011100011111000: color_data = Z;
		19'b1000011100011111001: color_data = Z;
		19'b1000011100011111010: color_data = Z;
		19'b1000011100011111011: color_data = Z;
		19'b1000011100011111100: color_data = Z;
		19'b1000011100011111101: color_data = Z;
		19'b1000011100011111110: color_data = Z;
		19'b1000011100011111111: color_data = Z;
		19'b1000011100100000000: color_data = Z;
		19'b1000011100100000001: color_data = Z;
		19'b1000011100100000010: color_data = Z;
		19'b1000011100100000011: color_data = Z;
		19'b1000011100100000100: color_data = Z;
		19'b1000011100100000101: color_data = Z;
		19'b1000011100100000110: color_data = Z;
		19'b1000011100100000111: color_data = Z;
		19'b1000011100100001000: color_data = Z;
		19'b1000011100100001001: color_data = Z;
		19'b1000011100100001010: color_data = Z;
		19'b1000011100100001011: color_data = Z;
		19'b1000011100100001100: color_data = Z;
		19'b1000011100100001101: color_data = Z;
		19'b1000011100100001110: color_data = Z;
		19'b1000011100100001111: color_data = Z;
		19'b1000011100100010000: color_data = Z;
		19'b1000011100100010001: color_data = Z;
		19'b1000011100100010010: color_data = Z;
		19'b1000011100100010011: color_data = Z;
		19'b1000011100100010100: color_data = Z;
		19'b1000011100100010101: color_data = Z;
		19'b1000011100100010110: color_data = Z;
		19'b1000011100100010111: color_data = Z;
		19'b1000011100100011000: color_data = Z;
		19'b1000011100100011001: color_data = Z;
		19'b1000011100100011010: color_data = Z;
		19'b1000011100100011011: color_data = Z;
		19'b1000011100100011100: color_data = Z;
		19'b1000011100100011101: color_data = Z;
		19'b1000011100100011110: color_data = Z;
		19'b1000011100100011111: color_data = Z;
		19'b1000011100100100000: color_data = Z;
		19'b1000011100100100001: color_data = Z;
		19'b1000011100100100010: color_data = Z;
		19'b1000011100100100011: color_data = Z;
		19'b1000011100100100100: color_data = Z;
		19'b1000011100100100101: color_data = Z;
		19'b1000011100100100110: color_data = Z;
		19'b1000011100100100111: color_data = Z;
		19'b1000011100100101000: color_data = Z;
		19'b1000011100100101001: color_data = Z;
		19'b1000011100100101101: color_data = Z;
		19'b1000011100100101110: color_data = Z;
		19'b1000011100100101111: color_data = Z;
		19'b1000011100101010100: color_data = Z;
		19'b1000011100101010101: color_data = Z;
		19'b1000011100101010110: color_data = Z;
		19'b1000011100101100111: color_data = Z;
		19'b1000011100101101000: color_data = Z;
		19'b1000011100101101001: color_data = Z;
		19'b1000011100101101010: color_data = Z;
		19'b1000011100101101011: color_data = Z;
		19'b1000011100101101100: color_data = Z;
		19'b1000011100101101101: color_data = Z;
		19'b1000011100101101110: color_data = Z;
		19'b1000011100101101111: color_data = Z;
		19'b1000011100101110000: color_data = Z;
		19'b1000011100101110001: color_data = Z;
		19'b1000011100101110010: color_data = Z;
		19'b1000011100101110011: color_data = Z;
		19'b1000011100101110100: color_data = Z;
		19'b1000011100101110101: color_data = Z;
		19'b1000011100101110110: color_data = Z;
		19'b1000011100101110111: color_data = Z;
		19'b1000011100101111000: color_data = Z;
		19'b1000011100101111001: color_data = Z;
		19'b1000011100101111010: color_data = Z;
		19'b1000011100101111011: color_data = Z;
		19'b1000011100101111100: color_data = Z;
		19'b1000011100101111101: color_data = Z;
		19'b1000011100101111110: color_data = Z;
		19'b1000011100101111111: color_data = Z;
		19'b1000011100110000000: color_data = Z;
		19'b1000011100110000001: color_data = Z;
		19'b1000011100110000010: color_data = Z;
		19'b1000011100110000011: color_data = Z;
		19'b1000011100110000100: color_data = Z;
		19'b1000011100110000101: color_data = Z;
		19'b1000011100110000110: color_data = Z;
		19'b1000011100110000111: color_data = Z;
		19'b1000011100110001000: color_data = Z;
		19'b1000011100110001001: color_data = Z;
		19'b1000011100110001010: color_data = Z;
		19'b1000011100110001011: color_data = Z;
		19'b1000011100110001100: color_data = Z;
		19'b1000011100110001101: color_data = Z;
		19'b1000011100110001110: color_data = Z;
		19'b1000011100110001111: color_data = Z;
		19'b1000011100110010000: color_data = Z;
		19'b1000011100110010001: color_data = Z;
		19'b1000011100110010010: color_data = Z;
		19'b1000011100110010011: color_data = Z;
		19'b1000011100110010100: color_data = Z;
		19'b1000011100110010101: color_data = Z;
		19'b1000011100110010110: color_data = Z;
		19'b1000011100110010111: color_data = Z;
		19'b1000011100110011000: color_data = Z;
		19'b1000011100110011001: color_data = Z;
		19'b1000011100110011010: color_data = Z;
		19'b1000011100110011011: color_data = Z;
		19'b1000011100110011100: color_data = Z;
		19'b1000011100110011101: color_data = Z;
		19'b1000011100110011110: color_data = Z;
		19'b1000011100110011111: color_data = Z;
		19'b1000011100110100000: color_data = Z;
		19'b1000011100110100001: color_data = Z;
		19'b1000011100110100010: color_data = Z;
		19'b1000011100110100011: color_data = Z;
		19'b1000011100110100100: color_data = Z;
		19'b1000011100110100101: color_data = Z;
		19'b1000011100110100110: color_data = Z;
		19'b1000011100110100111: color_data = Z;
		19'b1000011100110101000: color_data = Z;
		19'b1000011100110101001: color_data = Z;
		19'b1000011100110101010: color_data = Z;
		19'b1000011100110101011: color_data = Z;
		19'b1000011100110101100: color_data = Z;
		19'b1000011100110101101: color_data = Z;
		19'b1000011100110101110: color_data = Z;
		19'b1000011100110101111: color_data = Z;
		19'b1000011100110110000: color_data = Z;
		19'b1000011100110110001: color_data = Z;
		19'b1000011100110110010: color_data = Z;
		19'b1000011100110110011: color_data = Z;
		19'b1000011100110110100: color_data = Z;
		19'b1000011100110110101: color_data = Z;
		19'b1000011100110110110: color_data = Z;
		19'b1000011100110110111: color_data = Z;
		19'b1000011100110111000: color_data = Z;
		19'b1000011100110111001: color_data = Z;
		19'b1000011100110111010: color_data = Z;
		19'b1000011100110111011: color_data = Z;
		19'b1000011100110111100: color_data = Z;
		19'b1000011100110111101: color_data = Z;
		19'b1000011100111000110: color_data = Z;
		19'b1000011100111000111: color_data = Z;
		19'b1000011100111001000: color_data = Z;
		19'b1000011100111001001: color_data = Z;
		19'b1000011100111001010: color_data = Z;
		19'b1000011100111001011: color_data = Z;
		19'b1000011100111001100: color_data = Z;
		19'b1000011110010111110: color_data = Z;
		19'b1000011110010111111: color_data = Z;
		19'b1000011110011000000: color_data = Z;
		19'b1000011110011000001: color_data = Z;
		19'b1000011110011000010: color_data = Z;
		19'b1000011110011000011: color_data = Z;
		19'b1000011110011000100: color_data = Z;
		19'b1000011110011000101: color_data = Z;
		19'b1000011110011000110: color_data = Z;
		19'b1000011110011000111: color_data = Z;
		19'b1000011110011001000: color_data = Z;
		19'b1000011110011001001: color_data = Z;
		19'b1000011110011001010: color_data = Z;
		19'b1000011110011001011: color_data = Z;
		19'b1000011110011001100: color_data = Z;
		19'b1000011110011001101: color_data = Z;
		19'b1000011110011001110: color_data = Z;
		19'b1000011110011001111: color_data = Z;
		19'b1000011110011010000: color_data = Z;
		19'b1000011110011010001: color_data = Z;
		19'b1000011110011010010: color_data = Z;
		19'b1000011110011010011: color_data = Z;
		19'b1000011110011010100: color_data = Z;
		19'b1000011110011010101: color_data = Z;
		19'b1000011110011010110: color_data = Z;
		19'b1000011110011010111: color_data = Z;
		19'b1000011110011011000: color_data = Z;
		19'b1000011110011011001: color_data = Z;
		19'b1000011110011011010: color_data = Z;
		19'b1000011110011011011: color_data = Z;
		19'b1000011110011011100: color_data = Z;
		19'b1000011110011011101: color_data = Z;
		19'b1000011110011011110: color_data = Z;
		19'b1000011110011011111: color_data = Z;
		19'b1000011110011100000: color_data = Z;
		19'b1000011110011100001: color_data = Z;
		19'b1000011110011100010: color_data = Z;
		19'b1000011110011100011: color_data = Z;
		19'b1000011110011100100: color_data = Z;
		19'b1000011110011101110: color_data = Z;
		19'b1000011110011101111: color_data = Z;
		19'b1000011110011110000: color_data = Z;
		19'b1000011110011110001: color_data = Z;
		19'b1000011110011110010: color_data = Z;
		19'b1000011110011110011: color_data = Z;
		19'b1000011110011110100: color_data = Z;
		19'b1000011110011110101: color_data = Z;
		19'b1000011110011110110: color_data = Z;
		19'b1000011110011110111: color_data = Z;
		19'b1000011110011111000: color_data = Z;
		19'b1000011110011111001: color_data = Z;
		19'b1000011110011111010: color_data = Z;
		19'b1000011110011111011: color_data = Z;
		19'b1000011110011111100: color_data = Z;
		19'b1000011110011111101: color_data = Z;
		19'b1000011110011111110: color_data = Z;
		19'b1000011110011111111: color_data = Z;
		19'b1000011110100000000: color_data = Z;
		19'b1000011110100000001: color_data = Z;
		19'b1000011110100000010: color_data = Z;
		19'b1000011110100000011: color_data = Z;
		19'b1000011110100000100: color_data = Z;
		19'b1000011110100000101: color_data = Z;
		19'b1000011110100000110: color_data = Z;
		19'b1000011110100000111: color_data = Z;
		19'b1000011110100001000: color_data = Z;
		19'b1000011110100001001: color_data = Z;
		19'b1000011110100001010: color_data = Z;
		19'b1000011110100001011: color_data = Z;
		19'b1000011110100001100: color_data = Z;
		19'b1000011110100001101: color_data = Z;
		19'b1000011110100001110: color_data = Z;
		19'b1000011110100001111: color_data = Z;
		19'b1000011110100010000: color_data = Z;
		19'b1000011110100010001: color_data = Z;
		19'b1000011110100010010: color_data = Z;
		19'b1000011110100010011: color_data = Z;
		19'b1000011110100010100: color_data = Z;
		19'b1000011110100010101: color_data = Z;
		19'b1000011110100010110: color_data = Z;
		19'b1000011110100010111: color_data = Z;
		19'b1000011110100011000: color_data = Z;
		19'b1000011110100011001: color_data = Z;
		19'b1000011110100011010: color_data = Z;
		19'b1000011110100011011: color_data = Z;
		19'b1000011110100011100: color_data = Z;
		19'b1000011110100011101: color_data = Z;
		19'b1000011110100011110: color_data = Z;
		19'b1000011110100011111: color_data = Z;
		19'b1000011110100100000: color_data = Z;
		19'b1000011110100100001: color_data = Z;
		19'b1000011110100100010: color_data = Z;
		19'b1000011110100100011: color_data = Z;
		19'b1000011110100100100: color_data = Z;
		19'b1000011110100100101: color_data = Z;
		19'b1000011110100100110: color_data = Z;
		19'b1000011110100100111: color_data = Z;
		19'b1000011110100101000: color_data = Z;
		19'b1000011110100101001: color_data = Z;
		19'b1000011110100101111: color_data = Z;
		19'b1000011110100110000: color_data = Z;
		19'b1000011110100110001: color_data = Z;
		19'b1000011110101010100: color_data = Z;
		19'b1000011110101010101: color_data = Z;
		19'b1000011110101010110: color_data = Z;
		19'b1000011110101100110: color_data = Z;
		19'b1000011110101100111: color_data = Z;
		19'b1000011110101101000: color_data = Z;
		19'b1000011110101101001: color_data = Z;
		19'b1000011110101101010: color_data = Z;
		19'b1000011110101101011: color_data = Z;
		19'b1000011110101101100: color_data = Z;
		19'b1000011110101101101: color_data = Z;
		19'b1000011110101101110: color_data = Z;
		19'b1000011110101101111: color_data = Z;
		19'b1000011110101110000: color_data = Z;
		19'b1000011110101110001: color_data = Z;
		19'b1000011110101110010: color_data = Z;
		19'b1000011110101110011: color_data = Z;
		19'b1000011110101110100: color_data = Z;
		19'b1000011110101110101: color_data = Z;
		19'b1000011110101110110: color_data = Z;
		19'b1000011110101110111: color_data = Z;
		19'b1000011110101111000: color_data = Z;
		19'b1000011110101111001: color_data = Z;
		19'b1000011110101111010: color_data = Z;
		19'b1000011110101111011: color_data = Z;
		19'b1000011110101111100: color_data = Z;
		19'b1000011110101111101: color_data = Z;
		19'b1000011110101111110: color_data = Z;
		19'b1000011110101111111: color_data = Z;
		19'b1000011110110000000: color_data = Z;
		19'b1000011110110000001: color_data = Z;
		19'b1000011110110000010: color_data = Z;
		19'b1000011110110000011: color_data = Z;
		19'b1000011110110000100: color_data = Z;
		19'b1000011110110000101: color_data = Z;
		19'b1000011110110000110: color_data = Z;
		19'b1000011110110000111: color_data = Z;
		19'b1000011110110001000: color_data = Z;
		19'b1000011110110001001: color_data = Z;
		19'b1000011110110001010: color_data = Z;
		19'b1000011110110001011: color_data = Z;
		19'b1000011110110001100: color_data = Z;
		19'b1000011110110001101: color_data = Z;
		19'b1000011110110001110: color_data = Z;
		19'b1000011110110001111: color_data = Z;
		19'b1000011110110010000: color_data = Z;
		19'b1000011110110010001: color_data = Z;
		19'b1000011110110010010: color_data = Z;
		19'b1000011110110010011: color_data = Z;
		19'b1000011110110010100: color_data = Z;
		19'b1000011110110010101: color_data = Z;
		19'b1000011110110010110: color_data = Z;
		19'b1000011110110010111: color_data = Z;
		19'b1000011110110011000: color_data = Z;
		19'b1000011110110011001: color_data = Z;
		19'b1000011110110011010: color_data = Z;
		19'b1000011110110011011: color_data = Z;
		19'b1000011110110011100: color_data = Z;
		19'b1000011110110011101: color_data = Z;
		19'b1000011110110011110: color_data = Z;
		19'b1000011110110011111: color_data = Z;
		19'b1000011110110100000: color_data = Z;
		19'b1000011110110100001: color_data = Z;
		19'b1000011110110100010: color_data = Z;
		19'b1000011110110100011: color_data = Z;
		19'b1000011110110100100: color_data = Z;
		19'b1000011110110100101: color_data = Z;
		19'b1000011110110100110: color_data = Z;
		19'b1000011110110100111: color_data = Z;
		19'b1000011110110101000: color_data = Z;
		19'b1000011110110101001: color_data = Z;
		19'b1000011110110101010: color_data = Z;
		19'b1000011110110101011: color_data = Z;
		19'b1000011110110101100: color_data = Z;
		19'b1000011110110101101: color_data = Z;
		19'b1000011110110101110: color_data = Z;
		19'b1000011110110101111: color_data = Z;
		19'b1000011110110110000: color_data = Z;
		19'b1000011110110110001: color_data = Z;
		19'b1000011110110110010: color_data = Z;
		19'b1000011110110110011: color_data = Z;
		19'b1000011110110110100: color_data = Z;
		19'b1000011110110110101: color_data = Z;
		19'b1000011110110110110: color_data = Z;
		19'b1000011110110110111: color_data = Z;
		19'b1000011110110111000: color_data = Z;
		19'b1000011110110111001: color_data = Z;
		19'b1000011110110111010: color_data = Z;
		19'b1000011110110111011: color_data = Z;
		19'b1000011110110111100: color_data = Z;
		19'b1000011110110111101: color_data = Z;
		19'b1000011110111000110: color_data = Z;
		19'b1000011110111000111: color_data = Z;
		19'b1000011110111001000: color_data = Z;
		19'b1000011110111001001: color_data = Z;
		19'b1000011110111001010: color_data = Z;
		19'b1000011110111001011: color_data = Z;
		19'b1000011110111001100: color_data = Z;
		19'b1000100000010111110: color_data = Z;
		19'b1000100000010111111: color_data = Z;
		19'b1000100000011000000: color_data = Z;
		19'b1000100000011000001: color_data = Z;
		19'b1000100000011000010: color_data = Z;
		19'b1000100000011000011: color_data = Z;
		19'b1000100000011000100: color_data = Z;
		19'b1000100000011000101: color_data = Z;
		19'b1000100000011000110: color_data = Z;
		19'b1000100000011000111: color_data = Z;
		19'b1000100000011001000: color_data = Z;
		19'b1000100000011001001: color_data = Z;
		19'b1000100000011001010: color_data = Z;
		19'b1000100000011001011: color_data = Z;
		19'b1000100000011001100: color_data = Z;
		19'b1000100000011001101: color_data = Z;
		19'b1000100000011001110: color_data = Z;
		19'b1000100000011001111: color_data = Z;
		19'b1000100000011010000: color_data = Z;
		19'b1000100000011010001: color_data = Z;
		19'b1000100000011010010: color_data = Z;
		19'b1000100000011010011: color_data = Z;
		19'b1000100000011010100: color_data = Z;
		19'b1000100000011010101: color_data = Z;
		19'b1000100000011010110: color_data = Z;
		19'b1000100000011010111: color_data = Z;
		19'b1000100000011011000: color_data = Z;
		19'b1000100000011011001: color_data = Z;
		19'b1000100000011011010: color_data = Z;
		19'b1000100000011011011: color_data = Z;
		19'b1000100000011011100: color_data = Z;
		19'b1000100000011011101: color_data = Z;
		19'b1000100000011011110: color_data = Z;
		19'b1000100000011011111: color_data = Z;
		19'b1000100000011100000: color_data = Z;
		19'b1000100000011100001: color_data = Z;
		19'b1000100000011100010: color_data = Z;
		19'b1000100000011100011: color_data = Z;
		19'b1000100000011100100: color_data = Z;
		19'b1000100000011100101: color_data = Z;
		19'b1000100000011101100: color_data = Z;
		19'b1000100000011101101: color_data = Z;
		19'b1000100000011101110: color_data = Z;
		19'b1000100000011101111: color_data = Z;
		19'b1000100000011110000: color_data = Z;
		19'b1000100000011110001: color_data = Z;
		19'b1000100000011110010: color_data = Z;
		19'b1000100000011110011: color_data = Z;
		19'b1000100000011110100: color_data = Z;
		19'b1000100000011110101: color_data = Z;
		19'b1000100000011110110: color_data = Z;
		19'b1000100000011110111: color_data = Z;
		19'b1000100000011111000: color_data = Z;
		19'b1000100000011111001: color_data = Z;
		19'b1000100000011111010: color_data = Z;
		19'b1000100000011111011: color_data = Z;
		19'b1000100000011111100: color_data = Z;
		19'b1000100000011111101: color_data = Z;
		19'b1000100000011111110: color_data = Z;
		19'b1000100000011111111: color_data = Z;
		19'b1000100000100000000: color_data = Z;
		19'b1000100000100000001: color_data = Z;
		19'b1000100000100000010: color_data = Z;
		19'b1000100000100000011: color_data = Z;
		19'b1000100000100000100: color_data = Z;
		19'b1000100000100000101: color_data = Z;
		19'b1000100000100000110: color_data = Z;
		19'b1000100000100000111: color_data = Z;
		19'b1000100000100001000: color_data = Z;
		19'b1000100000100001001: color_data = Z;
		19'b1000100000100001010: color_data = Z;
		19'b1000100000100001011: color_data = Z;
		19'b1000100000100001100: color_data = Z;
		19'b1000100000100001101: color_data = Z;
		19'b1000100000100001110: color_data = Z;
		19'b1000100000100001111: color_data = Z;
		19'b1000100000100010000: color_data = Z;
		19'b1000100000100010001: color_data = Z;
		19'b1000100000100010010: color_data = Z;
		19'b1000100000100010011: color_data = Z;
		19'b1000100000100010100: color_data = Z;
		19'b1000100000100010101: color_data = Z;
		19'b1000100000100010110: color_data = Z;
		19'b1000100000100010111: color_data = Z;
		19'b1000100000100011000: color_data = Z;
		19'b1000100000100011001: color_data = Z;
		19'b1000100000100011010: color_data = Z;
		19'b1000100000100011011: color_data = Z;
		19'b1000100000100011100: color_data = Z;
		19'b1000100000100011101: color_data = Z;
		19'b1000100000100011110: color_data = Z;
		19'b1000100000100011111: color_data = Z;
		19'b1000100000100100000: color_data = Z;
		19'b1000100000100100001: color_data = Z;
		19'b1000100000100100010: color_data = Z;
		19'b1000100000100100011: color_data = Z;
		19'b1000100000100100100: color_data = Z;
		19'b1000100000100100101: color_data = Z;
		19'b1000100000100100110: color_data = Z;
		19'b1000100000100100111: color_data = Z;
		19'b1000100000100101000: color_data = Z;
		19'b1000100000100101001: color_data = Z;
		19'b1000100000100101111: color_data = Z;
		19'b1000100000100110000: color_data = Z;
		19'b1000100000100110001: color_data = Z;
		19'b1000100000100110010: color_data = Z;
		19'b1000100000101010100: color_data = Z;
		19'b1000100000101010101: color_data = Z;
		19'b1000100000101100101: color_data = Z;
		19'b1000100000101100110: color_data = Z;
		19'b1000100000101100111: color_data = Z;
		19'b1000100000101101000: color_data = Z;
		19'b1000100000101101001: color_data = Z;
		19'b1000100000101101010: color_data = Z;
		19'b1000100000101101011: color_data = Z;
		19'b1000100000101101100: color_data = Z;
		19'b1000100000101101101: color_data = Z;
		19'b1000100000101101110: color_data = Z;
		19'b1000100000101101111: color_data = Z;
		19'b1000100000101110000: color_data = Z;
		19'b1000100000101110001: color_data = Z;
		19'b1000100000101110010: color_data = Z;
		19'b1000100000101110011: color_data = Z;
		19'b1000100000101110100: color_data = Z;
		19'b1000100000101110101: color_data = Z;
		19'b1000100000101110110: color_data = Z;
		19'b1000100000101110111: color_data = Z;
		19'b1000100000101111000: color_data = Z;
		19'b1000100000101111001: color_data = Z;
		19'b1000100000101111010: color_data = Z;
		19'b1000100000101111011: color_data = Z;
		19'b1000100000101111100: color_data = Z;
		19'b1000100000101111101: color_data = Z;
		19'b1000100000101111110: color_data = Z;
		19'b1000100000101111111: color_data = Z;
		19'b1000100000110000000: color_data = Z;
		19'b1000100000110000001: color_data = Z;
		19'b1000100000110000010: color_data = Z;
		19'b1000100000110000011: color_data = Z;
		19'b1000100000110000100: color_data = Z;
		19'b1000100000110000101: color_data = Z;
		19'b1000100000110000110: color_data = Z;
		19'b1000100000110000111: color_data = Z;
		19'b1000100000110001000: color_data = Z;
		19'b1000100000110001001: color_data = Z;
		19'b1000100000110001010: color_data = Z;
		19'b1000100000110001011: color_data = Z;
		19'b1000100000110001100: color_data = Z;
		19'b1000100000110001101: color_data = Z;
		19'b1000100000110001110: color_data = Z;
		19'b1000100000110001111: color_data = Z;
		19'b1000100000110010000: color_data = Z;
		19'b1000100000110010001: color_data = Z;
		19'b1000100000110010010: color_data = Z;
		19'b1000100000110010011: color_data = Z;
		19'b1000100000110010100: color_data = Z;
		19'b1000100000110010101: color_data = Z;
		19'b1000100000110010110: color_data = Z;
		19'b1000100000110010111: color_data = Z;
		19'b1000100000110011000: color_data = Z;
		19'b1000100000110011001: color_data = Z;
		19'b1000100000110011010: color_data = Z;
		19'b1000100000110011011: color_data = Z;
		19'b1000100000110011100: color_data = Z;
		19'b1000100000110011101: color_data = Z;
		19'b1000100000110011110: color_data = Z;
		19'b1000100000110011111: color_data = Z;
		19'b1000100000110100000: color_data = Z;
		19'b1000100000110100001: color_data = Z;
		19'b1000100000110100010: color_data = Z;
		19'b1000100000110100011: color_data = Z;
		19'b1000100000110100100: color_data = Z;
		19'b1000100000110100101: color_data = Z;
		19'b1000100000110100110: color_data = Z;
		19'b1000100000110100111: color_data = Z;
		19'b1000100000110101000: color_data = Z;
		19'b1000100000110101001: color_data = Z;
		19'b1000100000110101010: color_data = Z;
		19'b1000100000110101011: color_data = Z;
		19'b1000100000110101100: color_data = Z;
		19'b1000100000110101101: color_data = Z;
		19'b1000100000110101110: color_data = Z;
		19'b1000100000110101111: color_data = Z;
		19'b1000100000110110000: color_data = Z;
		19'b1000100000110110001: color_data = Z;
		19'b1000100000110110010: color_data = Z;
		19'b1000100000110110011: color_data = Z;
		19'b1000100000110110100: color_data = Z;
		19'b1000100000110110101: color_data = Z;
		19'b1000100000110110110: color_data = Z;
		19'b1000100000110110111: color_data = Z;
		19'b1000100000110111000: color_data = Z;
		19'b1000100000110111001: color_data = Z;
		19'b1000100000110111010: color_data = Z;
		19'b1000100000110111011: color_data = Z;
		19'b1000100000110111100: color_data = Z;
		19'b1000100000110111101: color_data = Z;
		19'b1000100000111000111: color_data = Z;
		19'b1000100000111001000: color_data = Z;
		19'b1000100000111001001: color_data = Z;
		19'b1000100000111001010: color_data = Z;
		19'b1000100000111001011: color_data = Z;
		19'b1000100000111001100: color_data = Z;
		19'b1000100000111001101: color_data = Z;
		19'b1000100010010111111: color_data = Z;
		19'b1000100010011000000: color_data = Z;
		19'b1000100010011000001: color_data = Z;
		19'b1000100010011000010: color_data = Z;
		19'b1000100010011000011: color_data = Z;
		19'b1000100010011000100: color_data = Z;
		19'b1000100010011000101: color_data = Z;
		19'b1000100010011000110: color_data = Z;
		19'b1000100010011000111: color_data = Z;
		19'b1000100010011001000: color_data = Z;
		19'b1000100010011001001: color_data = Z;
		19'b1000100010011001010: color_data = Z;
		19'b1000100010011001011: color_data = Z;
		19'b1000100010011001100: color_data = Z;
		19'b1000100010011001101: color_data = Z;
		19'b1000100010011001110: color_data = Z;
		19'b1000100010011001111: color_data = Z;
		19'b1000100010011010000: color_data = Z;
		19'b1000100010011010001: color_data = Z;
		19'b1000100010011010010: color_data = Z;
		19'b1000100010011010011: color_data = Z;
		19'b1000100010011010100: color_data = Z;
		19'b1000100010011010101: color_data = Z;
		19'b1000100010011010110: color_data = Z;
		19'b1000100010011010111: color_data = Z;
		19'b1000100010011011000: color_data = Z;
		19'b1000100010011011001: color_data = Z;
		19'b1000100010011011010: color_data = Z;
		19'b1000100010011011011: color_data = Z;
		19'b1000100010011011100: color_data = Z;
		19'b1000100010011011101: color_data = Z;
		19'b1000100010011011110: color_data = Z;
		19'b1000100010011011111: color_data = Z;
		19'b1000100010011100000: color_data = Z;
		19'b1000100010011100001: color_data = Z;
		19'b1000100010011100010: color_data = Z;
		19'b1000100010011100011: color_data = Z;
		19'b1000100010011100100: color_data = Z;
		19'b1000100010011100101: color_data = Z;
		19'b1000100010011100110: color_data = Z;
		19'b1000100010011100111: color_data = Z;
		19'b1000100010011101000: color_data = Z;
		19'b1000100010011101001: color_data = Z;
		19'b1000100010011101010: color_data = Z;
		19'b1000100010011101011: color_data = Z;
		19'b1000100010011101100: color_data = Z;
		19'b1000100010011101101: color_data = Z;
		19'b1000100010011101110: color_data = Z;
		19'b1000100010011101111: color_data = Z;
		19'b1000100010011110000: color_data = Z;
		19'b1000100010011110001: color_data = Z;
		19'b1000100010011110010: color_data = Z;
		19'b1000100010011110011: color_data = Z;
		19'b1000100010011110100: color_data = Z;
		19'b1000100010011110101: color_data = Z;
		19'b1000100010011110110: color_data = Z;
		19'b1000100010011110111: color_data = Z;
		19'b1000100010011111000: color_data = Z;
		19'b1000100010011111001: color_data = Z;
		19'b1000100010011111010: color_data = Z;
		19'b1000100010011111011: color_data = Z;
		19'b1000100010011111100: color_data = Z;
		19'b1000100010011111101: color_data = Z;
		19'b1000100010011111110: color_data = Z;
		19'b1000100010011111111: color_data = Z;
		19'b1000100010100000000: color_data = Z;
		19'b1000100010100000001: color_data = Z;
		19'b1000100010100000010: color_data = Z;
		19'b1000100010100000011: color_data = Z;
		19'b1000100010100000100: color_data = Z;
		19'b1000100010100000101: color_data = Z;
		19'b1000100010100000110: color_data = Z;
		19'b1000100010100000111: color_data = Z;
		19'b1000100010100001000: color_data = Z;
		19'b1000100010100001001: color_data = Z;
		19'b1000100010100001010: color_data = Z;
		19'b1000100010100001011: color_data = Z;
		19'b1000100010100001100: color_data = Z;
		19'b1000100010100001101: color_data = Z;
		19'b1000100010100001110: color_data = Z;
		19'b1000100010100001111: color_data = Z;
		19'b1000100010100010000: color_data = Z;
		19'b1000100010100010001: color_data = Z;
		19'b1000100010100010010: color_data = Z;
		19'b1000100010100010011: color_data = Z;
		19'b1000100010100010100: color_data = Z;
		19'b1000100010100010101: color_data = Z;
		19'b1000100010100010110: color_data = Z;
		19'b1000100010100010111: color_data = Z;
		19'b1000100010100011000: color_data = Z;
		19'b1000100010100011001: color_data = Z;
		19'b1000100010100011010: color_data = Z;
		19'b1000100010100011011: color_data = Z;
		19'b1000100010100011100: color_data = Z;
		19'b1000100010100011101: color_data = Z;
		19'b1000100010100011110: color_data = Z;
		19'b1000100010100011111: color_data = Z;
		19'b1000100010100100000: color_data = Z;
		19'b1000100010100100001: color_data = Z;
		19'b1000100010100100010: color_data = Z;
		19'b1000100010100100011: color_data = Z;
		19'b1000100010100100100: color_data = Z;
		19'b1000100010100100101: color_data = Z;
		19'b1000100010100100110: color_data = Z;
		19'b1000100010100100111: color_data = Z;
		19'b1000100010100101000: color_data = Z;
		19'b1000100010100101001: color_data = Z;
		19'b1000100010100101010: color_data = Z;
		19'b1000100010100101111: color_data = Z;
		19'b1000100010100110000: color_data = Z;
		19'b1000100010100110001: color_data = Z;
		19'b1000100010100110010: color_data = Z;
		19'b1000100010100110011: color_data = Z;
		19'b1000100010101100011: color_data = Z;
		19'b1000100010101100100: color_data = Z;
		19'b1000100010101100101: color_data = Z;
		19'b1000100010101100110: color_data = Z;
		19'b1000100010101100111: color_data = Z;
		19'b1000100010101101000: color_data = Z;
		19'b1000100010101101001: color_data = Z;
		19'b1000100010101101010: color_data = Z;
		19'b1000100010101101011: color_data = Z;
		19'b1000100010101101100: color_data = Z;
		19'b1000100010101101101: color_data = Z;
		19'b1000100010101101110: color_data = Z;
		19'b1000100010101101111: color_data = Z;
		19'b1000100010101110000: color_data = Z;
		19'b1000100010101110001: color_data = Z;
		19'b1000100010101110010: color_data = Z;
		19'b1000100010101110011: color_data = Z;
		19'b1000100010101110100: color_data = Z;
		19'b1000100010101110101: color_data = Z;
		19'b1000100010101110110: color_data = Z;
		19'b1000100010101110111: color_data = Z;
		19'b1000100010101111000: color_data = Z;
		19'b1000100010101111001: color_data = Z;
		19'b1000100010101111010: color_data = Z;
		19'b1000100010101111011: color_data = Z;
		19'b1000100010101111100: color_data = Z;
		19'b1000100010101111101: color_data = Z;
		19'b1000100010101111110: color_data = Z;
		19'b1000100010101111111: color_data = Z;
		19'b1000100010110000000: color_data = Z;
		19'b1000100010110000001: color_data = Z;
		19'b1000100010110000010: color_data = Z;
		19'b1000100010110000011: color_data = Z;
		19'b1000100010110000100: color_data = Z;
		19'b1000100010110000101: color_data = Z;
		19'b1000100010110000110: color_data = Z;
		19'b1000100010110000111: color_data = Z;
		19'b1000100010110001000: color_data = Z;
		19'b1000100010110001001: color_data = Z;
		19'b1000100010110001010: color_data = Z;
		19'b1000100010110001011: color_data = Z;
		19'b1000100010110001100: color_data = Z;
		19'b1000100010110001101: color_data = Z;
		19'b1000100010110001110: color_data = Z;
		19'b1000100010110001111: color_data = Z;
		19'b1000100010110010000: color_data = Z;
		19'b1000100010110010001: color_data = Z;
		19'b1000100010110010010: color_data = Z;
		19'b1000100010110010011: color_data = Z;
		19'b1000100010110010100: color_data = Z;
		19'b1000100010110010101: color_data = Z;
		19'b1000100010110010110: color_data = Z;
		19'b1000100010110010111: color_data = Z;
		19'b1000100010110011000: color_data = Z;
		19'b1000100010110011001: color_data = Z;
		19'b1000100010110011010: color_data = Z;
		19'b1000100010110011011: color_data = Z;
		19'b1000100010110011100: color_data = Z;
		19'b1000100010110011101: color_data = Z;
		19'b1000100010110011110: color_data = Z;
		19'b1000100010110011111: color_data = Z;
		19'b1000100010110100000: color_data = Z;
		19'b1000100010110100001: color_data = Z;
		19'b1000100010110100010: color_data = Z;
		19'b1000100010110100011: color_data = Z;
		19'b1000100010110100100: color_data = Z;
		19'b1000100010110100101: color_data = Z;
		19'b1000100010110100110: color_data = Z;
		19'b1000100010110100111: color_data = Z;
		19'b1000100010110101000: color_data = Z;
		19'b1000100010110101001: color_data = Z;
		19'b1000100010110101010: color_data = Z;
		19'b1000100010110101011: color_data = Z;
		19'b1000100010110101100: color_data = Z;
		19'b1000100010110101101: color_data = Z;
		19'b1000100010110101110: color_data = Z;
		19'b1000100010110101111: color_data = Z;
		19'b1000100010110110000: color_data = Z;
		19'b1000100010110110001: color_data = Z;
		19'b1000100010110110010: color_data = Z;
		19'b1000100010110110011: color_data = Z;
		19'b1000100010110110100: color_data = Z;
		19'b1000100010110110101: color_data = Z;
		19'b1000100010110110110: color_data = Z;
		19'b1000100010110110111: color_data = Z;
		19'b1000100010110111000: color_data = Z;
		19'b1000100010110111001: color_data = Z;
		19'b1000100010110111010: color_data = Z;
		19'b1000100010110111011: color_data = Z;
		19'b1000100010110111100: color_data = Z;
		19'b1000100010110111101: color_data = Z;
		19'b1000100010111000111: color_data = Z;
		19'b1000100010111001000: color_data = Z;
		19'b1000100010111001001: color_data = Z;
		19'b1000100010111001010: color_data = Z;
		19'b1000100010111001011: color_data = Z;
		19'b1000100010111001100: color_data = Z;
		19'b1000100010111001101: color_data = Z;
		19'b1000100100011000000: color_data = Z;
		19'b1000100100011000001: color_data = Z;
		19'b1000100100011000010: color_data = Z;
		19'b1000100100011000011: color_data = Z;
		19'b1000100100011000100: color_data = Z;
		19'b1000100100011000101: color_data = Z;
		19'b1000100100011000110: color_data = Z;
		19'b1000100100011000111: color_data = Z;
		19'b1000100100011001000: color_data = Z;
		19'b1000100100011001001: color_data = Z;
		19'b1000100100011001010: color_data = Z;
		19'b1000100100011001011: color_data = Z;
		19'b1000100100011001100: color_data = Z;
		19'b1000100100011001101: color_data = Z;
		19'b1000100100011001110: color_data = Z;
		19'b1000100100011001111: color_data = Z;
		19'b1000100100011010000: color_data = Z;
		19'b1000100100011010001: color_data = Z;
		19'b1000100100011010010: color_data = Z;
		19'b1000100100011010011: color_data = Z;
		19'b1000100100011010100: color_data = Z;
		19'b1000100100011010101: color_data = Z;
		19'b1000100100011010110: color_data = Z;
		19'b1000100100011010111: color_data = Z;
		19'b1000100100011011000: color_data = Z;
		19'b1000100100011011001: color_data = Z;
		19'b1000100100011011010: color_data = Z;
		19'b1000100100011011011: color_data = Z;
		19'b1000100100011011100: color_data = Z;
		19'b1000100100011011101: color_data = Z;
		19'b1000100100011011110: color_data = Z;
		19'b1000100100011011111: color_data = Z;
		19'b1000100100011100000: color_data = Z;
		19'b1000100100011100001: color_data = Z;
		19'b1000100100011100010: color_data = Z;
		19'b1000100100011100011: color_data = Z;
		19'b1000100100011100100: color_data = Z;
		19'b1000100100011100101: color_data = Z;
		19'b1000100100011100110: color_data = Z;
		19'b1000100100011100111: color_data = Z;
		19'b1000100100011101000: color_data = Z;
		19'b1000100100011101001: color_data = Z;
		19'b1000100100011101010: color_data = Z;
		19'b1000100100011101011: color_data = Z;
		19'b1000100100011101100: color_data = Z;
		19'b1000100100011101101: color_data = Z;
		19'b1000100100011101110: color_data = Z;
		19'b1000100100011101111: color_data = Z;
		19'b1000100100011110000: color_data = Z;
		19'b1000100100011110001: color_data = Z;
		19'b1000100100011110010: color_data = Z;
		19'b1000100100011110011: color_data = Z;
		19'b1000100100011110100: color_data = Z;
		19'b1000100100011110101: color_data = Z;
		19'b1000100100011110110: color_data = Z;
		19'b1000100100011110111: color_data = Z;
		19'b1000100100011111000: color_data = Z;
		19'b1000100100011111001: color_data = Z;
		19'b1000100100011111010: color_data = Z;
		19'b1000100100011111011: color_data = Z;
		19'b1000100100011111100: color_data = Z;
		19'b1000100100011111101: color_data = Z;
		19'b1000100100011111110: color_data = Z;
		19'b1000100100011111111: color_data = Z;
		19'b1000100100100000000: color_data = Z;
		19'b1000100100100000001: color_data = Z;
		19'b1000100100100000010: color_data = Z;
		19'b1000100100100000011: color_data = Z;
		19'b1000100100100000100: color_data = Z;
		19'b1000100100100000101: color_data = Z;
		19'b1000100100100000110: color_data = Z;
		19'b1000100100100000111: color_data = Z;
		19'b1000100100100001000: color_data = Z;
		19'b1000100100100001001: color_data = Z;
		19'b1000100100100001010: color_data = Z;
		19'b1000100100100001011: color_data = Z;
		19'b1000100100100001100: color_data = Z;
		19'b1000100100100001101: color_data = Z;
		19'b1000100100100001110: color_data = Z;
		19'b1000100100100001111: color_data = Z;
		19'b1000100100100010000: color_data = Z;
		19'b1000100100100010001: color_data = Z;
		19'b1000100100100010010: color_data = Z;
		19'b1000100100100010011: color_data = Z;
		19'b1000100100100010100: color_data = Z;
		19'b1000100100100010101: color_data = Z;
		19'b1000100100100010110: color_data = Z;
		19'b1000100100100010111: color_data = Z;
		19'b1000100100100011000: color_data = Z;
		19'b1000100100100011001: color_data = Z;
		19'b1000100100100011010: color_data = Z;
		19'b1000100100100011011: color_data = Z;
		19'b1000100100100011100: color_data = Z;
		19'b1000100100100011101: color_data = Z;
		19'b1000100100100100000: color_data = Z;
		19'b1000100100100100100: color_data = Z;
		19'b1000100100100100101: color_data = Z;
		19'b1000100100100100110: color_data = Z;
		19'b1000100100100100111: color_data = Z;
		19'b1000100100100101000: color_data = Z;
		19'b1000100100100101001: color_data = Z;
		19'b1000100100100101010: color_data = Z;
		19'b1000100100100101111: color_data = Z;
		19'b1000100100100110000: color_data = Z;
		19'b1000100100100110001: color_data = Z;
		19'b1000100100100110010: color_data = Z;
		19'b1000100100100110011: color_data = Z;
		19'b1000100100100110100: color_data = Z;
		19'b1000100100100110101: color_data = Z;
		19'b1000100100100110110: color_data = Z;
		19'b1000100100101011100: color_data = Z;
		19'b1000100100101100010: color_data = Z;
		19'b1000100100101100011: color_data = Z;
		19'b1000100100101100100: color_data = Z;
		19'b1000100100101100101: color_data = Z;
		19'b1000100100101100110: color_data = Z;
		19'b1000100100101100111: color_data = Z;
		19'b1000100100101101000: color_data = Z;
		19'b1000100100101101001: color_data = Z;
		19'b1000100100101101010: color_data = Z;
		19'b1000100100101101011: color_data = Z;
		19'b1000100100101101100: color_data = Z;
		19'b1000100100101101101: color_data = Z;
		19'b1000100100101101110: color_data = Z;
		19'b1000100100101101111: color_data = Z;
		19'b1000100100101110000: color_data = Z;
		19'b1000100100101110001: color_data = Z;
		19'b1000100100101110010: color_data = Z;
		19'b1000100100101110011: color_data = Z;
		19'b1000100100101110100: color_data = Z;
		19'b1000100100101110101: color_data = Z;
		19'b1000100100101110110: color_data = Z;
		19'b1000100100101110111: color_data = Z;
		19'b1000100100101111000: color_data = Z;
		19'b1000100100101111001: color_data = Z;
		19'b1000100100101111010: color_data = Z;
		19'b1000100100101111011: color_data = Z;
		19'b1000100100101111100: color_data = Z;
		19'b1000100100101111101: color_data = Z;
		19'b1000100100101111110: color_data = Z;
		19'b1000100100101111111: color_data = Z;
		19'b1000100100110000000: color_data = Z;
		19'b1000100100110000001: color_data = Z;
		19'b1000100100110000010: color_data = Z;
		19'b1000100100110000011: color_data = Z;
		19'b1000100100110000100: color_data = Z;
		19'b1000100100110000101: color_data = Z;
		19'b1000100100110000110: color_data = Z;
		19'b1000100100110000111: color_data = Z;
		19'b1000100100110001000: color_data = Z;
		19'b1000100100110001001: color_data = Z;
		19'b1000100100110001010: color_data = Z;
		19'b1000100100110001011: color_data = Z;
		19'b1000100100110001100: color_data = Z;
		19'b1000100100110001101: color_data = Z;
		19'b1000100100110001110: color_data = Z;
		19'b1000100100110001111: color_data = Z;
		19'b1000100100110010000: color_data = Z;
		19'b1000100100110010001: color_data = Z;
		19'b1000100100110010010: color_data = Z;
		19'b1000100100110010011: color_data = Z;
		19'b1000100100110010100: color_data = Z;
		19'b1000100100110010101: color_data = Z;
		19'b1000100100110010110: color_data = Z;
		19'b1000100100110010111: color_data = Z;
		19'b1000100100110011000: color_data = Z;
		19'b1000100100110011001: color_data = Z;
		19'b1000100100110011010: color_data = Z;
		19'b1000100100110011011: color_data = Z;
		19'b1000100100110011100: color_data = Z;
		19'b1000100100110011101: color_data = Z;
		19'b1000100100110011110: color_data = Z;
		19'b1000100100110011111: color_data = Z;
		19'b1000100100110100000: color_data = Z;
		19'b1000100100110100001: color_data = Z;
		19'b1000100100110100010: color_data = Z;
		19'b1000100100110100011: color_data = Z;
		19'b1000100100110100100: color_data = Z;
		19'b1000100100110100101: color_data = Z;
		19'b1000100100110100110: color_data = Z;
		19'b1000100100110100111: color_data = Z;
		19'b1000100100110101000: color_data = Z;
		19'b1000100100110101001: color_data = Z;
		19'b1000100100110101010: color_data = Z;
		19'b1000100100110101011: color_data = Z;
		19'b1000100100110101100: color_data = Z;
		19'b1000100100110101101: color_data = Z;
		19'b1000100100110101110: color_data = Z;
		19'b1000100100110101111: color_data = Z;
		19'b1000100100110110000: color_data = Z;
		19'b1000100100110110001: color_data = Z;
		19'b1000100100110110010: color_data = Z;
		19'b1000100100110110011: color_data = Z;
		19'b1000100100110110100: color_data = Z;
		19'b1000100100110110101: color_data = Z;
		19'b1000100100110110110: color_data = Z;
		19'b1000100100110110111: color_data = Z;
		19'b1000100100110111000: color_data = Z;
		19'b1000100100110111001: color_data = Z;
		19'b1000100100110111010: color_data = Z;
		19'b1000100100110111011: color_data = Z;
		19'b1000100100110111100: color_data = Z;
		19'b1000100100110111101: color_data = Z;
		19'b1000100100111000111: color_data = Z;
		19'b1000100100111001000: color_data = Z;
		19'b1000100100111001001: color_data = Z;
		19'b1000100100111001010: color_data = Z;
		19'b1000100100111001011: color_data = Z;
		19'b1000100100111001100: color_data = Z;
		19'b1000100100111001101: color_data = Z;
		19'b1000100110011000001: color_data = Z;
		19'b1000100110011000010: color_data = Z;
		19'b1000100110011000011: color_data = Z;
		19'b1000100110011000100: color_data = Z;
		19'b1000100110011000101: color_data = Z;
		19'b1000100110011000110: color_data = Z;
		19'b1000100110011000111: color_data = Z;
		19'b1000100110011001000: color_data = Z;
		19'b1000100110011001001: color_data = Z;
		19'b1000100110011001010: color_data = Z;
		19'b1000100110011001011: color_data = Z;
		19'b1000100110011001100: color_data = Z;
		19'b1000100110011001101: color_data = Z;
		19'b1000100110011001110: color_data = Z;
		19'b1000100110011001111: color_data = Z;
		19'b1000100110011010000: color_data = Z;
		19'b1000100110011010001: color_data = Z;
		19'b1000100110011010010: color_data = Z;
		19'b1000100110011010011: color_data = Z;
		19'b1000100110011010100: color_data = Z;
		19'b1000100110011010101: color_data = Z;
		19'b1000100110011010110: color_data = Z;
		19'b1000100110011010111: color_data = Z;
		19'b1000100110011011000: color_data = Z;
		19'b1000100110011011001: color_data = Z;
		19'b1000100110011011010: color_data = Z;
		19'b1000100110011011011: color_data = Z;
		19'b1000100110011011100: color_data = Z;
		19'b1000100110011011101: color_data = Z;
		19'b1000100110011011110: color_data = Z;
		19'b1000100110011011111: color_data = Z;
		19'b1000100110011100000: color_data = Z;
		19'b1000100110011100001: color_data = Z;
		19'b1000100110011100010: color_data = Z;
		19'b1000100110011100011: color_data = Z;
		19'b1000100110011100100: color_data = Z;
		19'b1000100110011100101: color_data = Z;
		19'b1000100110011100110: color_data = Z;
		19'b1000100110011100111: color_data = Z;
		19'b1000100110011101000: color_data = Z;
		19'b1000100110011101001: color_data = Z;
		19'b1000100110011101010: color_data = Z;
		19'b1000100110011101011: color_data = Z;
		19'b1000100110011101100: color_data = Z;
		19'b1000100110011101101: color_data = Z;
		19'b1000100110011101110: color_data = Z;
		19'b1000100110011101111: color_data = Z;
		19'b1000100110011110000: color_data = Z;
		19'b1000100110011110001: color_data = Z;
		19'b1000100110011110010: color_data = Z;
		19'b1000100110011110011: color_data = Z;
		19'b1000100110011110100: color_data = Z;
		19'b1000100110011110101: color_data = Z;
		19'b1000100110011110110: color_data = Z;
		19'b1000100110011110111: color_data = Z;
		19'b1000100110011111000: color_data = Z;
		19'b1000100110011111001: color_data = Z;
		19'b1000100110011111010: color_data = Z;
		19'b1000100110011111011: color_data = Z;
		19'b1000100110011111100: color_data = Z;
		19'b1000100110011111101: color_data = Z;
		19'b1000100110011111110: color_data = Z;
		19'b1000100110011111111: color_data = Z;
		19'b1000100110100000000: color_data = Z;
		19'b1000100110100000001: color_data = Z;
		19'b1000100110100000010: color_data = Z;
		19'b1000100110100000011: color_data = Z;
		19'b1000100110100000100: color_data = Z;
		19'b1000100110100000101: color_data = Z;
		19'b1000100110100000110: color_data = Z;
		19'b1000100110100000111: color_data = Z;
		19'b1000100110100001000: color_data = Z;
		19'b1000100110100001001: color_data = Z;
		19'b1000100110100001010: color_data = Z;
		19'b1000100110100001011: color_data = Z;
		19'b1000100110100001100: color_data = Z;
		19'b1000100110100001101: color_data = Z;
		19'b1000100110100001110: color_data = Z;
		19'b1000100110100001111: color_data = Z;
		19'b1000100110100010000: color_data = Z;
		19'b1000100110100010001: color_data = Z;
		19'b1000100110100010010: color_data = Z;
		19'b1000100110100010011: color_data = Z;
		19'b1000100110100010100: color_data = Z;
		19'b1000100110100010101: color_data = Z;
		19'b1000100110100010110: color_data = Z;
		19'b1000100110100010111: color_data = Z;
		19'b1000100110100011000: color_data = Z;
		19'b1000100110100011001: color_data = Z;
		19'b1000100110100011010: color_data = Z;
		19'b1000100110100011011: color_data = Z;
		19'b1000100110100011100: color_data = Z;
		19'b1000100110100100100: color_data = Z;
		19'b1000100110100100101: color_data = Z;
		19'b1000100110100100110: color_data = Z;
		19'b1000100110100100111: color_data = Z;
		19'b1000100110100101000: color_data = Z;
		19'b1000100110100101001: color_data = Z;
		19'b1000100110100101111: color_data = Z;
		19'b1000100110100110000: color_data = Z;
		19'b1000100110100110001: color_data = Z;
		19'b1000100110100110010: color_data = Z;
		19'b1000100110100110011: color_data = Z;
		19'b1000100110100110100: color_data = Z;
		19'b1000100110100110101: color_data = Z;
		19'b1000100110100110110: color_data = Z;
		19'b1000100110100110111: color_data = Z;
		19'b1000100110100111000: color_data = Z;
		19'b1000100110100111100: color_data = Z;
		19'b1000100110100111101: color_data = Z;
		19'b1000100110100111110: color_data = Z;
		19'b1000100110100111111: color_data = Z;
		19'b1000100110101011100: color_data = Z;
		19'b1000100110101100001: color_data = Z;
		19'b1000100110101100010: color_data = Z;
		19'b1000100110101100011: color_data = Z;
		19'b1000100110101100100: color_data = Z;
		19'b1000100110101100101: color_data = Z;
		19'b1000100110101100110: color_data = Z;
		19'b1000100110101100111: color_data = Z;
		19'b1000100110101101000: color_data = Z;
		19'b1000100110101101001: color_data = Z;
		19'b1000100110101101010: color_data = Z;
		19'b1000100110101101011: color_data = Z;
		19'b1000100110101101100: color_data = Z;
		19'b1000100110101101101: color_data = Z;
		19'b1000100110101101110: color_data = Z;
		19'b1000100110101101111: color_data = Z;
		19'b1000100110101110000: color_data = Z;
		19'b1000100110101110001: color_data = Z;
		19'b1000100110101110010: color_data = Z;
		19'b1000100110101110011: color_data = Z;
		19'b1000100110101110100: color_data = Z;
		19'b1000100110101110101: color_data = Z;
		19'b1000100110101110110: color_data = Z;
		19'b1000100110101110111: color_data = Z;
		19'b1000100110101111000: color_data = Z;
		19'b1000100110101111001: color_data = Z;
		19'b1000100110101111010: color_data = Z;
		19'b1000100110101111011: color_data = Z;
		19'b1000100110101111100: color_data = Z;
		19'b1000100110101111101: color_data = Z;
		19'b1000100110101111110: color_data = Z;
		19'b1000100110101111111: color_data = Z;
		19'b1000100110110000000: color_data = Z;
		19'b1000100110110000001: color_data = Z;
		19'b1000100110110000010: color_data = Z;
		19'b1000100110110000011: color_data = Z;
		19'b1000100110110000100: color_data = Z;
		19'b1000100110110000101: color_data = Z;
		19'b1000100110110000110: color_data = Z;
		19'b1000100110110000111: color_data = Z;
		19'b1000100110110001000: color_data = Z;
		19'b1000100110110001001: color_data = Z;
		19'b1000100110110001010: color_data = Z;
		19'b1000100110110001011: color_data = Z;
		19'b1000100110110001100: color_data = Z;
		19'b1000100110110001101: color_data = Z;
		19'b1000100110110001110: color_data = Z;
		19'b1000100110110001111: color_data = Z;
		19'b1000100110110010000: color_data = Z;
		19'b1000100110110010001: color_data = Z;
		19'b1000100110110010010: color_data = Z;
		19'b1000100110110010011: color_data = Z;
		19'b1000100110110010100: color_data = Z;
		19'b1000100110110010101: color_data = Z;
		19'b1000100110110010110: color_data = Z;
		19'b1000100110110010111: color_data = Z;
		19'b1000100110110011000: color_data = Z;
		19'b1000100110110011001: color_data = Z;
		19'b1000100110110011010: color_data = Z;
		19'b1000100110110011011: color_data = Z;
		19'b1000100110110011100: color_data = Z;
		19'b1000100110110011101: color_data = Z;
		19'b1000100110110011110: color_data = Z;
		19'b1000100110110011111: color_data = Z;
		19'b1000100110110100000: color_data = Z;
		19'b1000100110110100001: color_data = Z;
		19'b1000100110110100010: color_data = Z;
		19'b1000100110110100011: color_data = Z;
		19'b1000100110110100100: color_data = Z;
		19'b1000100110110100101: color_data = Z;
		19'b1000100110110100110: color_data = Z;
		19'b1000100110110100111: color_data = Z;
		19'b1000100110110101000: color_data = Z;
		19'b1000100110110101001: color_data = Z;
		19'b1000100110110101010: color_data = Z;
		19'b1000100110110101011: color_data = Z;
		19'b1000100110110101100: color_data = Z;
		19'b1000100110110101101: color_data = Z;
		19'b1000100110110101110: color_data = Z;
		19'b1000100110110101111: color_data = Z;
		19'b1000100110110110000: color_data = Z;
		19'b1000100110110110001: color_data = Z;
		19'b1000100110110110010: color_data = Z;
		19'b1000100110110110011: color_data = Z;
		19'b1000100110110110100: color_data = Z;
		19'b1000100110110110101: color_data = Z;
		19'b1000100110110110110: color_data = Z;
		19'b1000100110110110111: color_data = Z;
		19'b1000100110110111000: color_data = Z;
		19'b1000100110110111001: color_data = Z;
		19'b1000100110110111010: color_data = Z;
		19'b1000100110110111011: color_data = Z;
		19'b1000100110110111100: color_data = Z;
		19'b1000100110110111101: color_data = Z;
		19'b1000100110111000111: color_data = Z;
		19'b1000100110111001000: color_data = Z;
		19'b1000100110111001001: color_data = Z;
		19'b1000100110111001010: color_data = Z;
		19'b1000100110111001011: color_data = Z;
		19'b1000100110111001100: color_data = Z;
		19'b1000100110111001101: color_data = Z;
		19'b1000101000011000010: color_data = Z;
		19'b1000101000011000011: color_data = Z;
		19'b1000101000011000100: color_data = Z;
		19'b1000101000011000101: color_data = Z;
		19'b1000101000011000110: color_data = Z;
		19'b1000101000011000111: color_data = Z;
		19'b1000101000011001000: color_data = Z;
		19'b1000101000011001001: color_data = Z;
		19'b1000101000011001010: color_data = Z;
		19'b1000101000011001011: color_data = Z;
		19'b1000101000011001100: color_data = Z;
		19'b1000101000011001101: color_data = Z;
		19'b1000101000011001110: color_data = Z;
		19'b1000101000011001111: color_data = Z;
		19'b1000101000011010000: color_data = Z;
		19'b1000101000011010001: color_data = Z;
		19'b1000101000011010010: color_data = Z;
		19'b1000101000011010011: color_data = Z;
		19'b1000101000011010100: color_data = Z;
		19'b1000101000011010101: color_data = Z;
		19'b1000101000011010110: color_data = Z;
		19'b1000101000011010111: color_data = Z;
		19'b1000101000011011000: color_data = Z;
		19'b1000101000011011001: color_data = Z;
		19'b1000101000011011010: color_data = Z;
		19'b1000101000011011011: color_data = Z;
		19'b1000101000011011100: color_data = Z;
		19'b1000101000011011101: color_data = Z;
		19'b1000101000011011110: color_data = Z;
		19'b1000101000011011111: color_data = Z;
		19'b1000101000011100000: color_data = Z;
		19'b1000101000011100001: color_data = Z;
		19'b1000101000011100010: color_data = Z;
		19'b1000101000011100011: color_data = Z;
		19'b1000101000011100100: color_data = Z;
		19'b1000101000011100101: color_data = Z;
		19'b1000101000011100110: color_data = Z;
		19'b1000101000011100111: color_data = Z;
		19'b1000101000011101000: color_data = Z;
		19'b1000101000011101001: color_data = Z;
		19'b1000101000011101010: color_data = Z;
		19'b1000101000011101011: color_data = Z;
		19'b1000101000011101100: color_data = Z;
		19'b1000101000011101101: color_data = Z;
		19'b1000101000011101110: color_data = Z;
		19'b1000101000011101111: color_data = Z;
		19'b1000101000011110000: color_data = Z;
		19'b1000101000011110001: color_data = Z;
		19'b1000101000011110010: color_data = Z;
		19'b1000101000011110011: color_data = Z;
		19'b1000101000011110100: color_data = Z;
		19'b1000101000011110101: color_data = Z;
		19'b1000101000011110110: color_data = Z;
		19'b1000101000011110111: color_data = Z;
		19'b1000101000011111000: color_data = Z;
		19'b1000101000011111001: color_data = Z;
		19'b1000101000011111010: color_data = Z;
		19'b1000101000011111011: color_data = Z;
		19'b1000101000011111100: color_data = Z;
		19'b1000101000011111101: color_data = Z;
		19'b1000101000011111110: color_data = Z;
		19'b1000101000011111111: color_data = Z;
		19'b1000101000100000000: color_data = Z;
		19'b1000101000100000001: color_data = Z;
		19'b1000101000100000010: color_data = Z;
		19'b1000101000100000011: color_data = Z;
		19'b1000101000100000100: color_data = Z;
		19'b1000101000100000101: color_data = Z;
		19'b1000101000100000110: color_data = Z;
		19'b1000101000100000111: color_data = Z;
		19'b1000101000100001000: color_data = Z;
		19'b1000101000100001001: color_data = Z;
		19'b1000101000100001010: color_data = Z;
		19'b1000101000100001011: color_data = Z;
		19'b1000101000100001100: color_data = Z;
		19'b1000101000100001101: color_data = Z;
		19'b1000101000100001110: color_data = Z;
		19'b1000101000100001111: color_data = Z;
		19'b1000101000100010000: color_data = Z;
		19'b1000101000100010001: color_data = Z;
		19'b1000101000100010010: color_data = Z;
		19'b1000101000100010011: color_data = Z;
		19'b1000101000100010100: color_data = Z;
		19'b1000101000100010101: color_data = Z;
		19'b1000101000100010110: color_data = Z;
		19'b1000101000100010111: color_data = Z;
		19'b1000101000100011000: color_data = Z;
		19'b1000101000100100100: color_data = Z;
		19'b1000101000100100101: color_data = Z;
		19'b1000101000100100110: color_data = Z;
		19'b1000101000100100111: color_data = Z;
		19'b1000101000100101000: color_data = Z;
		19'b1000101000100101100: color_data = Z;
		19'b1000101000100101101: color_data = Z;
		19'b1000101000100101110: color_data = Z;
		19'b1000101000100101111: color_data = Z;
		19'b1000101000100110000: color_data = Z;
		19'b1000101000100110001: color_data = Z;
		19'b1000101000100110010: color_data = Z;
		19'b1000101000100110011: color_data = Z;
		19'b1000101000100110100: color_data = Z;
		19'b1000101000100110101: color_data = Z;
		19'b1000101000100110110: color_data = Z;
		19'b1000101000100110111: color_data = Z;
		19'b1000101000100111000: color_data = Z;
		19'b1000101000100111001: color_data = Z;
		19'b1000101000100111010: color_data = Z;
		19'b1000101000100111011: color_data = Z;
		19'b1000101000100111100: color_data = Z;
		19'b1000101000100111101: color_data = Z;
		19'b1000101000100111110: color_data = Z;
		19'b1000101000100111111: color_data = Z;
		19'b1000101000101000000: color_data = Z;
		19'b1000101000101100000: color_data = Z;
		19'b1000101000101100001: color_data = Z;
		19'b1000101000101100010: color_data = Z;
		19'b1000101000101100011: color_data = Z;
		19'b1000101000101100100: color_data = Z;
		19'b1000101000101100101: color_data = Z;
		19'b1000101000101100110: color_data = Z;
		19'b1000101000101100111: color_data = Z;
		19'b1000101000101101000: color_data = Z;
		19'b1000101000101101001: color_data = Z;
		19'b1000101000101101010: color_data = Z;
		19'b1000101000101101011: color_data = Z;
		19'b1000101000101101100: color_data = Z;
		19'b1000101000101101101: color_data = Z;
		19'b1000101000101101110: color_data = Z;
		19'b1000101000101101111: color_data = Z;
		19'b1000101000101110000: color_data = Z;
		19'b1000101000101110001: color_data = Z;
		19'b1000101000101110010: color_data = Z;
		19'b1000101000101110011: color_data = Z;
		19'b1000101000101110100: color_data = Z;
		19'b1000101000101110101: color_data = Z;
		19'b1000101000101110110: color_data = Z;
		19'b1000101000101110111: color_data = Z;
		19'b1000101000101111000: color_data = Z;
		19'b1000101000101111001: color_data = Z;
		19'b1000101000101111010: color_data = Z;
		19'b1000101000101111011: color_data = Z;
		19'b1000101000101111100: color_data = Z;
		19'b1000101000101111101: color_data = Z;
		19'b1000101000101111110: color_data = Z;
		19'b1000101000101111111: color_data = Z;
		19'b1000101000110000000: color_data = Z;
		19'b1000101000110000001: color_data = Z;
		19'b1000101000110000010: color_data = Z;
		19'b1000101000110000011: color_data = Z;
		19'b1000101000110000100: color_data = Z;
		19'b1000101000110000101: color_data = Z;
		19'b1000101000110000110: color_data = Z;
		19'b1000101000110000111: color_data = Z;
		19'b1000101000110001000: color_data = Z;
		19'b1000101000110001001: color_data = Z;
		19'b1000101000110001010: color_data = Z;
		19'b1000101000110001011: color_data = Z;
		19'b1000101000110001100: color_data = Z;
		19'b1000101000110001101: color_data = Z;
		19'b1000101000110001110: color_data = Z;
		19'b1000101000110001111: color_data = Z;
		19'b1000101000110010000: color_data = Z;
		19'b1000101000110010001: color_data = Z;
		19'b1000101000110010010: color_data = Z;
		19'b1000101000110010011: color_data = Z;
		19'b1000101000110010100: color_data = Z;
		19'b1000101000110010101: color_data = Z;
		19'b1000101000110010110: color_data = Z;
		19'b1000101000110010111: color_data = Z;
		19'b1000101000110011000: color_data = Z;
		19'b1000101000110011001: color_data = Z;
		19'b1000101000110011010: color_data = Z;
		19'b1000101000110011011: color_data = Z;
		19'b1000101000110011100: color_data = Z;
		19'b1000101000110011101: color_data = Z;
		19'b1000101000110011110: color_data = Z;
		19'b1000101000110011111: color_data = Z;
		19'b1000101000110100000: color_data = Z;
		19'b1000101000110100001: color_data = Z;
		19'b1000101000110100010: color_data = Z;
		19'b1000101000110100011: color_data = Z;
		19'b1000101000110100100: color_data = Z;
		19'b1000101000110100101: color_data = Z;
		19'b1000101000110100110: color_data = Z;
		19'b1000101000110100111: color_data = Z;
		19'b1000101000110101000: color_data = Z;
		19'b1000101000110101001: color_data = Z;
		19'b1000101000110101010: color_data = Z;
		19'b1000101000110101011: color_data = Z;
		19'b1000101000110101100: color_data = Z;
		19'b1000101000110101101: color_data = Z;
		19'b1000101000110101110: color_data = Z;
		19'b1000101000110101111: color_data = Z;
		19'b1000101000110110000: color_data = Z;
		19'b1000101000110110001: color_data = Z;
		19'b1000101000110110010: color_data = Z;
		19'b1000101000110110011: color_data = Z;
		19'b1000101000110110100: color_data = Z;
		19'b1000101000110110101: color_data = Z;
		19'b1000101000110110110: color_data = Z;
		19'b1000101000110110111: color_data = Z;
		19'b1000101000110111000: color_data = Z;
		19'b1000101000110111001: color_data = Z;
		19'b1000101000110111010: color_data = Z;
		19'b1000101000110111011: color_data = Z;
		19'b1000101000110111100: color_data = Z;
		19'b1000101000110111101: color_data = Z;
		19'b1000101000111000111: color_data = Z;
		19'b1000101000111001000: color_data = Z;
		19'b1000101000111001001: color_data = Z;
		19'b1000101000111001010: color_data = Z;
		19'b1000101000111001011: color_data = Z;
		19'b1000101000111001100: color_data = Z;
		19'b1000101000111001101: color_data = Z;
		19'b1000101010011000011: color_data = Z;
		19'b1000101010011000100: color_data = Z;
		19'b1000101010011000101: color_data = Z;
		19'b1000101010011000110: color_data = Z;
		19'b1000101010011000111: color_data = Z;
		19'b1000101010011001000: color_data = Z;
		19'b1000101010011001001: color_data = Z;
		19'b1000101010011001010: color_data = Z;
		19'b1000101010011001011: color_data = Z;
		19'b1000101010011001100: color_data = Z;
		19'b1000101010011001101: color_data = Z;
		19'b1000101010011001110: color_data = Z;
		19'b1000101010011001111: color_data = Z;
		19'b1000101010011010000: color_data = Z;
		19'b1000101010011010001: color_data = Z;
		19'b1000101010011010010: color_data = Z;
		19'b1000101010011010011: color_data = Z;
		19'b1000101010011010100: color_data = Z;
		19'b1000101010011010101: color_data = Z;
		19'b1000101010011010110: color_data = Z;
		19'b1000101010011010111: color_data = Z;
		19'b1000101010011011000: color_data = Z;
		19'b1000101010011011001: color_data = Z;
		19'b1000101010011011010: color_data = Z;
		19'b1000101010011011011: color_data = Z;
		19'b1000101010011011100: color_data = Z;
		19'b1000101010011011101: color_data = Z;
		19'b1000101010011011110: color_data = Z;
		19'b1000101010011011111: color_data = Z;
		19'b1000101010011100000: color_data = Z;
		19'b1000101010011100001: color_data = Z;
		19'b1000101010011100010: color_data = Z;
		19'b1000101010011100011: color_data = Z;
		19'b1000101010011100100: color_data = Z;
		19'b1000101010011100101: color_data = Z;
		19'b1000101010011100110: color_data = Z;
		19'b1000101010011100111: color_data = Z;
		19'b1000101010011101000: color_data = Z;
		19'b1000101010011101001: color_data = Z;
		19'b1000101010011101010: color_data = Z;
		19'b1000101010011101011: color_data = Z;
		19'b1000101010011101100: color_data = Z;
		19'b1000101010011101101: color_data = Z;
		19'b1000101010011101110: color_data = Z;
		19'b1000101010011101111: color_data = Z;
		19'b1000101010011110000: color_data = Z;
		19'b1000101010011110001: color_data = Z;
		19'b1000101010011110010: color_data = Z;
		19'b1000101010011110011: color_data = Z;
		19'b1000101010011110100: color_data = Z;
		19'b1000101010011110101: color_data = Z;
		19'b1000101010011110110: color_data = Z;
		19'b1000101010011110111: color_data = Z;
		19'b1000101010011111000: color_data = Z;
		19'b1000101010011111001: color_data = Z;
		19'b1000101010011111010: color_data = Z;
		19'b1000101010011111011: color_data = Z;
		19'b1000101010011111100: color_data = Z;
		19'b1000101010011111101: color_data = Z;
		19'b1000101010011111110: color_data = Z;
		19'b1000101010011111111: color_data = Z;
		19'b1000101010100000000: color_data = Z;
		19'b1000101010100000001: color_data = Z;
		19'b1000101010100000010: color_data = Z;
		19'b1000101010100000011: color_data = Z;
		19'b1000101010100000100: color_data = Z;
		19'b1000101010100000101: color_data = Z;
		19'b1000101010100000110: color_data = Z;
		19'b1000101010100000111: color_data = Z;
		19'b1000101010100001000: color_data = Z;
		19'b1000101010100001001: color_data = Z;
		19'b1000101010100001010: color_data = Z;
		19'b1000101010100001011: color_data = Z;
		19'b1000101010100001100: color_data = Z;
		19'b1000101010100001101: color_data = Z;
		19'b1000101010100001110: color_data = Z;
		19'b1000101010100001111: color_data = Z;
		19'b1000101010100010000: color_data = Z;
		19'b1000101010100010001: color_data = Z;
		19'b1000101010100010010: color_data = Z;
		19'b1000101010100010011: color_data = Z;
		19'b1000101010100010100: color_data = Z;
		19'b1000101010100010101: color_data = Z;
		19'b1000101010100010111: color_data = Z;
		19'b1000101010100011000: color_data = Z;
		19'b1000101010100101100: color_data = Z;
		19'b1000101010100101101: color_data = Z;
		19'b1000101010100101110: color_data = Z;
		19'b1000101010100101111: color_data = Z;
		19'b1000101010100110000: color_data = Z;
		19'b1000101010100110001: color_data = Z;
		19'b1000101010100110010: color_data = Z;
		19'b1000101010100110011: color_data = Z;
		19'b1000101010100110100: color_data = Z;
		19'b1000101010100110101: color_data = Z;
		19'b1000101010100110110: color_data = Z;
		19'b1000101010100110111: color_data = Z;
		19'b1000101010100111000: color_data = Z;
		19'b1000101010100111001: color_data = Z;
		19'b1000101010100111010: color_data = Z;
		19'b1000101010100111011: color_data = Z;
		19'b1000101010100111100: color_data = Z;
		19'b1000101010100111101: color_data = Z;
		19'b1000101010100111110: color_data = Z;
		19'b1000101010100111111: color_data = Z;
		19'b1000101010101000000: color_data = Z;
		19'b1000101010101000001: color_data = Z;
		19'b1000101010101011011: color_data = Z;
		19'b1000101010101011100: color_data = Z;
		19'b1000101010101011101: color_data = Z;
		19'b1000101010101011110: color_data = Z;
		19'b1000101010101011111: color_data = Z;
		19'b1000101010101100000: color_data = Z;
		19'b1000101010101100001: color_data = Z;
		19'b1000101010101100010: color_data = Z;
		19'b1000101010101100011: color_data = Z;
		19'b1000101010101100100: color_data = Z;
		19'b1000101010101100101: color_data = Z;
		19'b1000101010101100110: color_data = Z;
		19'b1000101010101100111: color_data = Z;
		19'b1000101010101101000: color_data = Z;
		19'b1000101010101101001: color_data = Z;
		19'b1000101010101101010: color_data = Z;
		19'b1000101010101101011: color_data = Z;
		19'b1000101010101101100: color_data = Z;
		19'b1000101010101101101: color_data = Z;
		19'b1000101010101101110: color_data = Z;
		19'b1000101010101101111: color_data = Z;
		19'b1000101010101110000: color_data = Z;
		19'b1000101010101110001: color_data = Z;
		19'b1000101010101110010: color_data = Z;
		19'b1000101010101110011: color_data = Z;
		19'b1000101010101110100: color_data = Z;
		19'b1000101010101110101: color_data = Z;
		19'b1000101010101110110: color_data = Z;
		19'b1000101010101110111: color_data = Z;
		19'b1000101010101111000: color_data = Z;
		19'b1000101010101111001: color_data = Z;
		19'b1000101010101111010: color_data = Z;
		19'b1000101010101111011: color_data = Z;
		19'b1000101010101111100: color_data = Z;
		19'b1000101010101111101: color_data = Z;
		19'b1000101010101111110: color_data = Z;
		19'b1000101010101111111: color_data = Z;
		19'b1000101010110000000: color_data = Z;
		19'b1000101010110000001: color_data = Z;
		19'b1000101010110000010: color_data = Z;
		19'b1000101010110000011: color_data = Z;
		19'b1000101010110000100: color_data = Z;
		19'b1000101010110000101: color_data = Z;
		19'b1000101010110000110: color_data = Z;
		19'b1000101010110000111: color_data = Z;
		19'b1000101010110001000: color_data = Z;
		19'b1000101010110001001: color_data = Z;
		19'b1000101010110001010: color_data = Z;
		19'b1000101010110001011: color_data = Z;
		19'b1000101010110001100: color_data = Z;
		19'b1000101010110001101: color_data = Z;
		19'b1000101010110001110: color_data = Z;
		19'b1000101010110001111: color_data = Z;
		19'b1000101010110010000: color_data = Z;
		19'b1000101010110010001: color_data = Z;
		19'b1000101010110010010: color_data = Z;
		19'b1000101010110010011: color_data = Z;
		19'b1000101010110010100: color_data = Z;
		19'b1000101010110010101: color_data = Z;
		19'b1000101010110010110: color_data = Z;
		19'b1000101010110010111: color_data = Z;
		19'b1000101010110011000: color_data = Z;
		19'b1000101010110011001: color_data = Z;
		19'b1000101010110011010: color_data = Z;
		19'b1000101010110011011: color_data = Z;
		19'b1000101010110011100: color_data = Z;
		19'b1000101010110011101: color_data = Z;
		19'b1000101010110100000: color_data = Z;
		19'b1000101010110100001: color_data = Z;
		19'b1000101010110100010: color_data = Z;
		19'b1000101010110100011: color_data = Z;
		19'b1000101010110100100: color_data = Z;
		19'b1000101010110100101: color_data = Z;
		19'b1000101010110100110: color_data = Z;
		19'b1000101010110100111: color_data = Z;
		19'b1000101010110101000: color_data = Z;
		19'b1000101010110101001: color_data = Z;
		19'b1000101010110101010: color_data = Z;
		19'b1000101010110101011: color_data = Z;
		19'b1000101010110101100: color_data = Z;
		19'b1000101010110101101: color_data = Z;
		19'b1000101010110101110: color_data = Z;
		19'b1000101010110101111: color_data = Z;
		19'b1000101010110110000: color_data = Z;
		19'b1000101010110110001: color_data = Z;
		19'b1000101010110110010: color_data = Z;
		19'b1000101010110110011: color_data = Z;
		19'b1000101010110110100: color_data = Z;
		19'b1000101010110110101: color_data = Z;
		19'b1000101010110110110: color_data = Z;
		19'b1000101010110110111: color_data = Z;
		19'b1000101010110111000: color_data = Z;
		19'b1000101010110111001: color_data = Z;
		19'b1000101010110111010: color_data = Z;
		19'b1000101010110111011: color_data = Z;
		19'b1000101010110111100: color_data = Z;
		19'b1000101010110111101: color_data = Z;
		19'b1000101010111000111: color_data = Z;
		19'b1000101010111001000: color_data = Z;
		19'b1000101010111001001: color_data = Z;
		19'b1000101010111001010: color_data = Z;
		19'b1000101010111001011: color_data = Z;
		19'b1000101010111001100: color_data = Z;
		19'b1000101010111001101: color_data = Z;
		19'b1000101010111001110: color_data = Z;
		19'b1000101100011000100: color_data = Z;
		19'b1000101100011000101: color_data = Z;
		19'b1000101100011000110: color_data = Z;
		19'b1000101100011000111: color_data = Z;
		19'b1000101100011001000: color_data = Z;
		19'b1000101100011001001: color_data = Z;
		19'b1000101100011001010: color_data = Z;
		19'b1000101100011001011: color_data = Z;
		19'b1000101100011001100: color_data = Z;
		19'b1000101100011001101: color_data = Z;
		19'b1000101100011001110: color_data = Z;
		19'b1000101100011001111: color_data = Z;
		19'b1000101100011010000: color_data = Z;
		19'b1000101100011010001: color_data = Z;
		19'b1000101100011010010: color_data = Z;
		19'b1000101100011010011: color_data = Z;
		19'b1000101100011010100: color_data = Z;
		19'b1000101100011010101: color_data = Z;
		19'b1000101100011010110: color_data = Z;
		19'b1000101100011010111: color_data = Z;
		19'b1000101100011011000: color_data = Z;
		19'b1000101100011011001: color_data = Z;
		19'b1000101100011011010: color_data = Z;
		19'b1000101100011011011: color_data = Z;
		19'b1000101100011011100: color_data = Z;
		19'b1000101100011011101: color_data = Z;
		19'b1000101100011011110: color_data = Z;
		19'b1000101100011011111: color_data = Z;
		19'b1000101100011100000: color_data = Z;
		19'b1000101100011100001: color_data = Z;
		19'b1000101100011100010: color_data = Z;
		19'b1000101100011100011: color_data = Z;
		19'b1000101100011100100: color_data = Z;
		19'b1000101100011100101: color_data = Z;
		19'b1000101100011100110: color_data = Z;
		19'b1000101100011100111: color_data = Z;
		19'b1000101100011101000: color_data = Z;
		19'b1000101100011101001: color_data = Z;
		19'b1000101100011101010: color_data = Z;
		19'b1000101100011101011: color_data = Z;
		19'b1000101100011101100: color_data = Z;
		19'b1000101100011101101: color_data = Z;
		19'b1000101100011101110: color_data = Z;
		19'b1000101100011101111: color_data = Z;
		19'b1000101100011110000: color_data = Z;
		19'b1000101100011110001: color_data = Z;
		19'b1000101100011110010: color_data = Z;
		19'b1000101100011110011: color_data = Z;
		19'b1000101100011110100: color_data = Z;
		19'b1000101100011110101: color_data = Z;
		19'b1000101100011110110: color_data = Z;
		19'b1000101100011110111: color_data = Z;
		19'b1000101100011111000: color_data = Z;
		19'b1000101100011111001: color_data = Z;
		19'b1000101100011111010: color_data = Z;
		19'b1000101100011111011: color_data = Z;
		19'b1000101100011111100: color_data = Z;
		19'b1000101100011111101: color_data = Z;
		19'b1000101100011111110: color_data = Z;
		19'b1000101100011111111: color_data = Z;
		19'b1000101100100000000: color_data = Z;
		19'b1000101100100000001: color_data = Z;
		19'b1000101100100000010: color_data = Z;
		19'b1000101100100000011: color_data = Z;
		19'b1000101100100000100: color_data = Z;
		19'b1000101100100000101: color_data = Z;
		19'b1000101100100000110: color_data = Z;
		19'b1000101100100000111: color_data = Z;
		19'b1000101100100001000: color_data = Z;
		19'b1000101100100001001: color_data = Z;
		19'b1000101100100001010: color_data = Z;
		19'b1000101100100001011: color_data = Z;
		19'b1000101100100001100: color_data = Z;
		19'b1000101100100001101: color_data = Z;
		19'b1000101100100001110: color_data = Z;
		19'b1000101100100001111: color_data = Z;
		19'b1000101100100010000: color_data = Z;
		19'b1000101100100010001: color_data = Z;
		19'b1000101100100010010: color_data = Z;
		19'b1000101100100010011: color_data = Z;
		19'b1000101100100010100: color_data = Z;
		19'b1000101100100010101: color_data = Z;
		19'b1000101100100010110: color_data = Z;
		19'b1000101100100010111: color_data = Z;
		19'b1000101100100011000: color_data = Z;
		19'b1000101100100101011: color_data = Z;
		19'b1000101100100101100: color_data = Z;
		19'b1000101100100101101: color_data = Z;
		19'b1000101100100101110: color_data = Z;
		19'b1000101100100101111: color_data = Z;
		19'b1000101100100110000: color_data = Z;
		19'b1000101100100110001: color_data = Z;
		19'b1000101100100110010: color_data = Z;
		19'b1000101100100110011: color_data = Z;
		19'b1000101100100110100: color_data = Z;
		19'b1000101100100110101: color_data = Z;
		19'b1000101100100110110: color_data = Z;
		19'b1000101100100110111: color_data = Z;
		19'b1000101100100111000: color_data = Z;
		19'b1000101100100111001: color_data = Z;
		19'b1000101100100111010: color_data = Z;
		19'b1000101100100111011: color_data = Z;
		19'b1000101100100111100: color_data = Z;
		19'b1000101100100111101: color_data = Z;
		19'b1000101100100111110: color_data = Z;
		19'b1000101100100111111: color_data = Z;
		19'b1000101100101000000: color_data = Z;
		19'b1000101100101000001: color_data = Z;
		19'b1000101100101000010: color_data = Z;
		19'b1000101100101011010: color_data = Z;
		19'b1000101100101011011: color_data = Z;
		19'b1000101100101011100: color_data = Z;
		19'b1000101100101011101: color_data = Z;
		19'b1000101100101011110: color_data = Z;
		19'b1000101100101011111: color_data = Z;
		19'b1000101100101100000: color_data = Z;
		19'b1000101100101100001: color_data = Z;
		19'b1000101100101100010: color_data = Z;
		19'b1000101100101100011: color_data = Z;
		19'b1000101100101100100: color_data = Z;
		19'b1000101100101100101: color_data = Z;
		19'b1000101100101100110: color_data = Z;
		19'b1000101100101100111: color_data = Z;
		19'b1000101100101101000: color_data = Z;
		19'b1000101100101101001: color_data = Z;
		19'b1000101100101101010: color_data = Z;
		19'b1000101100101101011: color_data = Z;
		19'b1000101100101101100: color_data = Z;
		19'b1000101100101101101: color_data = Z;
		19'b1000101100101101110: color_data = Z;
		19'b1000101100101101111: color_data = Z;
		19'b1000101100101110000: color_data = Z;
		19'b1000101100101110001: color_data = Z;
		19'b1000101100101110010: color_data = Z;
		19'b1000101100101110011: color_data = Z;
		19'b1000101100101110100: color_data = Z;
		19'b1000101100101110101: color_data = Z;
		19'b1000101100101110110: color_data = Z;
		19'b1000101100101110111: color_data = Z;
		19'b1000101100101111000: color_data = Z;
		19'b1000101100101111001: color_data = Z;
		19'b1000101100101111010: color_data = Z;
		19'b1000101100101111011: color_data = Z;
		19'b1000101100101111100: color_data = Z;
		19'b1000101100101111101: color_data = Z;
		19'b1000101100101111110: color_data = Z;
		19'b1000101100101111111: color_data = Z;
		19'b1000101100110000000: color_data = Z;
		19'b1000101100110000001: color_data = Z;
		19'b1000101100110000010: color_data = Z;
		19'b1000101100110000011: color_data = Z;
		19'b1000101100110000100: color_data = Z;
		19'b1000101100110000101: color_data = Z;
		19'b1000101100110000110: color_data = Z;
		19'b1000101100110000111: color_data = Z;
		19'b1000101100110001000: color_data = Z;
		19'b1000101100110001001: color_data = Z;
		19'b1000101100110001010: color_data = Z;
		19'b1000101100110001011: color_data = Z;
		19'b1000101100110001100: color_data = Z;
		19'b1000101100110001101: color_data = Z;
		19'b1000101100110001110: color_data = Z;
		19'b1000101100110001111: color_data = Z;
		19'b1000101100110010000: color_data = Z;
		19'b1000101100110010001: color_data = Z;
		19'b1000101100110010010: color_data = Z;
		19'b1000101100110010011: color_data = Z;
		19'b1000101100110010100: color_data = Z;
		19'b1000101100110010101: color_data = Z;
		19'b1000101100110010110: color_data = Z;
		19'b1000101100110010111: color_data = Z;
		19'b1000101100110100100: color_data = Z;
		19'b1000101100110100101: color_data = Z;
		19'b1000101100110100110: color_data = Z;
		19'b1000101100110100111: color_data = Z;
		19'b1000101100110101000: color_data = Z;
		19'b1000101100110101001: color_data = Z;
		19'b1000101100110101010: color_data = Z;
		19'b1000101100110101011: color_data = Z;
		19'b1000101100110101100: color_data = Z;
		19'b1000101100110101101: color_data = Z;
		19'b1000101100110101110: color_data = Z;
		19'b1000101100110101111: color_data = Z;
		19'b1000101100110110000: color_data = Z;
		19'b1000101100110110001: color_data = Z;
		19'b1000101100110110010: color_data = Z;
		19'b1000101100110110011: color_data = Z;
		19'b1000101100110110100: color_data = Z;
		19'b1000101100110110101: color_data = Z;
		19'b1000101100110110110: color_data = Z;
		19'b1000101100110110111: color_data = Z;
		19'b1000101100110111000: color_data = Z;
		19'b1000101100110111001: color_data = Z;
		19'b1000101100110111010: color_data = Z;
		19'b1000101100110111011: color_data = Z;
		19'b1000101100110111100: color_data = Z;
		19'b1000101100110111101: color_data = Z;
		19'b1000101100111000111: color_data = Z;
		19'b1000101100111001000: color_data = Z;
		19'b1000101100111001001: color_data = Z;
		19'b1000101100111001010: color_data = Z;
		19'b1000101100111001011: color_data = Z;
		19'b1000101100111001100: color_data = Z;
		19'b1000101100111001101: color_data = Z;
		19'b1000101100111001110: color_data = Z;
		19'b1000101110011000110: color_data = Z;
		19'b1000101110011000111: color_data = Z;
		19'b1000101110011001000: color_data = Z;
		19'b1000101110011001001: color_data = Z;
		19'b1000101110011001010: color_data = Z;
		19'b1000101110011001011: color_data = Z;
		19'b1000101110011001100: color_data = Z;
		19'b1000101110011001101: color_data = Z;
		19'b1000101110011001110: color_data = Z;
		19'b1000101110011001111: color_data = Z;
		19'b1000101110011010000: color_data = Z;
		19'b1000101110011010001: color_data = Z;
		19'b1000101110011010010: color_data = Z;
		19'b1000101110011010011: color_data = Z;
		19'b1000101110011010100: color_data = Z;
		19'b1000101110011010101: color_data = Z;
		19'b1000101110011010110: color_data = Z;
		19'b1000101110011010111: color_data = Z;
		19'b1000101110011011000: color_data = Z;
		19'b1000101110011011001: color_data = Z;
		19'b1000101110011011010: color_data = Z;
		19'b1000101110011011011: color_data = Z;
		19'b1000101110011011100: color_data = Z;
		19'b1000101110011011101: color_data = Z;
		19'b1000101110011011110: color_data = Z;
		19'b1000101110011011111: color_data = Z;
		19'b1000101110011100000: color_data = Z;
		19'b1000101110011100001: color_data = Z;
		19'b1000101110011100010: color_data = Z;
		19'b1000101110011100011: color_data = Z;
		19'b1000101110011100100: color_data = Z;
		19'b1000101110011100101: color_data = Z;
		19'b1000101110011100110: color_data = Z;
		19'b1000101110011100111: color_data = Z;
		19'b1000101110011101000: color_data = Z;
		19'b1000101110011101001: color_data = Z;
		19'b1000101110011101010: color_data = Z;
		19'b1000101110011101011: color_data = Z;
		19'b1000101110011101100: color_data = Z;
		19'b1000101110011101101: color_data = Z;
		19'b1000101110011101110: color_data = Z;
		19'b1000101110011101111: color_data = Z;
		19'b1000101110011110000: color_data = Z;
		19'b1000101110011110001: color_data = Z;
		19'b1000101110011110010: color_data = Z;
		19'b1000101110011110011: color_data = Z;
		19'b1000101110011110100: color_data = Z;
		19'b1000101110011110101: color_data = Z;
		19'b1000101110011110110: color_data = Z;
		19'b1000101110011110111: color_data = Z;
		19'b1000101110011111000: color_data = Z;
		19'b1000101110011111001: color_data = Z;
		19'b1000101110011111010: color_data = Z;
		19'b1000101110011111011: color_data = Z;
		19'b1000101110011111100: color_data = Z;
		19'b1000101110011111101: color_data = Z;
		19'b1000101110011111110: color_data = Z;
		19'b1000101110011111111: color_data = Z;
		19'b1000101110100000000: color_data = Z;
		19'b1000101110100000001: color_data = Z;
		19'b1000101110100000010: color_data = Z;
		19'b1000101110100000011: color_data = Z;
		19'b1000101110100000100: color_data = Z;
		19'b1000101110100000101: color_data = Z;
		19'b1000101110100000110: color_data = Z;
		19'b1000101110100000111: color_data = Z;
		19'b1000101110100001000: color_data = Z;
		19'b1000101110100001001: color_data = Z;
		19'b1000101110100001010: color_data = Z;
		19'b1000101110100001011: color_data = Z;
		19'b1000101110100001100: color_data = Z;
		19'b1000101110100001101: color_data = Z;
		19'b1000101110100001110: color_data = Z;
		19'b1000101110100001111: color_data = Z;
		19'b1000101110100010000: color_data = Z;
		19'b1000101110100010001: color_data = Z;
		19'b1000101110100010010: color_data = Z;
		19'b1000101110100010011: color_data = Z;
		19'b1000101110100010100: color_data = Z;
		19'b1000101110100010101: color_data = Z;
		19'b1000101110100010110: color_data = Z;
		19'b1000101110100010111: color_data = Z;
		19'b1000101110100101100: color_data = Z;
		19'b1000101110100101101: color_data = Z;
		19'b1000101110100101110: color_data = Z;
		19'b1000101110100101111: color_data = Z;
		19'b1000101110100110000: color_data = Z;
		19'b1000101110100110001: color_data = Z;
		19'b1000101110100110010: color_data = Z;
		19'b1000101110100110011: color_data = Z;
		19'b1000101110100110100: color_data = Z;
		19'b1000101110100110101: color_data = Z;
		19'b1000101110100110110: color_data = Z;
		19'b1000101110100110111: color_data = Z;
		19'b1000101110100111000: color_data = Z;
		19'b1000101110100111001: color_data = Z;
		19'b1000101110100111010: color_data = Z;
		19'b1000101110100111011: color_data = Z;
		19'b1000101110100111100: color_data = Z;
		19'b1000101110100111101: color_data = Z;
		19'b1000101110100111110: color_data = Z;
		19'b1000101110100111111: color_data = Z;
		19'b1000101110101000000: color_data = Z;
		19'b1000101110101000001: color_data = Z;
		19'b1000101110101000010: color_data = Z;
		19'b1000101110101000011: color_data = Z;
		19'b1000101110101011000: color_data = Z;
		19'b1000101110101011001: color_data = Z;
		19'b1000101110101011010: color_data = Z;
		19'b1000101110101011011: color_data = Z;
		19'b1000101110101011100: color_data = Z;
		19'b1000101110101011101: color_data = Z;
		19'b1000101110101011110: color_data = Z;
		19'b1000101110101011111: color_data = Z;
		19'b1000101110101100000: color_data = Z;
		19'b1000101110101100001: color_data = Z;
		19'b1000101110101100010: color_data = Z;
		19'b1000101110101100011: color_data = Z;
		19'b1000101110101100100: color_data = Z;
		19'b1000101110101100101: color_data = Z;
		19'b1000101110101100110: color_data = Z;
		19'b1000101110101100111: color_data = Z;
		19'b1000101110101101000: color_data = Z;
		19'b1000101110101101001: color_data = Z;
		19'b1000101110101101010: color_data = Z;
		19'b1000101110101101011: color_data = Z;
		19'b1000101110101101100: color_data = Z;
		19'b1000101110101101101: color_data = Z;
		19'b1000101110101101110: color_data = Z;
		19'b1000101110101101111: color_data = Z;
		19'b1000101110101110000: color_data = Z;
		19'b1000101110101110001: color_data = Z;
		19'b1000101110101110010: color_data = Z;
		19'b1000101110101110011: color_data = Z;
		19'b1000101110101110100: color_data = Z;
		19'b1000101110101110101: color_data = Z;
		19'b1000101110101110110: color_data = Z;
		19'b1000101110101110111: color_data = Z;
		19'b1000101110101111000: color_data = Z;
		19'b1000101110101111001: color_data = Z;
		19'b1000101110101111010: color_data = Z;
		19'b1000101110101111011: color_data = Z;
		19'b1000101110101111100: color_data = Z;
		19'b1000101110101111101: color_data = Z;
		19'b1000101110101111110: color_data = Z;
		19'b1000101110101111111: color_data = Z;
		19'b1000101110110000000: color_data = Z;
		19'b1000101110110000001: color_data = Z;
		19'b1000101110110000010: color_data = Z;
		19'b1000101110110000011: color_data = Z;
		19'b1000101110110000100: color_data = Z;
		19'b1000101110110000101: color_data = Z;
		19'b1000101110110000110: color_data = Z;
		19'b1000101110110000111: color_data = Z;
		19'b1000101110110001000: color_data = Z;
		19'b1000101110110001001: color_data = Z;
		19'b1000101110110001010: color_data = Z;
		19'b1000101110110001011: color_data = Z;
		19'b1000101110110001100: color_data = Z;
		19'b1000101110110001101: color_data = Z;
		19'b1000101110110001110: color_data = Z;
		19'b1000101110110001111: color_data = Z;
		19'b1000101110110010000: color_data = Z;
		19'b1000101110110010001: color_data = Z;
		19'b1000101110110010010: color_data = Z;
		19'b1000101110110010011: color_data = Z;
		19'b1000101110110010100: color_data = Z;
		19'b1000101110110100101: color_data = Z;
		19'b1000101110110100110: color_data = Z;
		19'b1000101110110100111: color_data = Z;
		19'b1000101110110101000: color_data = Z;
		19'b1000101110110101001: color_data = Z;
		19'b1000101110110101010: color_data = Z;
		19'b1000101110110101011: color_data = Z;
		19'b1000101110110101100: color_data = Z;
		19'b1000101110110101101: color_data = Z;
		19'b1000101110110101110: color_data = Z;
		19'b1000101110110101111: color_data = Z;
		19'b1000101110110110000: color_data = Z;
		19'b1000101110110110001: color_data = Z;
		19'b1000101110110110010: color_data = Z;
		19'b1000101110110110011: color_data = Z;
		19'b1000101110110110100: color_data = Z;
		19'b1000101110110110101: color_data = Z;
		19'b1000101110110110110: color_data = Z;
		19'b1000101110110110111: color_data = Z;
		19'b1000101110110111000: color_data = Z;
		19'b1000101110110111001: color_data = Z;
		19'b1000101110110111010: color_data = Z;
		19'b1000101110110111011: color_data = Z;
		19'b1000101110110111100: color_data = Z;
		19'b1000101110110111101: color_data = Z;
		19'b1000101110111000111: color_data = Z;
		19'b1000101110111001000: color_data = Z;
		19'b1000101110111001001: color_data = Z;
		19'b1000101110111001010: color_data = Z;
		19'b1000101110111001011: color_data = Z;
		19'b1000101110111001100: color_data = Z;
		19'b1000101110111001101: color_data = Z;
		19'b1000101110111001110: color_data = Z;
		19'b1000110000011000111: color_data = Z;
		19'b1000110000011001000: color_data = Z;
		19'b1000110000011001001: color_data = Z;
		19'b1000110000011001010: color_data = Z;
		19'b1000110000011001011: color_data = Z;
		19'b1000110000011001100: color_data = Z;
		19'b1000110000011001101: color_data = Z;
		19'b1000110000011001110: color_data = Z;
		19'b1000110000011001111: color_data = Z;
		19'b1000110000011010000: color_data = Z;
		19'b1000110000011010001: color_data = Z;
		19'b1000110000011010010: color_data = Z;
		19'b1000110000011010011: color_data = Z;
		19'b1000110000011010100: color_data = Z;
		19'b1000110000011010101: color_data = Z;
		19'b1000110000011010110: color_data = Z;
		19'b1000110000011010111: color_data = Z;
		19'b1000110000011011000: color_data = Z;
		19'b1000110000011011001: color_data = Z;
		19'b1000110000011011010: color_data = Z;
		19'b1000110000011011011: color_data = Z;
		19'b1000110000011011100: color_data = Z;
		19'b1000110000011011101: color_data = Z;
		19'b1000110000011011110: color_data = Z;
		19'b1000110000011011111: color_data = Z;
		19'b1000110000011100000: color_data = Z;
		19'b1000110000011100001: color_data = Z;
		19'b1000110000011100010: color_data = Z;
		19'b1000110000011100011: color_data = Z;
		19'b1000110000011100100: color_data = Z;
		19'b1000110000011100101: color_data = Z;
		19'b1000110000011100110: color_data = Z;
		19'b1000110000011100111: color_data = Z;
		19'b1000110000011101000: color_data = Z;
		19'b1000110000011101001: color_data = Z;
		19'b1000110000011101010: color_data = Z;
		19'b1000110000011101011: color_data = Z;
		19'b1000110000011101100: color_data = Z;
		19'b1000110000011101101: color_data = Z;
		19'b1000110000011101110: color_data = Z;
		19'b1000110000011101111: color_data = Z;
		19'b1000110000011110000: color_data = Z;
		19'b1000110000011110001: color_data = Z;
		19'b1000110000011110010: color_data = Z;
		19'b1000110000011110011: color_data = Z;
		19'b1000110000011110100: color_data = Z;
		19'b1000110000011110101: color_data = Z;
		19'b1000110000011110110: color_data = Z;
		19'b1000110000011110111: color_data = Z;
		19'b1000110000011111000: color_data = Z;
		19'b1000110000011111001: color_data = Z;
		19'b1000110000011111010: color_data = Z;
		19'b1000110000011111011: color_data = Z;
		19'b1000110000011111100: color_data = Z;
		19'b1000110000011111101: color_data = Z;
		19'b1000110000011111110: color_data = Z;
		19'b1000110000011111111: color_data = Z;
		19'b1000110000100000000: color_data = Z;
		19'b1000110000100000001: color_data = Z;
		19'b1000110000100000010: color_data = Z;
		19'b1000110000100000011: color_data = Z;
		19'b1000110000100000100: color_data = Z;
		19'b1000110000100000101: color_data = Z;
		19'b1000110000100000110: color_data = Z;
		19'b1000110000100000111: color_data = Z;
		19'b1000110000100001000: color_data = Z;
		19'b1000110000100001001: color_data = Z;
		19'b1000110000100001010: color_data = Z;
		19'b1000110000100001011: color_data = Z;
		19'b1000110000100001100: color_data = Z;
		19'b1000110000100001101: color_data = Z;
		19'b1000110000100001110: color_data = Z;
		19'b1000110000100001111: color_data = Z;
		19'b1000110000100010000: color_data = Z;
		19'b1000110000100010001: color_data = Z;
		19'b1000110000100010010: color_data = Z;
		19'b1000110000100010011: color_data = Z;
		19'b1000110000100010100: color_data = Z;
		19'b1000110000100010101: color_data = Z;
		19'b1000110000100010110: color_data = Z;
		19'b1000110000100010111: color_data = Z;
		19'b1000110000100011000: color_data = Z;
		19'b1000110000100011001: color_data = Z;
		19'b1000110000100101110: color_data = Z;
		19'b1000110000100101111: color_data = Z;
		19'b1000110000100110000: color_data = Z;
		19'b1000110000100110001: color_data = Z;
		19'b1000110000100110010: color_data = Z;
		19'b1000110000100110011: color_data = Z;
		19'b1000110000100110100: color_data = Z;
		19'b1000110000100110101: color_data = Z;
		19'b1000110000100110110: color_data = Z;
		19'b1000110000100110111: color_data = Z;
		19'b1000110000100111000: color_data = Z;
		19'b1000110000100111001: color_data = Z;
		19'b1000110000100111010: color_data = Z;
		19'b1000110000100111011: color_data = Z;
		19'b1000110000100111100: color_data = Z;
		19'b1000110000100111101: color_data = Z;
		19'b1000110000100111110: color_data = Z;
		19'b1000110000100111111: color_data = Z;
		19'b1000110000101000000: color_data = Z;
		19'b1000110000101000001: color_data = Z;
		19'b1000110000101000010: color_data = Z;
		19'b1000110000101000011: color_data = Z;
		19'b1000110000101000100: color_data = Z;
		19'b1000110000101011000: color_data = Z;
		19'b1000110000101011001: color_data = Z;
		19'b1000110000101011010: color_data = Z;
		19'b1000110000101011011: color_data = Z;
		19'b1000110000101011100: color_data = Z;
		19'b1000110000101011101: color_data = Z;
		19'b1000110000101011110: color_data = Z;
		19'b1000110000101011111: color_data = Z;
		19'b1000110000101100000: color_data = Z;
		19'b1000110000101100001: color_data = Z;
		19'b1000110000101100010: color_data = Z;
		19'b1000110000101100011: color_data = Z;
		19'b1000110000101100100: color_data = Z;
		19'b1000110000101100101: color_data = Z;
		19'b1000110000101100110: color_data = Z;
		19'b1000110000101100111: color_data = Z;
		19'b1000110000101101000: color_data = Z;
		19'b1000110000101101001: color_data = Z;
		19'b1000110000101101010: color_data = Z;
		19'b1000110000101101011: color_data = Z;
		19'b1000110000101101100: color_data = Z;
		19'b1000110000101101101: color_data = Z;
		19'b1000110000101101110: color_data = Z;
		19'b1000110000101101111: color_data = Z;
		19'b1000110000101110000: color_data = Z;
		19'b1000110000101110001: color_data = Z;
		19'b1000110000101110010: color_data = Z;
		19'b1000110000101110011: color_data = Z;
		19'b1000110000101110100: color_data = Z;
		19'b1000110000101110101: color_data = Z;
		19'b1000110000101110110: color_data = Z;
		19'b1000110000101110111: color_data = Z;
		19'b1000110000101111000: color_data = Z;
		19'b1000110000101111001: color_data = Z;
		19'b1000110000101111010: color_data = Z;
		19'b1000110000101111011: color_data = Z;
		19'b1000110000101111100: color_data = Z;
		19'b1000110000101111101: color_data = Z;
		19'b1000110000101111110: color_data = Z;
		19'b1000110000101111111: color_data = Z;
		19'b1000110000110000000: color_data = Z;
		19'b1000110000110000001: color_data = Z;
		19'b1000110000110000010: color_data = Z;
		19'b1000110000110000011: color_data = Z;
		19'b1000110000110000100: color_data = Z;
		19'b1000110000110000101: color_data = Z;
		19'b1000110000110000110: color_data = Z;
		19'b1000110000110000111: color_data = Z;
		19'b1000110000110001000: color_data = Z;
		19'b1000110000110001001: color_data = Z;
		19'b1000110000110001010: color_data = Z;
		19'b1000110000110001011: color_data = Z;
		19'b1000110000110001100: color_data = Z;
		19'b1000110000110001101: color_data = Z;
		19'b1000110000110001110: color_data = Z;
		19'b1000110000110001111: color_data = Z;
		19'b1000110000110010000: color_data = Z;
		19'b1000110000110010001: color_data = Z;
		19'b1000110000110010010: color_data = Z;
		19'b1000110000110100110: color_data = Z;
		19'b1000110000110100111: color_data = Z;
		19'b1000110000110101000: color_data = Z;
		19'b1000110000110101001: color_data = Z;
		19'b1000110000110101010: color_data = Z;
		19'b1000110000110101011: color_data = Z;
		19'b1000110000110101100: color_data = Z;
		19'b1000110000110101101: color_data = Z;
		19'b1000110000110101110: color_data = Z;
		19'b1000110000110101111: color_data = Z;
		19'b1000110000110110000: color_data = Z;
		19'b1000110000110110001: color_data = Z;
		19'b1000110000110110010: color_data = Z;
		19'b1000110000110110011: color_data = Z;
		19'b1000110000110110100: color_data = Z;
		19'b1000110000110110101: color_data = Z;
		19'b1000110000110110110: color_data = Z;
		19'b1000110000110110111: color_data = Z;
		19'b1000110000110111000: color_data = Z;
		19'b1000110000110111001: color_data = Z;
		19'b1000110000110111010: color_data = Z;
		19'b1000110000110111011: color_data = Z;
		19'b1000110000110111100: color_data = Z;
		19'b1000110000110111101: color_data = Z;
		19'b1000110000111000111: color_data = Z;
		19'b1000110000111001000: color_data = Z;
		19'b1000110000111001001: color_data = Z;
		19'b1000110000111001010: color_data = Z;
		19'b1000110000111001011: color_data = Z;
		19'b1000110000111001100: color_data = Z;
		19'b1000110000111001101: color_data = Z;
		19'b1000110000111001110: color_data = Z;
		19'b1000110010011001010: color_data = Z;
		19'b1000110010011001011: color_data = Z;
		19'b1000110010011001100: color_data = Z;
		19'b1000110010011001101: color_data = Z;
		19'b1000110010011001110: color_data = Z;
		19'b1000110010011001111: color_data = Z;
		19'b1000110010011010000: color_data = Z;
		19'b1000110010011010001: color_data = Z;
		19'b1000110010011010010: color_data = Z;
		19'b1000110010011010011: color_data = Z;
		19'b1000110010011010100: color_data = Z;
		19'b1000110010011010101: color_data = Z;
		19'b1000110010011010110: color_data = Z;
		19'b1000110010011010111: color_data = Z;
		19'b1000110010011011000: color_data = Z;
		19'b1000110010011011001: color_data = Z;
		19'b1000110010011011010: color_data = Z;
		19'b1000110010011011011: color_data = Z;
		19'b1000110010011011100: color_data = Z;
		19'b1000110010011011101: color_data = Z;
		19'b1000110010011011110: color_data = Z;
		19'b1000110010011011111: color_data = Z;
		19'b1000110010011100000: color_data = Z;
		19'b1000110010011100001: color_data = Z;
		19'b1000110010011100010: color_data = Z;
		19'b1000110010011100011: color_data = Z;
		19'b1000110010011100100: color_data = Z;
		19'b1000110010011100101: color_data = Z;
		19'b1000110010011100110: color_data = Z;
		19'b1000110010011100111: color_data = Z;
		19'b1000110010011101000: color_data = Z;
		19'b1000110010011101001: color_data = Z;
		19'b1000110010011101010: color_data = Z;
		19'b1000110010011101011: color_data = Z;
		19'b1000110010011101100: color_data = Z;
		19'b1000110010011101101: color_data = Z;
		19'b1000110010011101110: color_data = Z;
		19'b1000110010011101111: color_data = Z;
		19'b1000110010011110000: color_data = Z;
		19'b1000110010011110001: color_data = Z;
		19'b1000110010011110010: color_data = Z;
		19'b1000110010011110011: color_data = Z;
		19'b1000110010011110100: color_data = Z;
		19'b1000110010011110101: color_data = Z;
		19'b1000110010011110110: color_data = Z;
		19'b1000110010011110111: color_data = Z;
		19'b1000110010011111000: color_data = Z;
		19'b1000110010011111001: color_data = Z;
		19'b1000110010011111010: color_data = Z;
		19'b1000110010011111011: color_data = Z;
		19'b1000110010011111100: color_data = Z;
		19'b1000110010011111101: color_data = Z;
		19'b1000110010011111110: color_data = Z;
		19'b1000110010011111111: color_data = Z;
		19'b1000110010100000000: color_data = Z;
		19'b1000110010100000001: color_data = Z;
		19'b1000110010100000010: color_data = Z;
		19'b1000110010100000011: color_data = Z;
		19'b1000110010100000100: color_data = Z;
		19'b1000110010100000101: color_data = Z;
		19'b1000110010100000110: color_data = Z;
		19'b1000110010100000111: color_data = Z;
		19'b1000110010100001000: color_data = Z;
		19'b1000110010100001001: color_data = Z;
		19'b1000110010100001010: color_data = Z;
		19'b1000110010100001011: color_data = Z;
		19'b1000110010100001100: color_data = Z;
		19'b1000110010100001101: color_data = Z;
		19'b1000110010100001110: color_data = Z;
		19'b1000110010100001111: color_data = Z;
		19'b1000110010100010000: color_data = Z;
		19'b1000110010100010001: color_data = Z;
		19'b1000110010100010010: color_data = Z;
		19'b1000110010100010011: color_data = Z;
		19'b1000110010100010100: color_data = Z;
		19'b1000110010100010101: color_data = Z;
		19'b1000110010100010110: color_data = Z;
		19'b1000110010100010111: color_data = Z;
		19'b1000110010100011000: color_data = Z;
		19'b1000110010100011001: color_data = Z;
		19'b1000110010100011010: color_data = Z;
		19'b1000110010100011011: color_data = Z;
		19'b1000110010100011100: color_data = Z;
		19'b1000110010100011101: color_data = Z;
		19'b1000110010100101111: color_data = Z;
		19'b1000110010100110000: color_data = Z;
		19'b1000110010100110001: color_data = Z;
		19'b1000110010100110010: color_data = Z;
		19'b1000110010100110011: color_data = Z;
		19'b1000110010100110100: color_data = Z;
		19'b1000110010100110101: color_data = Z;
		19'b1000110010100110110: color_data = Z;
		19'b1000110010100110111: color_data = Z;
		19'b1000110010100111000: color_data = Z;
		19'b1000110010100111001: color_data = Z;
		19'b1000110010100111010: color_data = Z;
		19'b1000110010100111011: color_data = Z;
		19'b1000110010100111100: color_data = Z;
		19'b1000110010100111101: color_data = Z;
		19'b1000110010100111110: color_data = Z;
		19'b1000110010100111111: color_data = Z;
		19'b1000110010101000000: color_data = Z;
		19'b1000110010101000001: color_data = Z;
		19'b1000110010101000010: color_data = Z;
		19'b1000110010101000011: color_data = Z;
		19'b1000110010101000100: color_data = Z;
		19'b1000110010101000101: color_data = Z;
		19'b1000110010101010110: color_data = Z;
		19'b1000110010101010111: color_data = Z;
		19'b1000110010101011000: color_data = Z;
		19'b1000110010101011001: color_data = Z;
		19'b1000110010101011010: color_data = Z;
		19'b1000110010101011011: color_data = Z;
		19'b1000110010101011100: color_data = Z;
		19'b1000110010101011101: color_data = Z;
		19'b1000110010101011110: color_data = Z;
		19'b1000110010101011111: color_data = Z;
		19'b1000110010101100000: color_data = Z;
		19'b1000110010101100001: color_data = Z;
		19'b1000110010101100010: color_data = Z;
		19'b1000110010101100011: color_data = Z;
		19'b1000110010101100100: color_data = Z;
		19'b1000110010101100101: color_data = Z;
		19'b1000110010101100110: color_data = Z;
		19'b1000110010101100111: color_data = Z;
		19'b1000110010101101000: color_data = Z;
		19'b1000110010101101001: color_data = Z;
		19'b1000110010101101010: color_data = Z;
		19'b1000110010101101011: color_data = Z;
		19'b1000110010101101100: color_data = Z;
		19'b1000110010101101101: color_data = Z;
		19'b1000110010101101110: color_data = Z;
		19'b1000110010101101111: color_data = Z;
		19'b1000110010101110000: color_data = Z;
		19'b1000110010101110001: color_data = Z;
		19'b1000110010101110010: color_data = Z;
		19'b1000110010101110011: color_data = Z;
		19'b1000110010101110100: color_data = Z;
		19'b1000110010101110101: color_data = Z;
		19'b1000110010101110110: color_data = Z;
		19'b1000110010101110111: color_data = Z;
		19'b1000110010101111000: color_data = Z;
		19'b1000110010101111001: color_data = Z;
		19'b1000110010101111010: color_data = Z;
		19'b1000110010101111011: color_data = Z;
		19'b1000110010101111100: color_data = Z;
		19'b1000110010101111101: color_data = Z;
		19'b1000110010101111110: color_data = Z;
		19'b1000110010101111111: color_data = Z;
		19'b1000110010110000000: color_data = Z;
		19'b1000110010110000001: color_data = Z;
		19'b1000110010110000010: color_data = Z;
		19'b1000110010110000011: color_data = Z;
		19'b1000110010110000100: color_data = Z;
		19'b1000110010110000101: color_data = Z;
		19'b1000110010110000110: color_data = Z;
		19'b1000110010110000111: color_data = Z;
		19'b1000110010110001000: color_data = Z;
		19'b1000110010110001001: color_data = Z;
		19'b1000110010110001010: color_data = Z;
		19'b1000110010110001011: color_data = Z;
		19'b1000110010110001100: color_data = Z;
		19'b1000110010110001101: color_data = Z;
		19'b1000110010110001110: color_data = Z;
		19'b1000110010110001111: color_data = Z;
		19'b1000110010110010000: color_data = Z;
		19'b1000110010110100111: color_data = Z;
		19'b1000110010110101000: color_data = Z;
		19'b1000110010110101001: color_data = Z;
		19'b1000110010110101010: color_data = Z;
		19'b1000110010110101011: color_data = Z;
		19'b1000110010110101100: color_data = Z;
		19'b1000110010110101101: color_data = Z;
		19'b1000110010110101110: color_data = Z;
		19'b1000110010110101111: color_data = Z;
		19'b1000110010110110000: color_data = Z;
		19'b1000110010110110001: color_data = Z;
		19'b1000110010110110010: color_data = Z;
		19'b1000110010110110011: color_data = Z;
		19'b1000110010110110100: color_data = Z;
		19'b1000110010110110101: color_data = Z;
		19'b1000110010110110110: color_data = Z;
		19'b1000110010110110111: color_data = Z;
		19'b1000110010110111000: color_data = Z;
		19'b1000110010110111001: color_data = Z;
		19'b1000110010110111010: color_data = Z;
		19'b1000110010110111011: color_data = Z;
		19'b1000110010110111100: color_data = Z;
		19'b1000110010110111101: color_data = Z;
		19'b1000110010111000111: color_data = Z;
		19'b1000110010111001000: color_data = Z;
		19'b1000110010111001001: color_data = Z;
		19'b1000110010111001010: color_data = Z;
		19'b1000110010111001011: color_data = Z;
		19'b1000110010111001100: color_data = Z;
		19'b1000110010111001101: color_data = Z;
		19'b1000110010111001110: color_data = Z;
		19'b1000110100011001100: color_data = Z;
		19'b1000110100011001101: color_data = Z;
		19'b1000110100011001110: color_data = Z;
		19'b1000110100011001111: color_data = Z;
		19'b1000110100011010000: color_data = Z;
		19'b1000110100011010001: color_data = Z;
		19'b1000110100011010010: color_data = Z;
		19'b1000110100011010011: color_data = Z;
		19'b1000110100011010100: color_data = Z;
		19'b1000110100011010101: color_data = Z;
		19'b1000110100011010110: color_data = Z;
		19'b1000110100011010111: color_data = Z;
		19'b1000110100011011000: color_data = Z;
		19'b1000110100011011001: color_data = Z;
		19'b1000110100011011010: color_data = Z;
		19'b1000110100011011011: color_data = Z;
		19'b1000110100011011100: color_data = Z;
		19'b1000110100011011101: color_data = Z;
		19'b1000110100011011110: color_data = Z;
		19'b1000110100011011111: color_data = Z;
		19'b1000110100011100000: color_data = Z;
		19'b1000110100011100001: color_data = Z;
		19'b1000110100011100010: color_data = Z;
		19'b1000110100011100011: color_data = Z;
		19'b1000110100011100100: color_data = Z;
		19'b1000110100011100101: color_data = Z;
		19'b1000110100011100110: color_data = Z;
		19'b1000110100011100111: color_data = Z;
		19'b1000110100011101000: color_data = Z;
		19'b1000110100011101001: color_data = Z;
		19'b1000110100011101010: color_data = Z;
		19'b1000110100011101011: color_data = Z;
		19'b1000110100011101100: color_data = Z;
		19'b1000110100011101101: color_data = Z;
		19'b1000110100011101110: color_data = Z;
		19'b1000110100011101111: color_data = Z;
		19'b1000110100011110000: color_data = Z;
		19'b1000110100011110001: color_data = Z;
		19'b1000110100011110010: color_data = Z;
		19'b1000110100011110011: color_data = Z;
		19'b1000110100011110100: color_data = Z;
		19'b1000110100011110101: color_data = Z;
		19'b1000110100011110110: color_data = Z;
		19'b1000110100011110111: color_data = Z;
		19'b1000110100011111000: color_data = Z;
		19'b1000110100011111001: color_data = Z;
		19'b1000110100011111010: color_data = Z;
		19'b1000110100011111011: color_data = Z;
		19'b1000110100011111100: color_data = Z;
		19'b1000110100011111101: color_data = Z;
		19'b1000110100011111110: color_data = Z;
		19'b1000110100011111111: color_data = Z;
		19'b1000110100100000000: color_data = Z;
		19'b1000110100100000001: color_data = Z;
		19'b1000110100100000010: color_data = Z;
		19'b1000110100100000011: color_data = Z;
		19'b1000110100100000100: color_data = Z;
		19'b1000110100100000101: color_data = Z;
		19'b1000110100100000110: color_data = Z;
		19'b1000110100100000111: color_data = Z;
		19'b1000110100100001000: color_data = Z;
		19'b1000110100100001001: color_data = Z;
		19'b1000110100100001010: color_data = Z;
		19'b1000110100100001011: color_data = Z;
		19'b1000110100100001100: color_data = Z;
		19'b1000110100100001101: color_data = Z;
		19'b1000110100100001110: color_data = Z;
		19'b1000110100100001111: color_data = Z;
		19'b1000110100100010000: color_data = Z;
		19'b1000110100100010001: color_data = Z;
		19'b1000110100100010010: color_data = Z;
		19'b1000110100100010011: color_data = Z;
		19'b1000110100100010100: color_data = Z;
		19'b1000110100100010101: color_data = Z;
		19'b1000110100100010110: color_data = Z;
		19'b1000110100100010111: color_data = Z;
		19'b1000110100100011000: color_data = Z;
		19'b1000110100100011001: color_data = Z;
		19'b1000110100100011010: color_data = Z;
		19'b1000110100100011011: color_data = Z;
		19'b1000110100100011100: color_data = Z;
		19'b1000110100100011101: color_data = Z;
		19'b1000110100100011110: color_data = Z;
		19'b1000110100100011111: color_data = Z;
		19'b1000110100100100000: color_data = Z;
		19'b1000110100100100001: color_data = Z;
		19'b1000110100100100010: color_data = Z;
		19'b1000110100100100011: color_data = Z;
		19'b1000110100100100100: color_data = Z;
		19'b1000110100100100101: color_data = Z;
		19'b1000110100100100110: color_data = Z;
		19'b1000110100100101111: color_data = Z;
		19'b1000110100100110000: color_data = Z;
		19'b1000110100100110001: color_data = Z;
		19'b1000110100100110010: color_data = Z;
		19'b1000110100100110011: color_data = Z;
		19'b1000110100100110100: color_data = Z;
		19'b1000110100100110101: color_data = Z;
		19'b1000110100100110110: color_data = Z;
		19'b1000110100100110111: color_data = Z;
		19'b1000110100100111000: color_data = Z;
		19'b1000110100100111001: color_data = Z;
		19'b1000110100100111010: color_data = Z;
		19'b1000110100100111011: color_data = Z;
		19'b1000110100100111100: color_data = Z;
		19'b1000110100100111101: color_data = Z;
		19'b1000110100100111110: color_data = Z;
		19'b1000110100100111111: color_data = Z;
		19'b1000110100101000000: color_data = Z;
		19'b1000110100101000001: color_data = Z;
		19'b1000110100101000010: color_data = Z;
		19'b1000110100101000011: color_data = Z;
		19'b1000110100101000100: color_data = Z;
		19'b1000110100101000101: color_data = Z;
		19'b1000110100101000110: color_data = Z;
		19'b1000110100101000111: color_data = Z;
		19'b1000110100101010101: color_data = Z;
		19'b1000110100101010110: color_data = Z;
		19'b1000110100101010111: color_data = Z;
		19'b1000110100101011000: color_data = Z;
		19'b1000110100101011001: color_data = Z;
		19'b1000110100101011010: color_data = Z;
		19'b1000110100101011011: color_data = Z;
		19'b1000110100101011100: color_data = Z;
		19'b1000110100101011101: color_data = Z;
		19'b1000110100101011110: color_data = Z;
		19'b1000110100101011111: color_data = Z;
		19'b1000110100101100000: color_data = Z;
		19'b1000110100101100001: color_data = Z;
		19'b1000110100101100010: color_data = Z;
		19'b1000110100101100011: color_data = Z;
		19'b1000110100101100100: color_data = Z;
		19'b1000110100101100101: color_data = Z;
		19'b1000110100101100110: color_data = Z;
		19'b1000110100101100111: color_data = Z;
		19'b1000110100101101000: color_data = Z;
		19'b1000110100101101001: color_data = Z;
		19'b1000110100101101010: color_data = Z;
		19'b1000110100101101011: color_data = Z;
		19'b1000110100101101100: color_data = Z;
		19'b1000110100101101101: color_data = Z;
		19'b1000110100101101110: color_data = Z;
		19'b1000110100101101111: color_data = Z;
		19'b1000110100101110000: color_data = Z;
		19'b1000110100101110001: color_data = Z;
		19'b1000110100101110010: color_data = Z;
		19'b1000110100101110011: color_data = Z;
		19'b1000110100101110100: color_data = Z;
		19'b1000110100101110101: color_data = Z;
		19'b1000110100101110110: color_data = Z;
		19'b1000110100101110111: color_data = Z;
		19'b1000110100101111000: color_data = Z;
		19'b1000110100101111001: color_data = Z;
		19'b1000110100101111010: color_data = Z;
		19'b1000110100101111011: color_data = Z;
		19'b1000110100101111100: color_data = Z;
		19'b1000110100101111101: color_data = Z;
		19'b1000110100101111110: color_data = Z;
		19'b1000110100101111111: color_data = Z;
		19'b1000110100110000000: color_data = Z;
		19'b1000110100110000001: color_data = Z;
		19'b1000110100110000010: color_data = Z;
		19'b1000110100110000011: color_data = Z;
		19'b1000110100110000100: color_data = Z;
		19'b1000110100110000101: color_data = Z;
		19'b1000110100110000110: color_data = Z;
		19'b1000110100110000111: color_data = Z;
		19'b1000110100110001000: color_data = Z;
		19'b1000110100110001001: color_data = Z;
		19'b1000110100110001010: color_data = Z;
		19'b1000110100110001011: color_data = Z;
		19'b1000110100110001100: color_data = Z;
		19'b1000110100110001101: color_data = Z;
		19'b1000110100110001110: color_data = Z;
		19'b1000110100110101000: color_data = Z;
		19'b1000110100110101001: color_data = Z;
		19'b1000110100110101010: color_data = Z;
		19'b1000110100110101011: color_data = Z;
		19'b1000110100110101100: color_data = Z;
		19'b1000110100110101101: color_data = Z;
		19'b1000110100110101110: color_data = Z;
		19'b1000110100110101111: color_data = Z;
		19'b1000110100110110000: color_data = Z;
		19'b1000110100110110001: color_data = Z;
		19'b1000110100110110010: color_data = Z;
		19'b1000110100110110011: color_data = Z;
		19'b1000110100110110100: color_data = Z;
		19'b1000110100110110101: color_data = Z;
		19'b1000110100110110110: color_data = Z;
		19'b1000110100110110111: color_data = Z;
		19'b1000110100110111000: color_data = Z;
		19'b1000110100110111001: color_data = Z;
		19'b1000110100110111010: color_data = Z;
		19'b1000110100110111011: color_data = Z;
		19'b1000110100110111100: color_data = Z;
		19'b1000110100110111101: color_data = Z;
		19'b1000110100111000111: color_data = Z;
		19'b1000110100111001001: color_data = Z;
		19'b1000110100111001010: color_data = Z;
		19'b1000110100111001011: color_data = Z;
		19'b1000110100111001100: color_data = Z;
		19'b1000110100111001101: color_data = Z;
		19'b1000110100111001110: color_data = Z;
		19'b1000110110011001110: color_data = Z;
		19'b1000110110011001111: color_data = Z;
		19'b1000110110011010000: color_data = Z;
		19'b1000110110011010001: color_data = Z;
		19'b1000110110011010010: color_data = Z;
		19'b1000110110011010011: color_data = Z;
		19'b1000110110011010100: color_data = Z;
		19'b1000110110011010101: color_data = Z;
		19'b1000110110011010110: color_data = Z;
		19'b1000110110011010111: color_data = Z;
		19'b1000110110011011000: color_data = Z;
		19'b1000110110011011001: color_data = Z;
		19'b1000110110011011010: color_data = Z;
		19'b1000110110011011011: color_data = Z;
		19'b1000110110011011100: color_data = Z;
		19'b1000110110011011101: color_data = Z;
		19'b1000110110011011110: color_data = Z;
		19'b1000110110011011111: color_data = Z;
		19'b1000110110011100000: color_data = Z;
		19'b1000110110011100001: color_data = Z;
		19'b1000110110011100010: color_data = Z;
		19'b1000110110011100011: color_data = Z;
		19'b1000110110011100100: color_data = Z;
		19'b1000110110011100101: color_data = Z;
		19'b1000110110011100110: color_data = Z;
		19'b1000110110011100111: color_data = Z;
		19'b1000110110011101000: color_data = Z;
		19'b1000110110011101001: color_data = Z;
		19'b1000110110011101010: color_data = Z;
		19'b1000110110011101011: color_data = Z;
		19'b1000110110011101100: color_data = Z;
		19'b1000110110011101101: color_data = Z;
		19'b1000110110011101110: color_data = Z;
		19'b1000110110011101111: color_data = Z;
		19'b1000110110011110000: color_data = Z;
		19'b1000110110011110001: color_data = Z;
		19'b1000110110011110010: color_data = Z;
		19'b1000110110011110011: color_data = Z;
		19'b1000110110011110100: color_data = Z;
		19'b1000110110011110101: color_data = Z;
		19'b1000110110011110110: color_data = Z;
		19'b1000110110011110111: color_data = Z;
		19'b1000110110011111000: color_data = Z;
		19'b1000110110011111001: color_data = Z;
		19'b1000110110011111010: color_data = Z;
		19'b1000110110011111011: color_data = Z;
		19'b1000110110011111100: color_data = Z;
		19'b1000110110011111101: color_data = Z;
		19'b1000110110011111110: color_data = Z;
		19'b1000110110011111111: color_data = Z;
		19'b1000110110100000000: color_data = Z;
		19'b1000110110100000001: color_data = Z;
		19'b1000110110100000010: color_data = Z;
		19'b1000110110100000011: color_data = Z;
		19'b1000110110100000100: color_data = Z;
		19'b1000110110100000101: color_data = Z;
		19'b1000110110100000110: color_data = Z;
		19'b1000110110100000111: color_data = Z;
		19'b1000110110100001000: color_data = Z;
		19'b1000110110100001001: color_data = Z;
		19'b1000110110100001010: color_data = Z;
		19'b1000110110100001011: color_data = Z;
		19'b1000110110100001100: color_data = Z;
		19'b1000110110100001101: color_data = Z;
		19'b1000110110100001110: color_data = Z;
		19'b1000110110100001111: color_data = Z;
		19'b1000110110100010000: color_data = Z;
		19'b1000110110100010001: color_data = Z;
		19'b1000110110100010010: color_data = Z;
		19'b1000110110100010011: color_data = Z;
		19'b1000110110100010100: color_data = Z;
		19'b1000110110100010101: color_data = Z;
		19'b1000110110100010110: color_data = Z;
		19'b1000110110100010111: color_data = Z;
		19'b1000110110100011000: color_data = Z;
		19'b1000110110100011001: color_data = Z;
		19'b1000110110100011010: color_data = Z;
		19'b1000110110100011011: color_data = Z;
		19'b1000110110100011100: color_data = Z;
		19'b1000110110100011101: color_data = Z;
		19'b1000110110100011110: color_data = Z;
		19'b1000110110100011111: color_data = Z;
		19'b1000110110100100000: color_data = Z;
		19'b1000110110100100001: color_data = Z;
		19'b1000110110100100010: color_data = Z;
		19'b1000110110100100011: color_data = Z;
		19'b1000110110100100100: color_data = Z;
		19'b1000110110100100101: color_data = Z;
		19'b1000110110100100110: color_data = Z;
		19'b1000110110100100111: color_data = Z;
		19'b1000110110100101000: color_data = Z;
		19'b1000110110100101001: color_data = Z;
		19'b1000110110100101010: color_data = Z;
		19'b1000110110100101011: color_data = Z;
		19'b1000110110100101100: color_data = Z;
		19'b1000110110100101101: color_data = Z;
		19'b1000110110100101110: color_data = Z;
		19'b1000110110100101111: color_data = Z;
		19'b1000110110100110000: color_data = Z;
		19'b1000110110100110001: color_data = Z;
		19'b1000110110100110010: color_data = Z;
		19'b1000110110100110011: color_data = Z;
		19'b1000110110100110100: color_data = Z;
		19'b1000110110100110101: color_data = Z;
		19'b1000110110100110110: color_data = Z;
		19'b1000110110100110111: color_data = Z;
		19'b1000110110100111000: color_data = Z;
		19'b1000110110100111001: color_data = Z;
		19'b1000110110100111010: color_data = Z;
		19'b1000110110100111011: color_data = Z;
		19'b1000110110100111100: color_data = Z;
		19'b1000110110100111101: color_data = Z;
		19'b1000110110100111110: color_data = Z;
		19'b1000110110100111111: color_data = Z;
		19'b1000110110101000000: color_data = Z;
		19'b1000110110101000001: color_data = Z;
		19'b1000110110101000010: color_data = Z;
		19'b1000110110101000011: color_data = Z;
		19'b1000110110101000100: color_data = Z;
		19'b1000110110101000101: color_data = Z;
		19'b1000110110101000110: color_data = Z;
		19'b1000110110101000111: color_data = Z;
		19'b1000110110101001000: color_data = Z;
		19'b1000110110101010010: color_data = Z;
		19'b1000110110101010011: color_data = Z;
		19'b1000110110101010100: color_data = Z;
		19'b1000110110101010101: color_data = Z;
		19'b1000110110101010110: color_data = Z;
		19'b1000110110101010111: color_data = Z;
		19'b1000110110101011000: color_data = Z;
		19'b1000110110101011001: color_data = Z;
		19'b1000110110101011010: color_data = Z;
		19'b1000110110101011011: color_data = Z;
		19'b1000110110101011100: color_data = Z;
		19'b1000110110101011101: color_data = Z;
		19'b1000110110101011110: color_data = Z;
		19'b1000110110101011111: color_data = Z;
		19'b1000110110101100000: color_data = Z;
		19'b1000110110101100001: color_data = Z;
		19'b1000110110101100010: color_data = Z;
		19'b1000110110101100011: color_data = Z;
		19'b1000110110101100100: color_data = Z;
		19'b1000110110101100101: color_data = Z;
		19'b1000110110101100110: color_data = Z;
		19'b1000110110101100111: color_data = Z;
		19'b1000110110101101000: color_data = Z;
		19'b1000110110101101001: color_data = Z;
		19'b1000110110101101010: color_data = Z;
		19'b1000110110101101011: color_data = Z;
		19'b1000110110101101100: color_data = Z;
		19'b1000110110101101101: color_data = Z;
		19'b1000110110101101110: color_data = Z;
		19'b1000110110101101111: color_data = Z;
		19'b1000110110101110000: color_data = Z;
		19'b1000110110101110001: color_data = Z;
		19'b1000110110101110010: color_data = Z;
		19'b1000110110101110011: color_data = Z;
		19'b1000110110101110100: color_data = Z;
		19'b1000110110101110101: color_data = Z;
		19'b1000110110101110110: color_data = Z;
		19'b1000110110101110111: color_data = Z;
		19'b1000110110101111000: color_data = Z;
		19'b1000110110101111001: color_data = Z;
		19'b1000110110101111010: color_data = Z;
		19'b1000110110101111011: color_data = Z;
		19'b1000110110101111100: color_data = Z;
		19'b1000110110101111101: color_data = Z;
		19'b1000110110101111110: color_data = Z;
		19'b1000110110101111111: color_data = Z;
		19'b1000110110110000000: color_data = Z;
		19'b1000110110110000001: color_data = Z;
		19'b1000110110110000010: color_data = Z;
		19'b1000110110110000011: color_data = Z;
		19'b1000110110110000100: color_data = Z;
		19'b1000110110110000101: color_data = Z;
		19'b1000110110110000110: color_data = Z;
		19'b1000110110110000111: color_data = Z;
		19'b1000110110110001000: color_data = Z;
		19'b1000110110110001001: color_data = Z;
		19'b1000110110110001010: color_data = Z;
		19'b1000110110110001011: color_data = Z;
		19'b1000110110110101001: color_data = Z;
		19'b1000110110110101010: color_data = Z;
		19'b1000110110110101011: color_data = Z;
		19'b1000110110110101100: color_data = Z;
		19'b1000110110110101101: color_data = Z;
		19'b1000110110110101110: color_data = Z;
		19'b1000110110110101111: color_data = Z;
		19'b1000110110110110000: color_data = Z;
		19'b1000110110110110001: color_data = Z;
		19'b1000110110110110010: color_data = Z;
		19'b1000110110110110011: color_data = Z;
		19'b1000110110110110100: color_data = Z;
		19'b1000110110110110101: color_data = Z;
		19'b1000110110110110110: color_data = Z;
		19'b1000110110110110111: color_data = Z;
		19'b1000110110110111000: color_data = Z;
		19'b1000110110110111001: color_data = Z;
		19'b1000110110110111010: color_data = Z;
		19'b1000110110110111011: color_data = Z;
		19'b1000110110110111100: color_data = Z;
		19'b1000110110110111101: color_data = Z;
		19'b1000110110111000111: color_data = Z;
		19'b1000110110111001001: color_data = Z;
		19'b1000110110111001010: color_data = Z;
		19'b1000110110111001011: color_data = Z;
		19'b1000110110111001100: color_data = Z;
		19'b1000110110111001101: color_data = Z;
		19'b1000110110111001110: color_data = Z;
		19'b1000111000011010000: color_data = Z;
		19'b1000111000011010001: color_data = Z;
		19'b1000111000011010010: color_data = Z;
		19'b1000111000011010011: color_data = Z;
		19'b1000111000011010100: color_data = Z;
		19'b1000111000011010101: color_data = Z;
		19'b1000111000011010110: color_data = Z;
		19'b1000111000011010111: color_data = Z;
		19'b1000111000011011000: color_data = Z;
		19'b1000111000011011001: color_data = Z;
		19'b1000111000011011010: color_data = Z;
		19'b1000111000011011011: color_data = Z;
		19'b1000111000011011100: color_data = Z;
		19'b1000111000011011101: color_data = Z;
		19'b1000111000011011110: color_data = Z;
		19'b1000111000011011111: color_data = Z;
		19'b1000111000011100000: color_data = Z;
		19'b1000111000011100001: color_data = Z;
		19'b1000111000011100010: color_data = Z;
		19'b1000111000011100011: color_data = Z;
		19'b1000111000011100100: color_data = Z;
		19'b1000111000011100101: color_data = Z;
		19'b1000111000011100110: color_data = Z;
		19'b1000111000011100111: color_data = Z;
		19'b1000111000011101000: color_data = Z;
		19'b1000111000011101001: color_data = Z;
		19'b1000111000011101010: color_data = Z;
		19'b1000111000011101011: color_data = Z;
		19'b1000111000011101100: color_data = Z;
		19'b1000111000011101101: color_data = Z;
		19'b1000111000011101110: color_data = Z;
		19'b1000111000011101111: color_data = Z;
		19'b1000111000011110000: color_data = Z;
		19'b1000111000011110001: color_data = Z;
		19'b1000111000011110010: color_data = Z;
		19'b1000111000011110011: color_data = Z;
		19'b1000111000011110100: color_data = Z;
		19'b1000111000011110101: color_data = Z;
		19'b1000111000011110110: color_data = Z;
		19'b1000111000011110111: color_data = Z;
		19'b1000111000011111000: color_data = Z;
		19'b1000111000011111001: color_data = Z;
		19'b1000111000011111010: color_data = Z;
		19'b1000111000011111011: color_data = Z;
		19'b1000111000011111100: color_data = Z;
		19'b1000111000011111101: color_data = Z;
		19'b1000111000011111110: color_data = Z;
		19'b1000111000011111111: color_data = Z;
		19'b1000111000100000000: color_data = Z;
		19'b1000111000100000001: color_data = Z;
		19'b1000111000100000010: color_data = Z;
		19'b1000111000100000011: color_data = Z;
		19'b1000111000100000100: color_data = Z;
		19'b1000111000100000101: color_data = Z;
		19'b1000111000100000110: color_data = Z;
		19'b1000111000100000111: color_data = Z;
		19'b1000111000100001000: color_data = Z;
		19'b1000111000100001001: color_data = Z;
		19'b1000111000100001010: color_data = Z;
		19'b1000111000100001011: color_data = Z;
		19'b1000111000100001100: color_data = Z;
		19'b1000111000100001101: color_data = Z;
		19'b1000111000100001110: color_data = Z;
		19'b1000111000100001111: color_data = Z;
		19'b1000111000100010000: color_data = Z;
		19'b1000111000100010001: color_data = Z;
		19'b1000111000100010010: color_data = Z;
		19'b1000111000100010011: color_data = Z;
		19'b1000111000100010100: color_data = Z;
		19'b1000111000100010101: color_data = Z;
		19'b1000111000100010110: color_data = Z;
		19'b1000111000100010111: color_data = Z;
		19'b1000111000100011000: color_data = Z;
		19'b1000111000100011001: color_data = Z;
		19'b1000111000100011010: color_data = Z;
		19'b1000111000100011011: color_data = Z;
		19'b1000111000100011100: color_data = Z;
		19'b1000111000100011101: color_data = Z;
		19'b1000111000100011110: color_data = Z;
		19'b1000111000100011111: color_data = Z;
		19'b1000111000100100000: color_data = Z;
		19'b1000111000100100001: color_data = Z;
		19'b1000111000100100010: color_data = Z;
		19'b1000111000100100011: color_data = Z;
		19'b1000111000100100100: color_data = Z;
		19'b1000111000100100101: color_data = Z;
		19'b1000111000100100110: color_data = Z;
		19'b1000111000100100111: color_data = Z;
		19'b1000111000100101000: color_data = Z;
		19'b1000111000100101001: color_data = Z;
		19'b1000111000100101010: color_data = Z;
		19'b1000111000100101011: color_data = Z;
		19'b1000111000100101100: color_data = Z;
		19'b1000111000100101101: color_data = Z;
		19'b1000111000100101110: color_data = Z;
		19'b1000111000100101111: color_data = Z;
		19'b1000111000100110000: color_data = Z;
		19'b1000111000100110001: color_data = Z;
		19'b1000111000100110010: color_data = Z;
		19'b1000111000100110011: color_data = Z;
		19'b1000111000100110100: color_data = Z;
		19'b1000111000100110101: color_data = Z;
		19'b1000111000100110110: color_data = Z;
		19'b1000111000100110111: color_data = Z;
		19'b1000111000100111000: color_data = Z;
		19'b1000111000100111001: color_data = Z;
		19'b1000111000100111010: color_data = Z;
		19'b1000111000100111011: color_data = Z;
		19'b1000111000100111100: color_data = Z;
		19'b1000111000100111101: color_data = Z;
		19'b1000111000100111110: color_data = Z;
		19'b1000111000100111111: color_data = Z;
		19'b1000111000101000000: color_data = Z;
		19'b1000111000101000001: color_data = Z;
		19'b1000111000101000010: color_data = Z;
		19'b1000111000101000011: color_data = Z;
		19'b1000111000101000100: color_data = Z;
		19'b1000111000101000101: color_data = Z;
		19'b1000111000101000110: color_data = Z;
		19'b1000111000101000111: color_data = Z;
		19'b1000111000101001000: color_data = Z;
		19'b1000111000101001001: color_data = Z;
		19'b1000111000101001010: color_data = Z;
		19'b1000111000101001011: color_data = Z;
		19'b1000111000101001100: color_data = Z;
		19'b1000111000101001101: color_data = Z;
		19'b1000111000101001110: color_data = Z;
		19'b1000111000101001111: color_data = Z;
		19'b1000111000101010000: color_data = Z;
		19'b1000111000101010001: color_data = Z;
		19'b1000111000101010010: color_data = Z;
		19'b1000111000101010011: color_data = Z;
		19'b1000111000101010100: color_data = Z;
		19'b1000111000101010101: color_data = Z;
		19'b1000111000101010110: color_data = Z;
		19'b1000111000101010111: color_data = Z;
		19'b1000111000101011000: color_data = Z;
		19'b1000111000101011001: color_data = Z;
		19'b1000111000101011010: color_data = Z;
		19'b1000111000101011011: color_data = Z;
		19'b1000111000101011100: color_data = Z;
		19'b1000111000101011101: color_data = Z;
		19'b1000111000101011110: color_data = Z;
		19'b1000111000101011111: color_data = Z;
		19'b1000111000101100000: color_data = Z;
		19'b1000111000101100001: color_data = Z;
		19'b1000111000101100010: color_data = Z;
		19'b1000111000101100011: color_data = Z;
		19'b1000111000101100100: color_data = Z;
		19'b1000111000101100101: color_data = Z;
		19'b1000111000101100110: color_data = Z;
		19'b1000111000101100111: color_data = Z;
		19'b1000111000101101000: color_data = Z;
		19'b1000111000101101001: color_data = Z;
		19'b1000111000101101010: color_data = Z;
		19'b1000111000101101011: color_data = Z;
		19'b1000111000101101100: color_data = Z;
		19'b1000111000101101101: color_data = Z;
		19'b1000111000101101110: color_data = Z;
		19'b1000111000101101111: color_data = Z;
		19'b1000111000101110000: color_data = Z;
		19'b1000111000101110001: color_data = Z;
		19'b1000111000101110010: color_data = Z;
		19'b1000111000101110011: color_data = Z;
		19'b1000111000101110100: color_data = Z;
		19'b1000111000101110101: color_data = Z;
		19'b1000111000101110110: color_data = Z;
		19'b1000111000101110111: color_data = Z;
		19'b1000111000101111000: color_data = Z;
		19'b1000111000101111001: color_data = Z;
		19'b1000111000101111010: color_data = Z;
		19'b1000111000101111011: color_data = Z;
		19'b1000111000101111100: color_data = Z;
		19'b1000111000101111101: color_data = Z;
		19'b1000111000101111110: color_data = Z;
		19'b1000111000101111111: color_data = Z;
		19'b1000111000110000000: color_data = Z;
		19'b1000111000110000001: color_data = Z;
		19'b1000111000110000010: color_data = Z;
		19'b1000111000110000011: color_data = Z;
		19'b1000111000110000100: color_data = Z;
		19'b1000111000110000101: color_data = Z;
		19'b1000111000110000110: color_data = Z;
		19'b1000111000110000111: color_data = Z;
		19'b1000111000110001000: color_data = Z;
		19'b1000111000110001001: color_data = Z;
		19'b1000111000110101001: color_data = Z;
		19'b1000111000110101010: color_data = Z;
		19'b1000111000110101011: color_data = Z;
		19'b1000111000110101100: color_data = Z;
		19'b1000111000110101101: color_data = Z;
		19'b1000111000110101110: color_data = Z;
		19'b1000111000110101111: color_data = Z;
		19'b1000111000110110000: color_data = Z;
		19'b1000111000110110001: color_data = Z;
		19'b1000111000110110010: color_data = Z;
		19'b1000111000110110011: color_data = Z;
		19'b1000111000110110100: color_data = Z;
		19'b1000111000110110101: color_data = Z;
		19'b1000111000110110110: color_data = Z;
		19'b1000111000110110111: color_data = Z;
		19'b1000111000110111000: color_data = Z;
		19'b1000111000110111001: color_data = Z;
		19'b1000111000110111010: color_data = Z;
		19'b1000111000110111011: color_data = Z;
		19'b1000111000110111100: color_data = Z;
		19'b1000111000110111101: color_data = Z;
		19'b1000111000111000111: color_data = Z;
		19'b1000111000111001001: color_data = Z;
		19'b1000111000111001010: color_data = Z;
		19'b1000111000111001011: color_data = Z;
		19'b1000111000111001100: color_data = Z;
		19'b1000111000111001101: color_data = Z;
		19'b1000111010011010010: color_data = Z;
		19'b1000111010011010011: color_data = Z;
		19'b1000111010011010100: color_data = Z;
		19'b1000111010011010101: color_data = Z;
		19'b1000111010011010110: color_data = Z;
		19'b1000111010011010111: color_data = Z;
		19'b1000111010011011000: color_data = Z;
		19'b1000111010011011001: color_data = Z;
		19'b1000111010011011010: color_data = Z;
		19'b1000111010011011011: color_data = Z;
		19'b1000111010011011100: color_data = Z;
		19'b1000111010011011101: color_data = Z;
		19'b1000111010011011110: color_data = Z;
		19'b1000111010011011111: color_data = Z;
		19'b1000111010011100000: color_data = Z;
		19'b1000111010011100001: color_data = Z;
		19'b1000111010011100010: color_data = Z;
		19'b1000111010011100011: color_data = Z;
		19'b1000111010011100100: color_data = Z;
		19'b1000111010011100101: color_data = Z;
		19'b1000111010011100110: color_data = Z;
		19'b1000111010011100111: color_data = Z;
		19'b1000111010011101000: color_data = Z;
		19'b1000111010011101001: color_data = Z;
		19'b1000111010011101010: color_data = Z;
		19'b1000111010011101011: color_data = Z;
		19'b1000111010011101100: color_data = Z;
		19'b1000111010011101101: color_data = Z;
		19'b1000111010011101110: color_data = Z;
		19'b1000111010011101111: color_data = Z;
		19'b1000111010011110000: color_data = Z;
		19'b1000111010011110001: color_data = Z;
		19'b1000111010011110010: color_data = Z;
		19'b1000111010011110011: color_data = Z;
		19'b1000111010011110100: color_data = Z;
		19'b1000111010011110101: color_data = Z;
		19'b1000111010011110110: color_data = Z;
		19'b1000111010011110111: color_data = Z;
		19'b1000111010011111000: color_data = Z;
		19'b1000111010011111001: color_data = Z;
		19'b1000111010011111010: color_data = Z;
		19'b1000111010011111011: color_data = Z;
		19'b1000111010011111100: color_data = Z;
		19'b1000111010011111101: color_data = Z;
		19'b1000111010011111110: color_data = Z;
		19'b1000111010011111111: color_data = Z;
		19'b1000111010100000000: color_data = Z;
		19'b1000111010100000001: color_data = Z;
		19'b1000111010100000010: color_data = Z;
		19'b1000111010100000011: color_data = Z;
		19'b1000111010100000100: color_data = Z;
		19'b1000111010100000101: color_data = Z;
		19'b1000111010100000110: color_data = Z;
		19'b1000111010100000111: color_data = Z;
		19'b1000111010100001000: color_data = Z;
		19'b1000111010100001001: color_data = Z;
		19'b1000111010100001010: color_data = Z;
		19'b1000111010100001011: color_data = Z;
		19'b1000111010100001100: color_data = Z;
		19'b1000111010100001101: color_data = Z;
		19'b1000111010100001110: color_data = Z;
		19'b1000111010100001111: color_data = Z;
		19'b1000111010100010000: color_data = Z;
		19'b1000111010100010001: color_data = Z;
		19'b1000111010100010010: color_data = Z;
		19'b1000111010100010011: color_data = Z;
		19'b1000111010100010100: color_data = Z;
		19'b1000111010100010101: color_data = Z;
		19'b1000111010100010110: color_data = Z;
		19'b1000111010100010111: color_data = Z;
		19'b1000111010100011000: color_data = Z;
		19'b1000111010100011001: color_data = Z;
		19'b1000111010100011010: color_data = Z;
		19'b1000111010100011011: color_data = Z;
		19'b1000111010100011100: color_data = Z;
		19'b1000111010100011101: color_data = Z;
		19'b1000111010100011110: color_data = Z;
		19'b1000111010100011111: color_data = Z;
		19'b1000111010100100000: color_data = Z;
		19'b1000111010100100001: color_data = Z;
		19'b1000111010100100010: color_data = Z;
		19'b1000111010100100011: color_data = Z;
		19'b1000111010100100100: color_data = Z;
		19'b1000111010100100101: color_data = Z;
		19'b1000111010100100110: color_data = Z;
		19'b1000111010100100111: color_data = Z;
		19'b1000111010100101000: color_data = Z;
		19'b1000111010100101001: color_data = Z;
		19'b1000111010100101010: color_data = Z;
		19'b1000111010100101011: color_data = Z;
		19'b1000111010100101100: color_data = Z;
		19'b1000111010100101101: color_data = Z;
		19'b1000111010100101110: color_data = Z;
		19'b1000111010100101111: color_data = Z;
		19'b1000111010100110000: color_data = Z;
		19'b1000111010100110001: color_data = Z;
		19'b1000111010100110010: color_data = Z;
		19'b1000111010100110011: color_data = Z;
		19'b1000111010100110100: color_data = Z;
		19'b1000111010100110101: color_data = Z;
		19'b1000111010100110110: color_data = Z;
		19'b1000111010100110111: color_data = Z;
		19'b1000111010100111000: color_data = Z;
		19'b1000111010100111001: color_data = Z;
		19'b1000111010100111010: color_data = Z;
		19'b1000111010100111011: color_data = Z;
		19'b1000111010100111100: color_data = Z;
		19'b1000111010100111101: color_data = Z;
		19'b1000111010100111110: color_data = Z;
		19'b1000111010100111111: color_data = Z;
		19'b1000111010101000000: color_data = Z;
		19'b1000111010101000001: color_data = Z;
		19'b1000111010101000010: color_data = Z;
		19'b1000111010101000011: color_data = Z;
		19'b1000111010101000100: color_data = Z;
		19'b1000111010101000101: color_data = Z;
		19'b1000111010101000110: color_data = Z;
		19'b1000111010101000111: color_data = Z;
		19'b1000111010101001000: color_data = Z;
		19'b1000111010101001001: color_data = Z;
		19'b1000111010101001010: color_data = Z;
		19'b1000111010101001011: color_data = Z;
		19'b1000111010101001100: color_data = Z;
		19'b1000111010101001101: color_data = Z;
		19'b1000111010101001110: color_data = Z;
		19'b1000111010101001111: color_data = Z;
		19'b1000111010101010000: color_data = Z;
		19'b1000111010101010001: color_data = Z;
		19'b1000111010101010010: color_data = Z;
		19'b1000111010101010011: color_data = Z;
		19'b1000111010101010100: color_data = Z;
		19'b1000111010101010101: color_data = Z;
		19'b1000111010101010110: color_data = Z;
		19'b1000111010101010111: color_data = Z;
		19'b1000111010101011000: color_data = Z;
		19'b1000111010101011001: color_data = Z;
		19'b1000111010101011010: color_data = Z;
		19'b1000111010101011011: color_data = Z;
		19'b1000111010101011100: color_data = Z;
		19'b1000111010101011101: color_data = Z;
		19'b1000111010101011110: color_data = Z;
		19'b1000111010101011111: color_data = Z;
		19'b1000111010101100000: color_data = Z;
		19'b1000111010101100001: color_data = Z;
		19'b1000111010101100010: color_data = Z;
		19'b1000111010101100011: color_data = Z;
		19'b1000111010101100100: color_data = Z;
		19'b1000111010101100101: color_data = Z;
		19'b1000111010101100110: color_data = Z;
		19'b1000111010101100111: color_data = Z;
		19'b1000111010101101000: color_data = Z;
		19'b1000111010101101001: color_data = Z;
		19'b1000111010101101010: color_data = Z;
		19'b1000111010101101011: color_data = Z;
		19'b1000111010101101100: color_data = Z;
		19'b1000111010101101101: color_data = Z;
		19'b1000111010101101110: color_data = Z;
		19'b1000111010101101111: color_data = Z;
		19'b1000111010101110000: color_data = Z;
		19'b1000111010101110001: color_data = Z;
		19'b1000111010101110010: color_data = Z;
		19'b1000111010101110011: color_data = Z;
		19'b1000111010101110100: color_data = Z;
		19'b1000111010101110101: color_data = Z;
		19'b1000111010101110110: color_data = Z;
		19'b1000111010101110111: color_data = Z;
		19'b1000111010101111000: color_data = Z;
		19'b1000111010101111001: color_data = Z;
		19'b1000111010101111010: color_data = Z;
		19'b1000111010101111011: color_data = Z;
		19'b1000111010101111100: color_data = Z;
		19'b1000111010101111101: color_data = Z;
		19'b1000111010101111110: color_data = Z;
		19'b1000111010101111111: color_data = Z;
		19'b1000111010110000000: color_data = Z;
		19'b1000111010110000001: color_data = Z;
		19'b1000111010110000010: color_data = Z;
		19'b1000111010110000011: color_data = Z;
		19'b1000111010110000100: color_data = Z;
		19'b1000111010110000101: color_data = Z;
		19'b1000111010110101010: color_data = Z;
		19'b1000111010110101011: color_data = Z;
		19'b1000111010110101100: color_data = Z;
		19'b1000111010110101101: color_data = Z;
		19'b1000111010110101110: color_data = Z;
		19'b1000111010110101111: color_data = Z;
		19'b1000111010110110000: color_data = Z;
		19'b1000111010110110001: color_data = Z;
		19'b1000111010110110010: color_data = Z;
		19'b1000111010110110011: color_data = Z;
		19'b1000111010110110100: color_data = Z;
		19'b1000111010110110101: color_data = Z;
		19'b1000111010110110110: color_data = Z;
		19'b1000111010110110111: color_data = Z;
		19'b1000111010110111000: color_data = Z;
		19'b1000111010110111001: color_data = Z;
		19'b1000111010110111010: color_data = Z;
		19'b1000111010110111011: color_data = Z;
		19'b1000111010110111100: color_data = Z;
		19'b1000111010110111101: color_data = Z;
		19'b1000111010111001001: color_data = Z;
		19'b1000111010111001010: color_data = Z;
		19'b1000111010111001011: color_data = Z;
		19'b1000111010111001100: color_data = Z;
		19'b1000111010111001101: color_data = Z;
		19'b1000111100011010100: color_data = Z;
		19'b1000111100011010101: color_data = Z;
		19'b1000111100011010110: color_data = Z;
		19'b1000111100011010111: color_data = Z;
		19'b1000111100011011000: color_data = Z;
		19'b1000111100011011001: color_data = Z;
		19'b1000111100011011010: color_data = Z;
		19'b1000111100011011011: color_data = Z;
		19'b1000111100011011100: color_data = Z;
		19'b1000111100011011101: color_data = Z;
		19'b1000111100011011110: color_data = Z;
		19'b1000111100011011111: color_data = Z;
		19'b1000111100011100000: color_data = Z;
		19'b1000111100011100001: color_data = Z;
		19'b1000111100011100010: color_data = Z;
		19'b1000111100011100011: color_data = Z;
		19'b1000111100011100100: color_data = Z;
		19'b1000111100011100101: color_data = Z;
		19'b1000111100011100110: color_data = Z;
		19'b1000111100011100111: color_data = Z;
		19'b1000111100011101000: color_data = Z;
		19'b1000111100011101001: color_data = Z;
		19'b1000111100011101010: color_data = Z;
		19'b1000111100011101011: color_data = Z;
		19'b1000111100011101100: color_data = Z;
		19'b1000111100011101101: color_data = Z;
		19'b1000111100011101110: color_data = Z;
		19'b1000111100011101111: color_data = Z;
		19'b1000111100011110000: color_data = Z;
		19'b1000111100011110001: color_data = Z;
		19'b1000111100011110010: color_data = Z;
		19'b1000111100011110011: color_data = Z;
		19'b1000111100011110100: color_data = Z;
		19'b1000111100011110101: color_data = Z;
		19'b1000111100011110110: color_data = Z;
		19'b1000111100011110111: color_data = Z;
		19'b1000111100011111000: color_data = Z;
		19'b1000111100011111001: color_data = Z;
		19'b1000111100011111010: color_data = Z;
		19'b1000111100011111011: color_data = Z;
		19'b1000111100011111100: color_data = Z;
		19'b1000111100011111101: color_data = Z;
		19'b1000111100011111110: color_data = Z;
		19'b1000111100011111111: color_data = Z;
		19'b1000111100100000000: color_data = Z;
		19'b1000111100100000001: color_data = Z;
		19'b1000111100100000010: color_data = Z;
		19'b1000111100100000011: color_data = Z;
		19'b1000111100100000100: color_data = Z;
		19'b1000111100100000101: color_data = Z;
		19'b1000111100100000110: color_data = Z;
		19'b1000111100100000111: color_data = Z;
		19'b1000111100100001000: color_data = Z;
		19'b1000111100100001001: color_data = Z;
		19'b1000111100100001010: color_data = Z;
		19'b1000111100100001011: color_data = Z;
		19'b1000111100100001100: color_data = Z;
		19'b1000111100100001101: color_data = Z;
		19'b1000111100100001110: color_data = Z;
		19'b1000111100100001111: color_data = Z;
		19'b1000111100100010000: color_data = Z;
		19'b1000111100100010001: color_data = Z;
		19'b1000111100100010010: color_data = Z;
		19'b1000111100100010011: color_data = Z;
		19'b1000111100100010100: color_data = Z;
		19'b1000111100100010101: color_data = Z;
		19'b1000111100100010110: color_data = Z;
		19'b1000111100100010111: color_data = Z;
		19'b1000111100100011000: color_data = Z;
		19'b1000111100100011001: color_data = Z;
		19'b1000111100100011010: color_data = Z;
		19'b1000111100100011011: color_data = Z;
		19'b1000111100100011100: color_data = Z;
		19'b1000111100100011101: color_data = Z;
		19'b1000111100100011110: color_data = Z;
		19'b1000111100100011111: color_data = Z;
		19'b1000111100100100000: color_data = Z;
		19'b1000111100100100001: color_data = Z;
		19'b1000111100100100010: color_data = Z;
		19'b1000111100100100011: color_data = Z;
		19'b1000111100100100100: color_data = Z;
		19'b1000111100100100101: color_data = Z;
		19'b1000111100100100110: color_data = Z;
		19'b1000111100100100111: color_data = Z;
		19'b1000111100100101000: color_data = Z;
		19'b1000111100100101001: color_data = Z;
		19'b1000111100100101010: color_data = Z;
		19'b1000111100100101011: color_data = Z;
		19'b1000111100100101100: color_data = Z;
		19'b1000111100100101101: color_data = Z;
		19'b1000111100100101110: color_data = Z;
		19'b1000111100100101111: color_data = Z;
		19'b1000111100100110000: color_data = Z;
		19'b1000111100100110001: color_data = Z;
		19'b1000111100100110010: color_data = Z;
		19'b1000111100100110011: color_data = Z;
		19'b1000111100100110100: color_data = Z;
		19'b1000111100100110101: color_data = Z;
		19'b1000111100100110110: color_data = Z;
		19'b1000111100100110111: color_data = Z;
		19'b1000111100100111000: color_data = Z;
		19'b1000111100100111001: color_data = Z;
		19'b1000111100100111010: color_data = Z;
		19'b1000111100100111011: color_data = Z;
		19'b1000111100100111100: color_data = Z;
		19'b1000111100100111101: color_data = Z;
		19'b1000111100100111110: color_data = Z;
		19'b1000111100100111111: color_data = Z;
		19'b1000111100101000000: color_data = Z;
		19'b1000111100101000001: color_data = Z;
		19'b1000111100101000010: color_data = Z;
		19'b1000111100101000011: color_data = Z;
		19'b1000111100101000100: color_data = Z;
		19'b1000111100101000101: color_data = Z;
		19'b1000111100101000110: color_data = Z;
		19'b1000111100101000111: color_data = Z;
		19'b1000111100101001000: color_data = Z;
		19'b1000111100101001001: color_data = Z;
		19'b1000111100101001010: color_data = Z;
		19'b1000111100101001011: color_data = Z;
		19'b1000111100101001100: color_data = Z;
		19'b1000111100101001101: color_data = Z;
		19'b1000111100101001110: color_data = Z;
		19'b1000111100101001111: color_data = Z;
		19'b1000111100101010000: color_data = Z;
		19'b1000111100101010001: color_data = Z;
		19'b1000111100101010010: color_data = Z;
		19'b1000111100101010011: color_data = Z;
		19'b1000111100101010100: color_data = Z;
		19'b1000111100101010101: color_data = Z;
		19'b1000111100101010110: color_data = Z;
		19'b1000111100101010111: color_data = Z;
		19'b1000111100101011000: color_data = Z;
		19'b1000111100101011001: color_data = Z;
		19'b1000111100101011010: color_data = Z;
		19'b1000111100101011011: color_data = Z;
		19'b1000111100101011100: color_data = Z;
		19'b1000111100101011101: color_data = Z;
		19'b1000111100101011110: color_data = Z;
		19'b1000111100101011111: color_data = Z;
		19'b1000111100101100000: color_data = Z;
		19'b1000111100101100001: color_data = Z;
		19'b1000111100101100010: color_data = Z;
		19'b1000111100101100011: color_data = Z;
		19'b1000111100101100100: color_data = Z;
		19'b1000111100101100101: color_data = Z;
		19'b1000111100101100110: color_data = Z;
		19'b1000111100101100111: color_data = Z;
		19'b1000111100101101000: color_data = Z;
		19'b1000111100101101001: color_data = Z;
		19'b1000111100101101010: color_data = Z;
		19'b1000111100101101011: color_data = Z;
		19'b1000111100101101100: color_data = Z;
		19'b1000111100101101101: color_data = Z;
		19'b1000111100101101110: color_data = Z;
		19'b1000111100101101111: color_data = Z;
		19'b1000111100101110000: color_data = Z;
		19'b1000111100101110001: color_data = Z;
		19'b1000111100101110010: color_data = Z;
		19'b1000111100101110011: color_data = Z;
		19'b1000111100101110100: color_data = Z;
		19'b1000111100101110101: color_data = Z;
		19'b1000111100101110110: color_data = Z;
		19'b1000111100101110111: color_data = Z;
		19'b1000111100101111000: color_data = Z;
		19'b1000111100101111001: color_data = Z;
		19'b1000111100101111010: color_data = Z;
		19'b1000111100101111011: color_data = Z;
		19'b1000111100101111100: color_data = Z;
		19'b1000111100101111101: color_data = Z;
		19'b1000111100101111110: color_data = Z;
		19'b1000111100101111111: color_data = Z;
		19'b1000111100110000000: color_data = Z;
		19'b1000111100110101011: color_data = Z;
		19'b1000111100110101100: color_data = Z;
		19'b1000111100110101101: color_data = Z;
		19'b1000111100110101110: color_data = Z;
		19'b1000111100110101111: color_data = Z;
		19'b1000111100110110000: color_data = Z;
		19'b1000111100110110001: color_data = Z;
		19'b1000111100110110010: color_data = Z;
		19'b1000111100110110011: color_data = Z;
		19'b1000111100110110100: color_data = Z;
		19'b1000111100110110101: color_data = Z;
		19'b1000111100110110110: color_data = Z;
		19'b1000111100110111000: color_data = Z;
		19'b1000111100110111001: color_data = Z;
		19'b1000111100110111010: color_data = Z;
		19'b1000111100110111011: color_data = Z;
		19'b1000111100110111100: color_data = Z;
		19'b1000111100110111101: color_data = Z;
		19'b1000111100111001001: color_data = Z;
		19'b1000111100111001010: color_data = Z;
		19'b1000111100111001011: color_data = Z;
		19'b1000111100111001100: color_data = Z;
		19'b1000111100111001101: color_data = Z;
		19'b1000111110011010110: color_data = Z;
		19'b1000111110011010111: color_data = Z;
		19'b1000111110011011000: color_data = Z;
		19'b1000111110011011001: color_data = Z;
		19'b1000111110011011010: color_data = Z;
		19'b1000111110011011011: color_data = Z;
		19'b1000111110011011100: color_data = Z;
		19'b1000111110011011101: color_data = Z;
		19'b1000111110011011110: color_data = Z;
		19'b1000111110011011111: color_data = Z;
		19'b1000111110011100000: color_data = Z;
		19'b1000111110011100001: color_data = Z;
		19'b1000111110011100010: color_data = Z;
		19'b1000111110011100011: color_data = Z;
		19'b1000111110011100100: color_data = Z;
		19'b1000111110011100101: color_data = Z;
		19'b1000111110011100110: color_data = Z;
		19'b1000111110011100111: color_data = Z;
		19'b1000111110011101000: color_data = Z;
		19'b1000111110011101001: color_data = Z;
		19'b1000111110011101010: color_data = Z;
		19'b1000111110011101011: color_data = Z;
		19'b1000111110011101100: color_data = Z;
		19'b1000111110011101101: color_data = Z;
		19'b1000111110011101110: color_data = Z;
		19'b1000111110011101111: color_data = Z;
		19'b1000111110011110000: color_data = Z;
		19'b1000111110011110001: color_data = Z;
		19'b1000111110011111010: color_data = Z;
		19'b1000111110011111011: color_data = Z;
		19'b1000111110011111100: color_data = Z;
		19'b1000111110011111101: color_data = Z;
		19'b1000111110011111110: color_data = Z;
		19'b1000111110011111111: color_data = Z;
		19'b1000111110100000000: color_data = Z;
		19'b1000111110100000001: color_data = Z;
		19'b1000111110100000010: color_data = Z;
		19'b1000111110100000011: color_data = Z;
		19'b1000111110100000100: color_data = Z;
		19'b1000111110100000101: color_data = Z;
		19'b1000111110100000110: color_data = Z;
		19'b1000111110100000111: color_data = Z;
		19'b1000111110100001000: color_data = Z;
		19'b1000111110100001001: color_data = Z;
		19'b1000111110100001010: color_data = Z;
		19'b1000111110100001011: color_data = Z;
		19'b1000111110100001100: color_data = Z;
		19'b1000111110100001101: color_data = Z;
		19'b1000111110100001110: color_data = Z;
		19'b1000111110100001111: color_data = Z;
		19'b1000111110100010000: color_data = Z;
		19'b1000111110100010001: color_data = Z;
		19'b1000111110100010010: color_data = Z;
		19'b1000111110100010011: color_data = Z;
		19'b1000111110100010100: color_data = Z;
		19'b1000111110100010101: color_data = Z;
		19'b1000111110100010110: color_data = Z;
		19'b1000111110100010111: color_data = Z;
		19'b1000111110100011000: color_data = Z;
		19'b1000111110100011001: color_data = Z;
		19'b1000111110100011010: color_data = Z;
		19'b1000111110100011011: color_data = Z;
		19'b1000111110100011100: color_data = Z;
		19'b1000111110100011101: color_data = Z;
		19'b1000111110100011110: color_data = Z;
		19'b1000111110100011111: color_data = Z;
		19'b1000111110100100000: color_data = Z;
		19'b1000111110100100001: color_data = Z;
		19'b1000111110100100010: color_data = Z;
		19'b1000111110100100011: color_data = Z;
		19'b1000111110100100100: color_data = Z;
		19'b1000111110100100101: color_data = Z;
		19'b1000111110100100110: color_data = Z;
		19'b1000111110100100111: color_data = Z;
		19'b1000111110100101000: color_data = Z;
		19'b1000111110100101001: color_data = Z;
		19'b1000111110100101010: color_data = Z;
		19'b1000111110100101011: color_data = Z;
		19'b1000111110100101100: color_data = Z;
		19'b1000111110100101101: color_data = Z;
		19'b1000111110100101110: color_data = Z;
		19'b1000111110100101111: color_data = Z;
		19'b1000111110100110000: color_data = Z;
		19'b1000111110100110001: color_data = Z;
		19'b1000111110100110010: color_data = Z;
		19'b1000111110100110011: color_data = Z;
		19'b1000111110100110100: color_data = Z;
		19'b1000111110100110101: color_data = Z;
		19'b1000111110100110110: color_data = Z;
		19'b1000111110100110111: color_data = Z;
		19'b1000111110100111000: color_data = Z;
		19'b1000111110100111001: color_data = Z;
		19'b1000111110100111010: color_data = Z;
		19'b1000111110100111011: color_data = Z;
		19'b1000111110100111100: color_data = Z;
		19'b1000111110100111101: color_data = Z;
		19'b1000111110100111110: color_data = Z;
		19'b1000111110100111111: color_data = Z;
		19'b1000111110101000000: color_data = Z;
		19'b1000111110101000001: color_data = Z;
		19'b1000111110101000010: color_data = Z;
		19'b1000111110101000011: color_data = Z;
		19'b1000111110101000100: color_data = Z;
		19'b1000111110101000101: color_data = Z;
		19'b1000111110101000110: color_data = Z;
		19'b1000111110101000111: color_data = Z;
		19'b1000111110101001000: color_data = Z;
		19'b1000111110101001001: color_data = Z;
		19'b1000111110101001010: color_data = Z;
		19'b1000111110101001011: color_data = Z;
		19'b1000111110101001100: color_data = Z;
		19'b1000111110101001101: color_data = Z;
		19'b1000111110101001110: color_data = Z;
		19'b1000111110101001111: color_data = Z;
		19'b1000111110101010000: color_data = Z;
		19'b1000111110101010001: color_data = Z;
		19'b1000111110101010010: color_data = Z;
		19'b1000111110101010011: color_data = Z;
		19'b1000111110101010100: color_data = Z;
		19'b1000111110101010101: color_data = Z;
		19'b1000111110101010110: color_data = Z;
		19'b1000111110101010111: color_data = Z;
		19'b1000111110101011000: color_data = Z;
		19'b1000111110101011001: color_data = Z;
		19'b1000111110101011010: color_data = Z;
		19'b1000111110101011011: color_data = Z;
		19'b1000111110101011100: color_data = Z;
		19'b1000111110101011101: color_data = Z;
		19'b1000111110101011110: color_data = Z;
		19'b1000111110101011111: color_data = Z;
		19'b1000111110101100000: color_data = Z;
		19'b1000111110101100001: color_data = Z;
		19'b1000111110101100010: color_data = Z;
		19'b1000111110101100011: color_data = Z;
		19'b1000111110101100100: color_data = Z;
		19'b1000111110101100101: color_data = Z;
		19'b1000111110101100110: color_data = Z;
		19'b1000111110101100111: color_data = Z;
		19'b1000111110101101000: color_data = Z;
		19'b1000111110101101001: color_data = Z;
		19'b1000111110101101010: color_data = Z;
		19'b1000111110101101011: color_data = Z;
		19'b1000111110101101100: color_data = Z;
		19'b1000111110101101101: color_data = Z;
		19'b1000111110101101110: color_data = Z;
		19'b1000111110101101111: color_data = Z;
		19'b1000111110101110000: color_data = Z;
		19'b1000111110101110001: color_data = Z;
		19'b1000111110101110010: color_data = Z;
		19'b1000111110101110011: color_data = Z;
		19'b1000111110101110100: color_data = Z;
		19'b1000111110101110101: color_data = Z;
		19'b1000111110101110110: color_data = Z;
		19'b1000111110101110111: color_data = Z;
		19'b1000111110101111000: color_data = Z;
		19'b1000111110101111001: color_data = Z;
		19'b1000111110101111010: color_data = Z;
		19'b1000111110101111011: color_data = Z;
		19'b1000111110110101100: color_data = Z;
		19'b1000111110110101101: color_data = Z;
		19'b1000111110110101110: color_data = Z;
		19'b1000111110110101111: color_data = Z;
		19'b1000111110110110000: color_data = Z;
		19'b1000111110110110001: color_data = Z;
		19'b1000111110110110010: color_data = Z;
		19'b1000111110110110011: color_data = Z;
		19'b1000111110110110100: color_data = Z;
		19'b1000111110110110101: color_data = Z;
		19'b1000111110110110110: color_data = Z;
		19'b1000111110110111000: color_data = Z;
		19'b1000111110110111001: color_data = Z;
		19'b1000111110110111010: color_data = Z;
		19'b1000111110110111011: color_data = Z;
		19'b1000111110110111100: color_data = Z;
		19'b1000111110111001001: color_data = Z;
		19'b1000111110111001010: color_data = Z;
		19'b1000111110111001011: color_data = Z;
		19'b1000111110111001100: color_data = Z;
		19'b1000111110111001101: color_data = Z;
		19'b1001000000011010110: color_data = Z;
		19'b1001000000011010111: color_data = Z;
		19'b1001000000011011000: color_data = Z;
		19'b1001000000011011001: color_data = Z;
		19'b1001000000011011010: color_data = Z;
		19'b1001000000011011011: color_data = Z;
		19'b1001000000011011100: color_data = Z;
		19'b1001000000011011101: color_data = Z;
		19'b1001000000011011110: color_data = Z;
		19'b1001000000011011111: color_data = Z;
		19'b1001000000011100000: color_data = Z;
		19'b1001000000011100001: color_data = Z;
		19'b1001000000011100010: color_data = Z;
		19'b1001000000011100011: color_data = Z;
		19'b1001000000011100100: color_data = Z;
		19'b1001000000011100101: color_data = Z;
		19'b1001000000011100110: color_data = Z;
		19'b1001000000011100111: color_data = Z;
		19'b1001000000011101000: color_data = Z;
		19'b1001000000011101001: color_data = Z;
		19'b1001000000011101010: color_data = Z;
		19'b1001000000011101100: color_data = Z;
		19'b1001000000011101101: color_data = Z;
		19'b1001000000011101110: color_data = Z;
		19'b1001000000011101111: color_data = Z;
		19'b1001000000011110000: color_data = Z;
		19'b1001000000011110001: color_data = Z;
		19'b1001000000011110011: color_data = Z;
		19'b1001000000011110100: color_data = Z;
		19'b1001000000011111110: color_data = Z;
		19'b1001000000011111111: color_data = Z;
		19'b1001000000100000000: color_data = Z;
		19'b1001000000100000001: color_data = Z;
		19'b1001000000100000010: color_data = Z;
		19'b1001000000100000011: color_data = Z;
		19'b1001000000100000100: color_data = Z;
		19'b1001000000100000101: color_data = Z;
		19'b1001000000100000110: color_data = Z;
		19'b1001000000100000111: color_data = Z;
		19'b1001000000100001000: color_data = Z;
		19'b1001000000100001001: color_data = Z;
		19'b1001000000100001010: color_data = Z;
		19'b1001000000100001011: color_data = Z;
		19'b1001000000100001100: color_data = Z;
		19'b1001000000100001101: color_data = Z;
		19'b1001000000100001110: color_data = Z;
		19'b1001000000100001111: color_data = Z;
		19'b1001000000100010000: color_data = Z;
		19'b1001000000100010001: color_data = Z;
		19'b1001000000100010010: color_data = Z;
		19'b1001000000100010011: color_data = Z;
		19'b1001000000100010100: color_data = Z;
		19'b1001000000100010101: color_data = Z;
		19'b1001000000100010110: color_data = Z;
		19'b1001000000100010111: color_data = Z;
		19'b1001000000100011000: color_data = Z;
		19'b1001000000100011001: color_data = Z;
		19'b1001000000100011010: color_data = Z;
		19'b1001000000100011011: color_data = Z;
		19'b1001000000100011100: color_data = Z;
		19'b1001000000100011101: color_data = Z;
		19'b1001000000100011110: color_data = Z;
		19'b1001000000100011111: color_data = Z;
		19'b1001000000100100000: color_data = Z;
		19'b1001000000100100001: color_data = Z;
		19'b1001000000100100010: color_data = Z;
		19'b1001000000100100011: color_data = Z;
		19'b1001000000100100100: color_data = Z;
		19'b1001000000100100101: color_data = Z;
		19'b1001000000100100110: color_data = Z;
		19'b1001000000100100111: color_data = Z;
		19'b1001000000100101000: color_data = Z;
		19'b1001000000100101001: color_data = Z;
		19'b1001000000100101010: color_data = Z;
		19'b1001000000100101011: color_data = Z;
		19'b1001000000100101100: color_data = Z;
		19'b1001000000100101101: color_data = Z;
		19'b1001000000100101110: color_data = Z;
		19'b1001000000100101111: color_data = Z;
		19'b1001000000100110000: color_data = Z;
		19'b1001000000100110001: color_data = Z;
		19'b1001000000100110010: color_data = Z;
		19'b1001000000100110011: color_data = Z;
		19'b1001000000100110100: color_data = Z;
		19'b1001000000100110101: color_data = Z;
		19'b1001000000100110110: color_data = Z;
		19'b1001000000100110111: color_data = Z;
		19'b1001000000100111000: color_data = Z;
		19'b1001000000100111001: color_data = Z;
		19'b1001000000100111010: color_data = Z;
		19'b1001000000100111011: color_data = Z;
		19'b1001000000100111100: color_data = Z;
		19'b1001000000100111101: color_data = Z;
		19'b1001000000100111110: color_data = Z;
		19'b1001000000100111111: color_data = Z;
		19'b1001000000101000000: color_data = Z;
		19'b1001000000101000001: color_data = Z;
		19'b1001000000101000010: color_data = Z;
		19'b1001000000101000011: color_data = Z;
		19'b1001000000101000100: color_data = Z;
		19'b1001000000101000101: color_data = Z;
		19'b1001000000101000110: color_data = Z;
		19'b1001000000101000111: color_data = Z;
		19'b1001000000101001000: color_data = Z;
		19'b1001000000101001001: color_data = Z;
		19'b1001000000101001010: color_data = Z;
		19'b1001000000101001011: color_data = Z;
		19'b1001000000101001100: color_data = Z;
		19'b1001000000101001101: color_data = Z;
		19'b1001000000101001110: color_data = Z;
		19'b1001000000101001111: color_data = Z;
		19'b1001000000101010000: color_data = Z;
		19'b1001000000101010001: color_data = Z;
		19'b1001000000101010010: color_data = Z;
		19'b1001000000101010011: color_data = Z;
		19'b1001000000101010100: color_data = Z;
		19'b1001000000101010101: color_data = Z;
		19'b1001000000101010110: color_data = Z;
		19'b1001000000101010111: color_data = Z;
		19'b1001000000101011000: color_data = Z;
		19'b1001000000101011001: color_data = Z;
		19'b1001000000101011010: color_data = Z;
		19'b1001000000101011011: color_data = Z;
		19'b1001000000101011100: color_data = Z;
		19'b1001000000101011101: color_data = Z;
		19'b1001000000101011110: color_data = Z;
		19'b1001000000101011111: color_data = Z;
		19'b1001000000101100000: color_data = Z;
		19'b1001000000101100001: color_data = Z;
		19'b1001000000101100010: color_data = Z;
		19'b1001000000101100011: color_data = Z;
		19'b1001000000101100100: color_data = Z;
		19'b1001000000101100101: color_data = Z;
		19'b1001000000101100110: color_data = Z;
		19'b1001000000101100111: color_data = Z;
		19'b1001000000101101000: color_data = Z;
		19'b1001000000101101001: color_data = Z;
		19'b1001000000101101010: color_data = Z;
		19'b1001000000101101011: color_data = Z;
		19'b1001000000101101100: color_data = Z;
		19'b1001000000101101101: color_data = Z;
		19'b1001000000101101110: color_data = Z;
		19'b1001000000101101111: color_data = Z;
		19'b1001000000101110000: color_data = Z;
		19'b1001000000101110001: color_data = Z;
		19'b1001000000101110010: color_data = Z;
		19'b1001000000101110011: color_data = Z;
		19'b1001000000101110100: color_data = Z;
		19'b1001000000101110101: color_data = Z;
		19'b1001000000101110110: color_data = Z;
		19'b1001000000101110111: color_data = Z;
		19'b1001000000101111000: color_data = Z;
		19'b1001000000101111001: color_data = Z;
		19'b1001000000110101100: color_data = Z;
		19'b1001000000110101101: color_data = Z;
		19'b1001000000110101110: color_data = Z;
		19'b1001000000110101111: color_data = Z;
		19'b1001000000110110000: color_data = Z;
		19'b1001000000110110001: color_data = Z;
		19'b1001000000110110010: color_data = Z;
		19'b1001000000110110011: color_data = Z;
		19'b1001000000110110100: color_data = Z;
		19'b1001000000110110101: color_data = Z;
		19'b1001000000110110110: color_data = Z;
		19'b1001000000110111000: color_data = Z;
		19'b1001000000110111001: color_data = Z;
		19'b1001000000110111010: color_data = Z;
		19'b1001000000110111011: color_data = Z;
		19'b1001000000111001001: color_data = Z;
		19'b1001000000111001010: color_data = Z;
		19'b1001000000111001011: color_data = Z;
		19'b1001000000111001100: color_data = Z;
		19'b1001000000111001101: color_data = Z;
		19'b1001000010011010110: color_data = Z;
		19'b1001000010011010111: color_data = Z;
		19'b1001000010011011000: color_data = Z;
		19'b1001000010011011001: color_data = Z;
		19'b1001000010011011010: color_data = Z;
		19'b1001000010011011011: color_data = Z;
		19'b1001000010011011100: color_data = Z;
		19'b1001000010011011101: color_data = Z;
		19'b1001000010011011110: color_data = Z;
		19'b1001000010011011111: color_data = Z;
		19'b1001000010011100000: color_data = Z;
		19'b1001000010011100001: color_data = Z;
		19'b1001000010011100010: color_data = Z;
		19'b1001000010011100011: color_data = Z;
		19'b1001000010011100100: color_data = Z;
		19'b1001000010011100101: color_data = Z;
		19'b1001000010011100110: color_data = Z;
		19'b1001000010011100111: color_data = Z;
		19'b1001000010011101000: color_data = Z;
		19'b1001000010011101001: color_data = Z;
		19'b1001000010011101100: color_data = Z;
		19'b1001000010011101101: color_data = Z;
		19'b1001000010011101110: color_data = Z;
		19'b1001000010011101111: color_data = Z;
		19'b1001000010011110000: color_data = Z;
		19'b1001000010011110001: color_data = Z;
		19'b1001000010011110010: color_data = Z;
		19'b1001000010011110011: color_data = Z;
		19'b1001000010011110100: color_data = Z;
		19'b1001000010011110101: color_data = Z;
		19'b1001000010011110110: color_data = Z;
		19'b1001000010100001001: color_data = Z;
		19'b1001000010100001010: color_data = Z;
		19'b1001000010100001011: color_data = Z;
		19'b1001000010100001100: color_data = Z;
		19'b1001000010100001101: color_data = Z;
		19'b1001000010100001110: color_data = Z;
		19'b1001000010100001111: color_data = Z;
		19'b1001000010100010000: color_data = Z;
		19'b1001000010100010001: color_data = Z;
		19'b1001000010100010010: color_data = Z;
		19'b1001000010100010011: color_data = Z;
		19'b1001000010100010100: color_data = Z;
		19'b1001000010100010101: color_data = Z;
		19'b1001000010100010110: color_data = Z;
		19'b1001000010100010111: color_data = Z;
		19'b1001000010100011000: color_data = Z;
		19'b1001000010100011001: color_data = Z;
		19'b1001000010100011010: color_data = Z;
		19'b1001000010100011011: color_data = Z;
		19'b1001000010100011100: color_data = Z;
		19'b1001000010100011101: color_data = Z;
		19'b1001000010100011110: color_data = Z;
		19'b1001000010100011111: color_data = Z;
		19'b1001000010100100000: color_data = Z;
		19'b1001000010100100001: color_data = Z;
		19'b1001000010100100010: color_data = Z;
		19'b1001000010100100011: color_data = Z;
		19'b1001000010100100100: color_data = Z;
		19'b1001000010100100101: color_data = Z;
		19'b1001000010100100110: color_data = Z;
		19'b1001000010100100111: color_data = Z;
		19'b1001000010100101000: color_data = Z;
		19'b1001000010100101001: color_data = Z;
		19'b1001000010100101010: color_data = Z;
		19'b1001000010100101011: color_data = Z;
		19'b1001000010100101100: color_data = Z;
		19'b1001000010100101101: color_data = Z;
		19'b1001000010100101110: color_data = Z;
		19'b1001000010100101111: color_data = Z;
		19'b1001000010100110000: color_data = Z;
		19'b1001000010100110001: color_data = Z;
		19'b1001000010100110010: color_data = Z;
		19'b1001000010100110011: color_data = Z;
		19'b1001000010100110100: color_data = Z;
		19'b1001000010100110101: color_data = Z;
		19'b1001000010100110110: color_data = Z;
		19'b1001000010100110111: color_data = Z;
		19'b1001000010100111000: color_data = Z;
		19'b1001000010100111001: color_data = Z;
		19'b1001000010100111010: color_data = Z;
		19'b1001000010100111011: color_data = Z;
		19'b1001000010100111100: color_data = Z;
		19'b1001000010100111101: color_data = Z;
		19'b1001000010100111110: color_data = Z;
		19'b1001000010100111111: color_data = Z;
		19'b1001000010101000000: color_data = Z;
		19'b1001000010101000001: color_data = Z;
		19'b1001000010101000010: color_data = Z;
		19'b1001000010101000011: color_data = Z;
		19'b1001000010101000100: color_data = Z;
		19'b1001000010101000101: color_data = Z;
		19'b1001000010101000110: color_data = Z;
		19'b1001000010101000111: color_data = Z;
		19'b1001000010101001000: color_data = Z;
		19'b1001000010101001001: color_data = Z;
		19'b1001000010101001010: color_data = Z;
		19'b1001000010101001011: color_data = Z;
		19'b1001000010101001100: color_data = Z;
		19'b1001000010101001101: color_data = Z;
		19'b1001000010101001110: color_data = Z;
		19'b1001000010101001111: color_data = Z;
		19'b1001000010101010000: color_data = Z;
		19'b1001000010101010001: color_data = Z;
		19'b1001000010101010010: color_data = Z;
		19'b1001000010101010011: color_data = Z;
		19'b1001000010101010100: color_data = Z;
		19'b1001000010101010101: color_data = Z;
		19'b1001000010101010110: color_data = Z;
		19'b1001000010101010111: color_data = Z;
		19'b1001000010101011000: color_data = Z;
		19'b1001000010101011001: color_data = Z;
		19'b1001000010101011010: color_data = Z;
		19'b1001000010101011011: color_data = Z;
		19'b1001000010101011100: color_data = Z;
		19'b1001000010101011101: color_data = Z;
		19'b1001000010101011110: color_data = Z;
		19'b1001000010101011111: color_data = Z;
		19'b1001000010101100000: color_data = Z;
		19'b1001000010101100001: color_data = Z;
		19'b1001000010101100010: color_data = Z;
		19'b1001000010101100011: color_data = Z;
		19'b1001000010101100100: color_data = Z;
		19'b1001000010101100101: color_data = Z;
		19'b1001000010101100110: color_data = Z;
		19'b1001000010101100111: color_data = Z;
		19'b1001000010101101000: color_data = Z;
		19'b1001000010101101001: color_data = Z;
		19'b1001000010101101010: color_data = Z;
		19'b1001000010101101011: color_data = Z;
		19'b1001000010101101100: color_data = Z;
		19'b1001000010101101101: color_data = Z;
		19'b1001000010101101110: color_data = Z;
		19'b1001000010101101111: color_data = Z;
		19'b1001000010101110000: color_data = Z;
		19'b1001000010101110001: color_data = Z;
		19'b1001000010101110010: color_data = Z;
		19'b1001000010101110011: color_data = Z;
		19'b1001000010101110100: color_data = Z;
		19'b1001000010101110101: color_data = Z;
		19'b1001000010101110110: color_data = Z;
		19'b1001000010101110111: color_data = Z;
		19'b1001000010110101101: color_data = Z;
		19'b1001000010110101110: color_data = Z;
		19'b1001000010110101111: color_data = Z;
		19'b1001000010110110000: color_data = Z;
		19'b1001000010110110001: color_data = Z;
		19'b1001000010110110010: color_data = Z;
		19'b1001000010110110011: color_data = Z;
		19'b1001000010110110100: color_data = Z;
		19'b1001000010110110101: color_data = Z;
		19'b1001000010110110110: color_data = Z;
		19'b1001000010110111001: color_data = Z;
		19'b1001000010110111010: color_data = Z;
		19'b1001000010110111011: color_data = Z;
		19'b1001000010111001000: color_data = Z;
		19'b1001000010111001001: color_data = Z;
		19'b1001000010111001010: color_data = Z;
		19'b1001000010111001011: color_data = Z;
		19'b1001000010111001100: color_data = Z;
		19'b1001000010111001101: color_data = Z;
		19'b1001000100011010110: color_data = Z;
		19'b1001000100011010111: color_data = Z;
		19'b1001000100011011000: color_data = Z;
		19'b1001000100011011001: color_data = Z;
		19'b1001000100011011010: color_data = Z;
		19'b1001000100011011011: color_data = Z;
		19'b1001000100011011100: color_data = Z;
		19'b1001000100011011101: color_data = Z;
		19'b1001000100011011110: color_data = Z;
		19'b1001000100011011111: color_data = Z;
		19'b1001000100011100000: color_data = Z;
		19'b1001000100011100001: color_data = Z;
		19'b1001000100011100010: color_data = Z;
		19'b1001000100011100011: color_data = Z;
		19'b1001000100011100100: color_data = Z;
		19'b1001000100011100101: color_data = Z;
		19'b1001000100011100110: color_data = Z;
		19'b1001000100011100111: color_data = Z;
		19'b1001000100011101000: color_data = Z;
		19'b1001000100011101011: color_data = Z;
		19'b1001000100011101100: color_data = Z;
		19'b1001000100011101101: color_data = Z;
		19'b1001000100011101110: color_data = Z;
		19'b1001000100011101111: color_data = Z;
		19'b1001000100011110000: color_data = Z;
		19'b1001000100011110001: color_data = Z;
		19'b1001000100011110010: color_data = Z;
		19'b1001000100011110011: color_data = Z;
		19'b1001000100011110100: color_data = Z;
		19'b1001000100011110101: color_data = Z;
		19'b1001000100100001100: color_data = Z;
		19'b1001000100100001101: color_data = Z;
		19'b1001000100100001110: color_data = Z;
		19'b1001000100100001111: color_data = Z;
		19'b1001000100100010001: color_data = Z;
		19'b1001000100100010010: color_data = Z;
		19'b1001000100100010011: color_data = Z;
		19'b1001000100100010100: color_data = Z;
		19'b1001000100100010101: color_data = Z;
		19'b1001000100100010110: color_data = Z;
		19'b1001000100100010111: color_data = Z;
		19'b1001000100100011000: color_data = Z;
		19'b1001000100100011001: color_data = Z;
		19'b1001000100100011010: color_data = Z;
		19'b1001000100100011011: color_data = Z;
		19'b1001000100100011100: color_data = Z;
		19'b1001000100100011101: color_data = Z;
		19'b1001000100100011110: color_data = Z;
		19'b1001000100100011111: color_data = Z;
		19'b1001000100100100000: color_data = Z;
		19'b1001000100100100001: color_data = Z;
		19'b1001000100100100010: color_data = Z;
		19'b1001000100100100011: color_data = Z;
		19'b1001000100100100100: color_data = Z;
		19'b1001000100100100101: color_data = Z;
		19'b1001000100100100110: color_data = Z;
		19'b1001000100100100111: color_data = Z;
		19'b1001000100100101000: color_data = Z;
		19'b1001000100100101001: color_data = Z;
		19'b1001000100100101010: color_data = Z;
		19'b1001000100100101011: color_data = Z;
		19'b1001000100100101100: color_data = Z;
		19'b1001000100100101101: color_data = Z;
		19'b1001000100100101110: color_data = Z;
		19'b1001000100100101111: color_data = Z;
		19'b1001000100100110000: color_data = Z;
		19'b1001000100100110001: color_data = Z;
		19'b1001000100100110010: color_data = Z;
		19'b1001000100100110011: color_data = Z;
		19'b1001000100100110100: color_data = Z;
		19'b1001000100100110101: color_data = Z;
		19'b1001000100100110110: color_data = Z;
		19'b1001000100100110111: color_data = Z;
		19'b1001000100100111000: color_data = Z;
		19'b1001000100100111001: color_data = Z;
		19'b1001000100100111010: color_data = Z;
		19'b1001000100100111011: color_data = Z;
		19'b1001000100100111100: color_data = Z;
		19'b1001000100100111101: color_data = Z;
		19'b1001000100100111110: color_data = Z;
		19'b1001000100100111111: color_data = Z;
		19'b1001000100101000000: color_data = Z;
		19'b1001000100101000001: color_data = Z;
		19'b1001000100101000010: color_data = Z;
		19'b1001000100101000011: color_data = Z;
		19'b1001000100101000100: color_data = Z;
		19'b1001000100101000101: color_data = Z;
		19'b1001000100101000110: color_data = Z;
		19'b1001000100101000111: color_data = Z;
		19'b1001000100101001000: color_data = Z;
		19'b1001000100101001001: color_data = Z;
		19'b1001000100101001010: color_data = Z;
		19'b1001000100101001011: color_data = Z;
		19'b1001000100101001100: color_data = Z;
		19'b1001000100101001101: color_data = Z;
		19'b1001000100101001110: color_data = Z;
		19'b1001000100101001111: color_data = Z;
		19'b1001000100101010000: color_data = Z;
		19'b1001000100101010001: color_data = Z;
		19'b1001000100101010010: color_data = Z;
		19'b1001000100101010011: color_data = Z;
		19'b1001000100101010100: color_data = Z;
		19'b1001000100101010101: color_data = Z;
		19'b1001000100101010110: color_data = Z;
		19'b1001000100101010111: color_data = Z;
		19'b1001000100101011000: color_data = Z;
		19'b1001000100101011001: color_data = Z;
		19'b1001000100101011010: color_data = Z;
		19'b1001000100101011011: color_data = Z;
		19'b1001000100101011100: color_data = Z;
		19'b1001000100101011101: color_data = Z;
		19'b1001000100101011110: color_data = Z;
		19'b1001000100101011111: color_data = Z;
		19'b1001000100101100000: color_data = Z;
		19'b1001000100101100001: color_data = Z;
		19'b1001000100101100010: color_data = Z;
		19'b1001000100101100011: color_data = Z;
		19'b1001000100101100100: color_data = Z;
		19'b1001000100101100101: color_data = Z;
		19'b1001000100101100110: color_data = Z;
		19'b1001000100101100111: color_data = Z;
		19'b1001000100101101000: color_data = Z;
		19'b1001000100101101001: color_data = Z;
		19'b1001000100101101010: color_data = Z;
		19'b1001000100101101011: color_data = Z;
		19'b1001000100101101100: color_data = Z;
		19'b1001000100101101101: color_data = Z;
		19'b1001000100101101110: color_data = Z;
		19'b1001000100101101111: color_data = Z;
		19'b1001000100101110000: color_data = Z;
		19'b1001000100101110001: color_data = Z;
		19'b1001000100101110010: color_data = Z;
		19'b1001000100101110011: color_data = Z;
		19'b1001000100101110100: color_data = Z;
		19'b1001000100101110101: color_data = Z;
		19'b1001000100101110110: color_data = Z;
		19'b1001000100110101101: color_data = Z;
		19'b1001000100110101110: color_data = Z;
		19'b1001000100110101111: color_data = Z;
		19'b1001000100110110000: color_data = Z;
		19'b1001000100110110001: color_data = Z;
		19'b1001000100110110010: color_data = Z;
		19'b1001000100110110011: color_data = Z;
		19'b1001000100110110100: color_data = Z;
		19'b1001000100110110101: color_data = Z;
		19'b1001000100110110110: color_data = Z;
		19'b1001000100110111001: color_data = Z;
		19'b1001000100110111010: color_data = Z;
		19'b1001000100110111011: color_data = Z;
		19'b1001000100111001000: color_data = Z;
		19'b1001000100111001001: color_data = Z;
		19'b1001000100111001010: color_data = Z;
		19'b1001000100111001011: color_data = Z;
		19'b1001000100111001100: color_data = Z;
		19'b1001000100111001101: color_data = Z;
		19'b1001000110011010101: color_data = Z;
		19'b1001000110011010110: color_data = Z;
		19'b1001000110011010111: color_data = Z;
		19'b1001000110011011000: color_data = Z;
		19'b1001000110011011001: color_data = Z;
		19'b1001000110011011010: color_data = Z;
		19'b1001000110011011011: color_data = Z;
		19'b1001000110011011100: color_data = Z;
		19'b1001000110011011101: color_data = Z;
		19'b1001000110011011110: color_data = Z;
		19'b1001000110011011111: color_data = Z;
		19'b1001000110011100000: color_data = Z;
		19'b1001000110011100001: color_data = Z;
		19'b1001000110011100010: color_data = Z;
		19'b1001000110011100011: color_data = Z;
		19'b1001000110011100100: color_data = Z;
		19'b1001000110011100101: color_data = Z;
		19'b1001000110011100110: color_data = Z;
		19'b1001000110011100111: color_data = Z;
		19'b1001000110011101011: color_data = Z;
		19'b1001000110011101100: color_data = Z;
		19'b1001000110011101101: color_data = Z;
		19'b1001000110011101110: color_data = Z;
		19'b1001000110011101111: color_data = Z;
		19'b1001000110011110001: color_data = Z;
		19'b1001000110011110010: color_data = Z;
		19'b1001000110011110011: color_data = Z;
		19'b1001000110011110100: color_data = Z;
		19'b1001000110100001110: color_data = Z;
		19'b1001000110100001111: color_data = Z;
		19'b1001000110100010111: color_data = Z;
		19'b1001000110100011000: color_data = Z;
		19'b1001000110100011001: color_data = Z;
		19'b1001000110100011010: color_data = Z;
		19'b1001000110100011011: color_data = Z;
		19'b1001000110100011100: color_data = Z;
		19'b1001000110100011101: color_data = Z;
		19'b1001000110100011110: color_data = Z;
		19'b1001000110100011111: color_data = Z;
		19'b1001000110100100000: color_data = Z;
		19'b1001000110100100001: color_data = Z;
		19'b1001000110100100010: color_data = Z;
		19'b1001000110100100011: color_data = Z;
		19'b1001000110100100100: color_data = Z;
		19'b1001000110100100101: color_data = Z;
		19'b1001000110100100110: color_data = Z;
		19'b1001000110100100111: color_data = Z;
		19'b1001000110100101000: color_data = Z;
		19'b1001000110100101001: color_data = Z;
		19'b1001000110100101010: color_data = Z;
		19'b1001000110100101011: color_data = Z;
		19'b1001000110100101100: color_data = Z;
		19'b1001000110100101101: color_data = Z;
		19'b1001000110100101110: color_data = Z;
		19'b1001000110100101111: color_data = Z;
		19'b1001000110100110000: color_data = Z;
		19'b1001000110100110001: color_data = Z;
		19'b1001000110100110010: color_data = Z;
		19'b1001000110100110011: color_data = Z;
		19'b1001000110100110100: color_data = Z;
		19'b1001000110100110101: color_data = Z;
		19'b1001000110100110110: color_data = Z;
		19'b1001000110100110111: color_data = Z;
		19'b1001000110100111000: color_data = Z;
		19'b1001000110100111001: color_data = Z;
		19'b1001000110100111010: color_data = Z;
		19'b1001000110100111011: color_data = Z;
		19'b1001000110100111100: color_data = Z;
		19'b1001000110100111101: color_data = Z;
		19'b1001000110100111110: color_data = Z;
		19'b1001000110100111111: color_data = Z;
		19'b1001000110101000000: color_data = Z;
		19'b1001000110101000001: color_data = Z;
		19'b1001000110101000010: color_data = Z;
		19'b1001000110101000011: color_data = Z;
		19'b1001000110101000100: color_data = Z;
		19'b1001000110101000101: color_data = Z;
		19'b1001000110101000110: color_data = Z;
		19'b1001000110101000111: color_data = Z;
		19'b1001000110101001000: color_data = Z;
		19'b1001000110101001001: color_data = Z;
		19'b1001000110101001010: color_data = Z;
		19'b1001000110101001011: color_data = Z;
		19'b1001000110101001100: color_data = Z;
		19'b1001000110101001101: color_data = Z;
		19'b1001000110101001110: color_data = Z;
		19'b1001000110101001111: color_data = Z;
		19'b1001000110101010000: color_data = Z;
		19'b1001000110101010001: color_data = Z;
		19'b1001000110101010010: color_data = Z;
		19'b1001000110101010011: color_data = Z;
		19'b1001000110101010100: color_data = Z;
		19'b1001000110101010101: color_data = Z;
		19'b1001000110101010110: color_data = Z;
		19'b1001000110101010111: color_data = Z;
		19'b1001000110101011000: color_data = Z;
		19'b1001000110101011001: color_data = Z;
		19'b1001000110101011010: color_data = Z;
		19'b1001000110101011011: color_data = Z;
		19'b1001000110101011100: color_data = Z;
		19'b1001000110101011101: color_data = Z;
		19'b1001000110101011110: color_data = Z;
		19'b1001000110101011111: color_data = Z;
		19'b1001000110101100000: color_data = Z;
		19'b1001000110101100001: color_data = Z;
		19'b1001000110101100010: color_data = Z;
		19'b1001000110101100011: color_data = Z;
		19'b1001000110101100100: color_data = Z;
		19'b1001000110101100101: color_data = Z;
		19'b1001000110101100110: color_data = Z;
		19'b1001000110101100111: color_data = Z;
		19'b1001000110101101000: color_data = Z;
		19'b1001000110101101001: color_data = Z;
		19'b1001000110101101010: color_data = Z;
		19'b1001000110101101011: color_data = Z;
		19'b1001000110101101100: color_data = Z;
		19'b1001000110101101101: color_data = Z;
		19'b1001000110101101110: color_data = Z;
		19'b1001000110101101111: color_data = Z;
		19'b1001000110101110000: color_data = Z;
		19'b1001000110101110001: color_data = Z;
		19'b1001000110101110010: color_data = Z;
		19'b1001000110101110011: color_data = Z;
		19'b1001000110101110100: color_data = Z;
		19'b1001000110101110101: color_data = Z;
		19'b1001000110110000110: color_data = Z;
		19'b1001000110110000111: color_data = Z;
		19'b1001000110110001000: color_data = Z;
		19'b1001000110110101110: color_data = Z;
		19'b1001000110110101111: color_data = Z;
		19'b1001000110110110000: color_data = Z;
		19'b1001000110110110001: color_data = Z;
		19'b1001000110110110010: color_data = Z;
		19'b1001000110110110011: color_data = Z;
		19'b1001000110110110100: color_data = Z;
		19'b1001000110110110101: color_data = Z;
		19'b1001000110110110110: color_data = Z;
		19'b1001000110110111010: color_data = Z;
		19'b1001000110110111011: color_data = Z;
		19'b1001000110111001000: color_data = Z;
		19'b1001000110111001001: color_data = Z;
		19'b1001000110111001010: color_data = Z;
		19'b1001000110111001011: color_data = Z;
		19'b1001000110111001100: color_data = Z;
		19'b1001000110111001101: color_data = Z;
		19'b1001001000011001001: color_data = Z;
		19'b1001001000011010101: color_data = Z;
		19'b1001001000011010110: color_data = Z;
		19'b1001001000011010111: color_data = Z;
		19'b1001001000011011000: color_data = Z;
		19'b1001001000011011001: color_data = Z;
		19'b1001001000011011010: color_data = Z;
		19'b1001001000011011011: color_data = Z;
		19'b1001001000011011100: color_data = Z;
		19'b1001001000011011101: color_data = Z;
		19'b1001001000011011110: color_data = Z;
		19'b1001001000011011111: color_data = Z;
		19'b1001001000011100000: color_data = Z;
		19'b1001001000011100001: color_data = Z;
		19'b1001001000011100010: color_data = Z;
		19'b1001001000011100011: color_data = Z;
		19'b1001001000011100100: color_data = Z;
		19'b1001001000011100101: color_data = Z;
		19'b1001001000011100110: color_data = Z;
		19'b1001001000011100111: color_data = Z;
		19'b1001001000011101010: color_data = Z;
		19'b1001001000011101011: color_data = Z;
		19'b1001001000011101100: color_data = Z;
		19'b1001001000011101101: color_data = Z;
		19'b1001001000011101110: color_data = Z;
		19'b1001001000011101111: color_data = Z;
		19'b1001001000011110000: color_data = Z;
		19'b1001001000011110001: color_data = Z;
		19'b1001001000011110010: color_data = Z;
		19'b1001001000011110011: color_data = Z;
		19'b1001001000100011000: color_data = Z;
		19'b1001001000100011110: color_data = Z;
		19'b1001001000100011111: color_data = Z;
		19'b1001001000100100000: color_data = Z;
		19'b1001001000100100001: color_data = Z;
		19'b1001001000100100010: color_data = Z;
		19'b1001001000100100011: color_data = Z;
		19'b1001001000100100100: color_data = Z;
		19'b1001001000100100101: color_data = Z;
		19'b1001001000100100110: color_data = Z;
		19'b1001001000100100111: color_data = Z;
		19'b1001001000100101000: color_data = Z;
		19'b1001001000100101001: color_data = Z;
		19'b1001001000100101010: color_data = Z;
		19'b1001001000100101011: color_data = Z;
		19'b1001001000100101100: color_data = Z;
		19'b1001001000100101101: color_data = Z;
		19'b1001001000100101110: color_data = Z;
		19'b1001001000100101111: color_data = Z;
		19'b1001001000100110000: color_data = Z;
		19'b1001001000100110001: color_data = Z;
		19'b1001001000100110010: color_data = Z;
		19'b1001001000100110011: color_data = Z;
		19'b1001001000100110100: color_data = Z;
		19'b1001001000100110101: color_data = Z;
		19'b1001001000100110110: color_data = Z;
		19'b1001001000100110111: color_data = Z;
		19'b1001001000100111000: color_data = Z;
		19'b1001001000100111001: color_data = Z;
		19'b1001001000100111010: color_data = Z;
		19'b1001001000100111011: color_data = Z;
		19'b1001001000100111100: color_data = Z;
		19'b1001001000100111101: color_data = Z;
		19'b1001001000100111110: color_data = Z;
		19'b1001001000100111111: color_data = Z;
		19'b1001001000101000000: color_data = Z;
		19'b1001001000101000001: color_data = Z;
		19'b1001001000101000010: color_data = Z;
		19'b1001001000101000011: color_data = Z;
		19'b1001001000101000100: color_data = Z;
		19'b1001001000101000101: color_data = Z;
		19'b1001001000101000110: color_data = Z;
		19'b1001001000101000111: color_data = Z;
		19'b1001001000101001000: color_data = Z;
		19'b1001001000101001001: color_data = Z;
		19'b1001001000101001010: color_data = Z;
		19'b1001001000101001011: color_data = Z;
		19'b1001001000101001100: color_data = Z;
		19'b1001001000101001101: color_data = Z;
		19'b1001001000101001110: color_data = Z;
		19'b1001001000101001111: color_data = Z;
		19'b1001001000101010000: color_data = Z;
		19'b1001001000101010001: color_data = Z;
		19'b1001001000101010010: color_data = Z;
		19'b1001001000101010011: color_data = Z;
		19'b1001001000101010100: color_data = Z;
		19'b1001001000101010101: color_data = Z;
		19'b1001001000101010110: color_data = Z;
		19'b1001001000101010111: color_data = Z;
		19'b1001001000101011000: color_data = Z;
		19'b1001001000101011001: color_data = Z;
		19'b1001001000101011010: color_data = Z;
		19'b1001001000101011011: color_data = Z;
		19'b1001001000101011100: color_data = Z;
		19'b1001001000101011101: color_data = Z;
		19'b1001001000101011110: color_data = Z;
		19'b1001001000101011111: color_data = Z;
		19'b1001001000101100000: color_data = Z;
		19'b1001001000101100001: color_data = Z;
		19'b1001001000101100010: color_data = Z;
		19'b1001001000101100011: color_data = Z;
		19'b1001001000101100100: color_data = Z;
		19'b1001001000101100101: color_data = Z;
		19'b1001001000101100110: color_data = Z;
		19'b1001001000101100111: color_data = Z;
		19'b1001001000101101000: color_data = Z;
		19'b1001001000101101001: color_data = Z;
		19'b1001001000101101010: color_data = Z;
		19'b1001001000101101011: color_data = Z;
		19'b1001001000101101100: color_data = Z;
		19'b1001001000101101101: color_data = Z;
		19'b1001001000101101110: color_data = Z;
		19'b1001001000101101111: color_data = Z;
		19'b1001001000101110000: color_data = Z;
		19'b1001001000101110001: color_data = Z;
		19'b1001001000110000100: color_data = Z;
		19'b1001001000110000101: color_data = Z;
		19'b1001001000110000110: color_data = Z;
		19'b1001001000110000111: color_data = Z;
		19'b1001001000110001000: color_data = Z;
		19'b1001001000110101111: color_data = Z;
		19'b1001001000110110000: color_data = Z;
		19'b1001001000110110001: color_data = Z;
		19'b1001001000110110010: color_data = Z;
		19'b1001001000110110011: color_data = Z;
		19'b1001001000110110100: color_data = Z;
		19'b1001001000110110101: color_data = Z;
		19'b1001001000110110110: color_data = Z;
		19'b1001001000110111011: color_data = Z;
		19'b1001001000111001000: color_data = Z;
		19'b1001001000111001001: color_data = Z;
		19'b1001001000111001010: color_data = Z;
		19'b1001001000111001011: color_data = Z;
		19'b1001001000111001100: color_data = Z;
		19'b1001001000111001101: color_data = Z;
		19'b1001001010011001000: color_data = Z;
		19'b1001001010011010101: color_data = Z;
		19'b1001001010011010110: color_data = Z;
		19'b1001001010011010111: color_data = Z;
		19'b1001001010011011000: color_data = Z;
		19'b1001001010011011001: color_data = Z;
		19'b1001001010011011010: color_data = Z;
		19'b1001001010011011011: color_data = Z;
		19'b1001001010011011100: color_data = Z;
		19'b1001001010011011101: color_data = Z;
		19'b1001001010011011110: color_data = Z;
		19'b1001001010011011111: color_data = Z;
		19'b1001001010011100000: color_data = Z;
		19'b1001001010011100001: color_data = Z;
		19'b1001001010011100010: color_data = Z;
		19'b1001001010011100011: color_data = Z;
		19'b1001001010011100100: color_data = Z;
		19'b1001001010011100101: color_data = Z;
		19'b1001001010011100110: color_data = Z;
		19'b1001001010011101010: color_data = Z;
		19'b1001001010011101011: color_data = Z;
		19'b1001001010011101100: color_data = Z;
		19'b1001001010011101101: color_data = Z;
		19'b1001001010011101110: color_data = Z;
		19'b1001001010011101111: color_data = Z;
		19'b1001001010011110000: color_data = Z;
		19'b1001001010011110001: color_data = Z;
		19'b1001001010011110010: color_data = Z;
		19'b1001001010100011110: color_data = Z;
		19'b1001001010100011111: color_data = Z;
		19'b1001001010100100000: color_data = Z;
		19'b1001001010100100001: color_data = Z;
		19'b1001001010100100010: color_data = Z;
		19'b1001001010100100011: color_data = Z;
		19'b1001001010100100100: color_data = Z;
		19'b1001001010100100101: color_data = Z;
		19'b1001001010100100110: color_data = Z;
		19'b1001001010100100111: color_data = Z;
		19'b1001001010100101000: color_data = Z;
		19'b1001001010100101001: color_data = Z;
		19'b1001001010100101010: color_data = Z;
		19'b1001001010100101011: color_data = Z;
		19'b1001001010100101100: color_data = Z;
		19'b1001001010100101101: color_data = Z;
		19'b1001001010100101110: color_data = Z;
		19'b1001001010100101111: color_data = Z;
		19'b1001001010100110000: color_data = Z;
		19'b1001001010100110001: color_data = Z;
		19'b1001001010100110010: color_data = Z;
		19'b1001001010100110011: color_data = Z;
		19'b1001001010100110100: color_data = Z;
		19'b1001001010100110101: color_data = Z;
		19'b1001001010100110110: color_data = Z;
		19'b1001001010100110111: color_data = Z;
		19'b1001001010100111000: color_data = Z;
		19'b1001001010100111001: color_data = Z;
		19'b1001001010100111010: color_data = Z;
		19'b1001001010100111011: color_data = Z;
		19'b1001001010100111100: color_data = Z;
		19'b1001001010100111101: color_data = Z;
		19'b1001001010100111110: color_data = Z;
		19'b1001001010100111111: color_data = Z;
		19'b1001001010101000000: color_data = Z;
		19'b1001001010101000001: color_data = Z;
		19'b1001001010101000010: color_data = Z;
		19'b1001001010101000011: color_data = Z;
		19'b1001001010101000100: color_data = Z;
		19'b1001001010101000101: color_data = Z;
		19'b1001001010101000110: color_data = Z;
		19'b1001001010101000111: color_data = Z;
		19'b1001001010101001000: color_data = Z;
		19'b1001001010101001001: color_data = Z;
		19'b1001001010101001010: color_data = Z;
		19'b1001001010101001011: color_data = Z;
		19'b1001001010101001100: color_data = Z;
		19'b1001001010101001101: color_data = Z;
		19'b1001001010101001110: color_data = Z;
		19'b1001001010101001111: color_data = Z;
		19'b1001001010101010000: color_data = Z;
		19'b1001001010101010001: color_data = Z;
		19'b1001001010101010010: color_data = Z;
		19'b1001001010101010011: color_data = Z;
		19'b1001001010101010100: color_data = Z;
		19'b1001001010101010101: color_data = Z;
		19'b1001001010101010110: color_data = Z;
		19'b1001001010101010111: color_data = Z;
		19'b1001001010101011000: color_data = Z;
		19'b1001001010101011001: color_data = Z;
		19'b1001001010101011010: color_data = Z;
		19'b1001001010101011011: color_data = Z;
		19'b1001001010101011100: color_data = Z;
		19'b1001001010101011101: color_data = Z;
		19'b1001001010101011110: color_data = Z;
		19'b1001001010101011111: color_data = Z;
		19'b1001001010101100000: color_data = Z;
		19'b1001001010101100001: color_data = Z;
		19'b1001001010101100010: color_data = Z;
		19'b1001001010101100011: color_data = Z;
		19'b1001001010101100100: color_data = Z;
		19'b1001001010101100101: color_data = Z;
		19'b1001001010101100110: color_data = Z;
		19'b1001001010101100111: color_data = Z;
		19'b1001001010101101000: color_data = Z;
		19'b1001001010101101001: color_data = Z;
		19'b1001001010101101010: color_data = Z;
		19'b1001001010101101011: color_data = Z;
		19'b1001001010101101100: color_data = Z;
		19'b1001001010101101101: color_data = Z;
		19'b1001001010101101110: color_data = Z;
		19'b1001001010101101111: color_data = Z;
		19'b1001001010110000010: color_data = Z;
		19'b1001001010110000011: color_data = Z;
		19'b1001001010110000100: color_data = Z;
		19'b1001001010110000101: color_data = Z;
		19'b1001001010110000110: color_data = Z;
		19'b1001001010110000111: color_data = Z;
		19'b1001001010110101111: color_data = Z;
		19'b1001001010110110000: color_data = Z;
		19'b1001001010110110001: color_data = Z;
		19'b1001001010110110010: color_data = Z;
		19'b1001001010110110011: color_data = Z;
		19'b1001001010110110100: color_data = Z;
		19'b1001001010110110101: color_data = Z;
		19'b1001001010110110110: color_data = Z;
		19'b1001001010111001000: color_data = Z;
		19'b1001001010111001001: color_data = Z;
		19'b1001001010111001010: color_data = Z;
		19'b1001001010111001011: color_data = Z;
		19'b1001001010111001100: color_data = Z;
		19'b1001001010111001101: color_data = Z;
		19'b1001001100011000111: color_data = Z;
		19'b1001001100011010101: color_data = Z;
		19'b1001001100011010110: color_data = Z;
		19'b1001001100011010111: color_data = Z;
		19'b1001001100011011000: color_data = Z;
		19'b1001001100011011001: color_data = Z;
		19'b1001001100011011010: color_data = Z;
		19'b1001001100011011011: color_data = Z;
		19'b1001001100011011100: color_data = Z;
		19'b1001001100011011101: color_data = Z;
		19'b1001001100011011110: color_data = Z;
		19'b1001001100011011111: color_data = Z;
		19'b1001001100011100000: color_data = Z;
		19'b1001001100011100001: color_data = Z;
		19'b1001001100011100010: color_data = Z;
		19'b1001001100011100011: color_data = Z;
		19'b1001001100011100100: color_data = Z;
		19'b1001001100011100101: color_data = Z;
		19'b1001001100011100110: color_data = Z;
		19'b1001001100011101010: color_data = Z;
		19'b1001001100011101011: color_data = Z;
		19'b1001001100011101100: color_data = Z;
		19'b1001001100011101101: color_data = Z;
		19'b1001001100011101110: color_data = Z;
		19'b1001001100011101111: color_data = Z;
		19'b1001001100011110000: color_data = Z;
		19'b1001001100011110001: color_data = Z;
		19'b1001001100100100001: color_data = Z;
		19'b1001001100100100010: color_data = Z;
		19'b1001001100100100011: color_data = Z;
		19'b1001001100100100100: color_data = Z;
		19'b1001001100100100101: color_data = Z;
		19'b1001001100100100110: color_data = Z;
		19'b1001001100100100111: color_data = Z;
		19'b1001001100100101000: color_data = Z;
		19'b1001001100100101001: color_data = Z;
		19'b1001001100100101010: color_data = Z;
		19'b1001001100100101011: color_data = Z;
		19'b1001001100100101100: color_data = Z;
		19'b1001001100100101101: color_data = Z;
		19'b1001001100100101110: color_data = Z;
		19'b1001001100100101111: color_data = Z;
		19'b1001001100100110000: color_data = Z;
		19'b1001001100100110001: color_data = Z;
		19'b1001001100100110010: color_data = Z;
		19'b1001001100100110011: color_data = Z;
		19'b1001001100100110100: color_data = Z;
		19'b1001001100100110101: color_data = Z;
		19'b1001001100100110110: color_data = Z;
		19'b1001001100100110111: color_data = Z;
		19'b1001001100100111000: color_data = Z;
		19'b1001001100100111001: color_data = Z;
		19'b1001001100100111010: color_data = Z;
		19'b1001001100100111011: color_data = Z;
		19'b1001001100100111100: color_data = Z;
		19'b1001001100100111101: color_data = Z;
		19'b1001001100100111110: color_data = Z;
		19'b1001001100100111111: color_data = Z;
		19'b1001001100101000000: color_data = Z;
		19'b1001001100101000001: color_data = Z;
		19'b1001001100101000010: color_data = Z;
		19'b1001001100101000011: color_data = Z;
		19'b1001001100101000100: color_data = Z;
		19'b1001001100101000101: color_data = Z;
		19'b1001001100101000110: color_data = Z;
		19'b1001001100101000111: color_data = Z;
		19'b1001001100101001000: color_data = Z;
		19'b1001001100101001001: color_data = Z;
		19'b1001001100101001010: color_data = Z;
		19'b1001001100101001011: color_data = Z;
		19'b1001001100101001100: color_data = Z;
		19'b1001001100101001101: color_data = Z;
		19'b1001001100101001110: color_data = Z;
		19'b1001001100101001111: color_data = Z;
		19'b1001001100101010000: color_data = Z;
		19'b1001001100101010001: color_data = Z;
		19'b1001001100101010010: color_data = Z;
		19'b1001001100101010011: color_data = Z;
		19'b1001001100101010100: color_data = Z;
		19'b1001001100101010101: color_data = Z;
		19'b1001001100101010110: color_data = Z;
		19'b1001001100101010111: color_data = Z;
		19'b1001001100101011000: color_data = Z;
		19'b1001001100101011001: color_data = Z;
		19'b1001001100101011010: color_data = Z;
		19'b1001001100101011011: color_data = Z;
		19'b1001001100101011100: color_data = Z;
		19'b1001001100101011101: color_data = Z;
		19'b1001001100101011110: color_data = Z;
		19'b1001001100101011111: color_data = Z;
		19'b1001001100101100000: color_data = Z;
		19'b1001001100101100001: color_data = Z;
		19'b1001001100101100010: color_data = Z;
		19'b1001001100101100011: color_data = Z;
		19'b1001001100101100100: color_data = Z;
		19'b1001001100101100101: color_data = Z;
		19'b1001001100101100110: color_data = Z;
		19'b1001001100101100111: color_data = Z;
		19'b1001001100101101000: color_data = Z;
		19'b1001001100110000001: color_data = Z;
		19'b1001001100110000010: color_data = Z;
		19'b1001001100110000011: color_data = Z;
		19'b1001001100110000100: color_data = Z;
		19'b1001001100110110000: color_data = Z;
		19'b1001001100110110001: color_data = Z;
		19'b1001001100110110010: color_data = Z;
		19'b1001001100110110011: color_data = Z;
		19'b1001001100110110100: color_data = Z;
		19'b1001001100110110101: color_data = Z;
		19'b1001001100110110110: color_data = Z;
		19'b1001001100111001001: color_data = Z;
		19'b1001001100111001010: color_data = Z;
		19'b1001001100111001011: color_data = Z;
		19'b1001001100111001100: color_data = Z;
		19'b1001001100111001101: color_data = Z;
		19'b1001001110011000111: color_data = Z;
		19'b1001001110011010101: color_data = Z;
		19'b1001001110011010110: color_data = Z;
		19'b1001001110011010111: color_data = Z;
		19'b1001001110011011000: color_data = Z;
		19'b1001001110011011001: color_data = Z;
		19'b1001001110011011010: color_data = Z;
		19'b1001001110011011011: color_data = Z;
		19'b1001001110011011100: color_data = Z;
		19'b1001001110011011101: color_data = Z;
		19'b1001001110011011110: color_data = Z;
		19'b1001001110011011111: color_data = Z;
		19'b1001001110011100000: color_data = Z;
		19'b1001001110011100001: color_data = Z;
		19'b1001001110011100010: color_data = Z;
		19'b1001001110011100011: color_data = Z;
		19'b1001001110011100100: color_data = Z;
		19'b1001001110011100101: color_data = Z;
		19'b1001001110011101001: color_data = Z;
		19'b1001001110011101010: color_data = Z;
		19'b1001001110011101011: color_data = Z;
		19'b1001001110011101100: color_data = Z;
		19'b1001001110011101101: color_data = Z;
		19'b1001001110011101110: color_data = Z;
		19'b1001001110011101111: color_data = Z;
		19'b1001001110100100010: color_data = Z;
		19'b1001001110100100011: color_data = Z;
		19'b1001001110100100100: color_data = Z;
		19'b1001001110100100101: color_data = Z;
		19'b1001001110100100110: color_data = Z;
		19'b1001001110100100111: color_data = Z;
		19'b1001001110100101000: color_data = Z;
		19'b1001001110100101001: color_data = Z;
		19'b1001001110100101010: color_data = Z;
		19'b1001001110100101011: color_data = Z;
		19'b1001001110100101100: color_data = Z;
		19'b1001001110100101101: color_data = Z;
		19'b1001001110100101110: color_data = Z;
		19'b1001001110100101111: color_data = Z;
		19'b1001001110100110000: color_data = Z;
		19'b1001001110100110001: color_data = Z;
		19'b1001001110100110010: color_data = Z;
		19'b1001001110100110011: color_data = Z;
		19'b1001001110100110100: color_data = Z;
		19'b1001001110100110101: color_data = Z;
		19'b1001001110100110110: color_data = Z;
		19'b1001001110100110111: color_data = Z;
		19'b1001001110100111000: color_data = Z;
		19'b1001001110100111001: color_data = Z;
		19'b1001001110100111010: color_data = Z;
		19'b1001001110100111011: color_data = Z;
		19'b1001001110100111100: color_data = Z;
		19'b1001001110100111101: color_data = Z;
		19'b1001001110100111110: color_data = Z;
		19'b1001001110100111111: color_data = Z;
		19'b1001001110101000000: color_data = Z;
		19'b1001001110101000001: color_data = Z;
		19'b1001001110101000010: color_data = Z;
		19'b1001001110101000011: color_data = Z;
		19'b1001001110101000100: color_data = Z;
		19'b1001001110101000101: color_data = Z;
		19'b1001001110101000110: color_data = Z;
		19'b1001001110101000111: color_data = Z;
		19'b1001001110101001000: color_data = Z;
		19'b1001001110101001001: color_data = Z;
		19'b1001001110101001010: color_data = Z;
		19'b1001001110101001011: color_data = Z;
		19'b1001001110101001100: color_data = Z;
		19'b1001001110101001101: color_data = Z;
		19'b1001001110101001110: color_data = Z;
		19'b1001001110101001111: color_data = Z;
		19'b1001001110101010000: color_data = Z;
		19'b1001001110101010001: color_data = Z;
		19'b1001001110101010010: color_data = Z;
		19'b1001001110101010011: color_data = Z;
		19'b1001001110101010100: color_data = Z;
		19'b1001001110101010101: color_data = Z;
		19'b1001001110101010110: color_data = Z;
		19'b1001001110101010111: color_data = Z;
		19'b1001001110101011000: color_data = Z;
		19'b1001001110101011001: color_data = Z;
		19'b1001001110101011010: color_data = Z;
		19'b1001001110101011011: color_data = Z;
		19'b1001001110101011100: color_data = Z;
		19'b1001001110101011101: color_data = Z;
		19'b1001001110101011110: color_data = Z;
		19'b1001001110101011111: color_data = Z;
		19'b1001001110101100000: color_data = Z;
		19'b1001001110101100001: color_data = Z;
		19'b1001001110101100010: color_data = Z;
		19'b1001001110101100011: color_data = Z;
		19'b1001001110101100100: color_data = Z;
		19'b1001001110110110000: color_data = Z;
		19'b1001001110110110001: color_data = Z;
		19'b1001001110110110010: color_data = Z;
		19'b1001001110110110011: color_data = Z;
		19'b1001001110110110100: color_data = Z;
		19'b1001001110110110101: color_data = Z;
		19'b1001001110110110110: color_data = Z;
		19'b1001001110111001001: color_data = Z;
		19'b1001001110111001010: color_data = Z;
		19'b1001001110111001011: color_data = Z;
		19'b1001001110111001100: color_data = Z;
		19'b1001001110111001101: color_data = Z;
		19'b1001010000011000111: color_data = Z;
		19'b1001010000011010100: color_data = Z;
		19'b1001010000011010101: color_data = Z;
		19'b1001010000011010110: color_data = Z;
		19'b1001010000011010111: color_data = Z;
		19'b1001010000011011000: color_data = Z;
		19'b1001010000011011001: color_data = Z;
		19'b1001010000011011010: color_data = Z;
		19'b1001010000011011011: color_data = Z;
		19'b1001010000011011100: color_data = Z;
		19'b1001010000011011101: color_data = Z;
		19'b1001010000011011110: color_data = Z;
		19'b1001010000011011111: color_data = Z;
		19'b1001010000011100000: color_data = Z;
		19'b1001010000011100001: color_data = Z;
		19'b1001010000011100010: color_data = Z;
		19'b1001010000011100011: color_data = Z;
		19'b1001010000011100100: color_data = Z;
		19'b1001010000011100101: color_data = Z;
		19'b1001010000011101001: color_data = Z;
		19'b1001010000011101010: color_data = Z;
		19'b1001010000011101011: color_data = Z;
		19'b1001010000011101100: color_data = Z;
		19'b1001010000011101101: color_data = Z;
		19'b1001010000100100011: color_data = Z;
		19'b1001010000100100100: color_data = Z;
		19'b1001010000100100101: color_data = Z;
		19'b1001010000100100110: color_data = Z;
		19'b1001010000100100111: color_data = Z;
		19'b1001010000100101000: color_data = Z;
		19'b1001010000100101001: color_data = Z;
		19'b1001010000100101010: color_data = Z;
		19'b1001010000100101011: color_data = Z;
		19'b1001010000100101100: color_data = Z;
		19'b1001010000100101101: color_data = Z;
		19'b1001010000100101110: color_data = Z;
		19'b1001010000100101111: color_data = Z;
		19'b1001010000100110000: color_data = Z;
		19'b1001010000100110001: color_data = Z;
		19'b1001010000100110010: color_data = Z;
		19'b1001010000100110011: color_data = Z;
		19'b1001010000100110100: color_data = Z;
		19'b1001010000100110101: color_data = Z;
		19'b1001010000100110110: color_data = Z;
		19'b1001010000100110111: color_data = Z;
		19'b1001010000100111000: color_data = Z;
		19'b1001010000100111001: color_data = Z;
		19'b1001010000100111010: color_data = Z;
		19'b1001010000100111011: color_data = Z;
		19'b1001010000100111100: color_data = Z;
		19'b1001010000100111101: color_data = Z;
		19'b1001010000100111110: color_data = Z;
		19'b1001010000100111111: color_data = Z;
		19'b1001010000101000000: color_data = Z;
		19'b1001010000101000001: color_data = Z;
		19'b1001010000101000010: color_data = Z;
		19'b1001010000101000011: color_data = Z;
		19'b1001010000101000100: color_data = Z;
		19'b1001010000101000101: color_data = Z;
		19'b1001010000101000110: color_data = Z;
		19'b1001010000101000111: color_data = Z;
		19'b1001010000101001000: color_data = Z;
		19'b1001010000101001001: color_data = Z;
		19'b1001010000101001010: color_data = Z;
		19'b1001010000101001011: color_data = Z;
		19'b1001010000101001100: color_data = Z;
		19'b1001010000101001101: color_data = Z;
		19'b1001010000101001110: color_data = Z;
		19'b1001010000101001111: color_data = Z;
		19'b1001010000101010000: color_data = Z;
		19'b1001010000101010001: color_data = Z;
		19'b1001010000101010010: color_data = Z;
		19'b1001010000101010011: color_data = Z;
		19'b1001010000101010100: color_data = Z;
		19'b1001010000101010101: color_data = Z;
		19'b1001010000101010110: color_data = Z;
		19'b1001010000101010111: color_data = Z;
		19'b1001010000101011000: color_data = Z;
		19'b1001010000101011001: color_data = Z;
		19'b1001010000101011010: color_data = Z;
		19'b1001010000101011011: color_data = Z;
		19'b1001010000101011100: color_data = Z;
		19'b1001010000110110000: color_data = Z;
		19'b1001010000110110001: color_data = Z;
		19'b1001010000110110010: color_data = Z;
		19'b1001010000110110011: color_data = Z;
		19'b1001010000110110100: color_data = Z;
		19'b1001010000110110101: color_data = Z;
		19'b1001010000110110110: color_data = Z;
		19'b1001010000110110111: color_data = Z;
		19'b1001010000111001001: color_data = Z;
		19'b1001010000111001010: color_data = Z;
		19'b1001010000111001011: color_data = Z;
		19'b1001010000111001100: color_data = Z;
		19'b1001010000111001101: color_data = Z;
		19'b1001010010011010100: color_data = Z;
		19'b1001010010011010101: color_data = Z;
		19'b1001010010011010110: color_data = Z;
		19'b1001010010011010111: color_data = Z;
		19'b1001010010011011000: color_data = Z;
		19'b1001010010011011001: color_data = Z;
		19'b1001010010011011010: color_data = Z;
		19'b1001010010011011011: color_data = Z;
		19'b1001010010011011100: color_data = Z;
		19'b1001010010011011101: color_data = Z;
		19'b1001010010011011110: color_data = Z;
		19'b1001010010011011111: color_data = Z;
		19'b1001010010011100000: color_data = Z;
		19'b1001010010011100001: color_data = Z;
		19'b1001010010011100010: color_data = Z;
		19'b1001010010011100011: color_data = Z;
		19'b1001010010011100100: color_data = Z;
		19'b1001010010011101001: color_data = Z;
		19'b1001010010011101010: color_data = Z;
		19'b1001010010011101011: color_data = Z;
		19'b1001010010011101100: color_data = Z;
		19'b1001010010100100101: color_data = Z;
		19'b1001010010100100110: color_data = Z;
		19'b1001010010100100111: color_data = Z;
		19'b1001010010100101000: color_data = Z;
		19'b1001010010100101001: color_data = Z;
		19'b1001010010100101010: color_data = Z;
		19'b1001010010100101011: color_data = Z;
		19'b1001010010100101100: color_data = Z;
		19'b1001010010100101101: color_data = Z;
		19'b1001010010100101110: color_data = Z;
		19'b1001010010100101111: color_data = Z;
		19'b1001010010100110000: color_data = Z;
		19'b1001010010100110001: color_data = Z;
		19'b1001010010100110010: color_data = Z;
		19'b1001010010100110011: color_data = Z;
		19'b1001010010100110100: color_data = Z;
		19'b1001010010100110101: color_data = Z;
		19'b1001010010100110110: color_data = Z;
		19'b1001010010100110111: color_data = Z;
		19'b1001010010100111000: color_data = Z;
		19'b1001010010100111001: color_data = Z;
		19'b1001010010100111010: color_data = Z;
		19'b1001010010100111011: color_data = Z;
		19'b1001010010100111100: color_data = Z;
		19'b1001010010100111101: color_data = Z;
		19'b1001010010100111110: color_data = Z;
		19'b1001010010100111111: color_data = Z;
		19'b1001010010101000000: color_data = Z;
		19'b1001010010101000001: color_data = Z;
		19'b1001010010101000010: color_data = Z;
		19'b1001010010101000011: color_data = Z;
		19'b1001010010101000100: color_data = Z;
		19'b1001010010101000101: color_data = Z;
		19'b1001010010101000110: color_data = Z;
		19'b1001010010101000111: color_data = Z;
		19'b1001010010101001000: color_data = Z;
		19'b1001010010101001001: color_data = Z;
		19'b1001010010101001010: color_data = Z;
		19'b1001010010101001011: color_data = Z;
		19'b1001010010101001100: color_data = Z;
		19'b1001010010101001101: color_data = Z;
		19'b1001010010101001110: color_data = Z;
		19'b1001010010101001111: color_data = Z;
		19'b1001010010101010000: color_data = Z;
		19'b1001010010101010001: color_data = Z;
		19'b1001010010101010010: color_data = Z;
		19'b1001010010101010011: color_data = Z;
		19'b1001010010101010100: color_data = Z;
		19'b1001010010101010101: color_data = Z;
		19'b1001010010101010110: color_data = Z;
		19'b1001010010101010111: color_data = Z;
		19'b1001010010101011000: color_data = Z;
		19'b1001010010110000100: color_data = Z;
		19'b1001010010110000101: color_data = Z;
		19'b1001010010110110001: color_data = Z;
		19'b1001010010110110010: color_data = Z;
		19'b1001010010110110011: color_data = Z;
		19'b1001010010110110100: color_data = Z;
		19'b1001010010110110101: color_data = Z;
		19'b1001010010110110110: color_data = Z;
		19'b1001010010110110111: color_data = Z;
		19'b1001010010111001001: color_data = Z;
		19'b1001010010111001010: color_data = Z;
		19'b1001010010111001011: color_data = Z;
		19'b1001010010111001100: color_data = Z;
		19'b1001010010111001101: color_data = Z;
		19'b1001010100011010100: color_data = Z;
		19'b1001010100011010101: color_data = Z;
		19'b1001010100011010110: color_data = Z;
		19'b1001010100011010111: color_data = Z;
		19'b1001010100011011000: color_data = Z;
		19'b1001010100011011001: color_data = Z;
		19'b1001010100011011010: color_data = Z;
		19'b1001010100011011011: color_data = Z;
		19'b1001010100011011100: color_data = Z;
		19'b1001010100011011101: color_data = Z;
		19'b1001010100011011110: color_data = Z;
		19'b1001010100011011111: color_data = Z;
		19'b1001010100011100000: color_data = Z;
		19'b1001010100011100001: color_data = Z;
		19'b1001010100011100010: color_data = Z;
		19'b1001010100011100011: color_data = Z;
		19'b1001010100011100100: color_data = Z;
		19'b1001010100011101001: color_data = Z;
		19'b1001010100011101010: color_data = Z;
		19'b1001010100011101011: color_data = Z;
		19'b1001010100100101010: color_data = Z;
		19'b1001010100100101011: color_data = Z;
		19'b1001010100100101100: color_data = Z;
		19'b1001010100100101110: color_data = Z;
		19'b1001010100100101111: color_data = Z;
		19'b1001010100100110000: color_data = Z;
		19'b1001010100100110001: color_data = Z;
		19'b1001010100100110010: color_data = Z;
		19'b1001010100100110011: color_data = Z;
		19'b1001010100100110100: color_data = Z;
		19'b1001010100100110101: color_data = Z;
		19'b1001010100100110110: color_data = Z;
		19'b1001010100100110111: color_data = Z;
		19'b1001010100100111000: color_data = Z;
		19'b1001010100100111001: color_data = Z;
		19'b1001010100100111010: color_data = Z;
		19'b1001010100100111011: color_data = Z;
		19'b1001010100100111100: color_data = Z;
		19'b1001010100100111101: color_data = Z;
		19'b1001010100100111110: color_data = Z;
		19'b1001010100100111111: color_data = Z;
		19'b1001010100101000000: color_data = Z;
		19'b1001010100101000001: color_data = Z;
		19'b1001010100101000010: color_data = Z;
		19'b1001010100101000011: color_data = Z;
		19'b1001010100101000100: color_data = Z;
		19'b1001010100101000101: color_data = Z;
		19'b1001010100101000110: color_data = Z;
		19'b1001010100101000111: color_data = Z;
		19'b1001010100101001000: color_data = Z;
		19'b1001010100101001001: color_data = Z;
		19'b1001010100101001010: color_data = Z;
		19'b1001010100101001011: color_data = Z;
		19'b1001010100101001100: color_data = Z;
		19'b1001010100101001101: color_data = Z;
		19'b1001010100101001110: color_data = Z;
		19'b1001010100101001111: color_data = Z;
		19'b1001010100101010000: color_data = Z;
		19'b1001010100101010001: color_data = Z;
		19'b1001010100101010010: color_data = Z;
		19'b1001010100101111111: color_data = Z;
		19'b1001010100110000000: color_data = Z;
		19'b1001010100110110001: color_data = Z;
		19'b1001010100110110010: color_data = Z;
		19'b1001010100110110011: color_data = Z;
		19'b1001010100110110101: color_data = Z;
		19'b1001010100110110110: color_data = Z;
		19'b1001010100110110111: color_data = Z;
		19'b1001010100111001010: color_data = Z;
		19'b1001010100111001011: color_data = Z;
		19'b1001010100111001100: color_data = Z;
		19'b1001010110011001000: color_data = Z;
		19'b1001010110011010011: color_data = Z;
		19'b1001010110011010100: color_data = Z;
		19'b1001010110011010101: color_data = Z;
		19'b1001010110011010110: color_data = Z;
		19'b1001010110011010111: color_data = Z;
		19'b1001010110011011000: color_data = Z;
		19'b1001010110011011001: color_data = Z;
		19'b1001010110011011010: color_data = Z;
		19'b1001010110011011011: color_data = Z;
		19'b1001010110011011100: color_data = Z;
		19'b1001010110011011101: color_data = Z;
		19'b1001010110011011110: color_data = Z;
		19'b1001010110011011111: color_data = Z;
		19'b1001010110011100000: color_data = Z;
		19'b1001010110011100001: color_data = Z;
		19'b1001010110011100010: color_data = Z;
		19'b1001010110011100011: color_data = Z;
		19'b1001010110011100100: color_data = Z;
		19'b1001010110011100101: color_data = Z;
		19'b1001010110011100111: color_data = Z;
		19'b1001010110011101000: color_data = Z;
		19'b1001010110011101001: color_data = Z;
		19'b1001010110011101010: color_data = Z;
		19'b1001010110100110001: color_data = Z;
		19'b1001010110100110010: color_data = Z;
		19'b1001010110100110011: color_data = Z;
		19'b1001010110100110100: color_data = Z;
		19'b1001010110100110101: color_data = Z;
		19'b1001010110100110110: color_data = Z;
		19'b1001010110100110111: color_data = Z;
		19'b1001010110100111000: color_data = Z;
		19'b1001010110100111001: color_data = Z;
		19'b1001010110100111010: color_data = Z;
		19'b1001010110100111011: color_data = Z;
		19'b1001010110100111100: color_data = Z;
		19'b1001010110100111101: color_data = Z;
		19'b1001010110100111110: color_data = Z;
		19'b1001010110100111111: color_data = Z;
		19'b1001010110101000000: color_data = Z;
		19'b1001010110101000001: color_data = Z;
		19'b1001010110101000010: color_data = Z;
		19'b1001010110101000011: color_data = Z;
		19'b1001010110101000100: color_data = Z;
		19'b1001010110101000101: color_data = Z;
		19'b1001010110101000110: color_data = Z;
		19'b1001010110101000111: color_data = Z;
		19'b1001010110101001000: color_data = Z;
		19'b1001010110101001001: color_data = Z;
		19'b1001010110101001010: color_data = Z;
		19'b1001010110101001011: color_data = Z;
		19'b1001010110101001100: color_data = Z;
		19'b1001010110101001101: color_data = Z;
		19'b1001010110101111101: color_data = Z;
		19'b1001010110101111110: color_data = Z;
		19'b1001010110101111111: color_data = Z;
		19'b1001010110110000000: color_data = Z;
		19'b1001010110110000001: color_data = Z;
		19'b1001010110110110001: color_data = Z;
		19'b1001010110110110010: color_data = Z;
		19'b1001010110110110011: color_data = Z;
		19'b1001010110110110101: color_data = Z;
		19'b1001010110110110110: color_data = Z;
		19'b1001010110110110111: color_data = Z;
		19'b1001010110111001010: color_data = Z;
		19'b1001010110111001011: color_data = Z;
		19'b1001010110111001100: color_data = Z;
		19'b1001011000011001000: color_data = Z;
		19'b1001011000011001001: color_data = Z;
		19'b1001011000011010011: color_data = Z;
		19'b1001011000011010100: color_data = Z;
		19'b1001011000011010101: color_data = Z;
		19'b1001011000011010110: color_data = Z;
		19'b1001011000011010111: color_data = Z;
		19'b1001011000011011000: color_data = Z;
		19'b1001011000011011001: color_data = Z;
		19'b1001011000011011010: color_data = Z;
		19'b1001011000011011011: color_data = Z;
		19'b1001011000011011100: color_data = Z;
		19'b1001011000011011101: color_data = Z;
		19'b1001011000011011110: color_data = Z;
		19'b1001011000011011111: color_data = Z;
		19'b1001011000011100000: color_data = Z;
		19'b1001011000011100001: color_data = Z;
		19'b1001011000011100010: color_data = Z;
		19'b1001011000011100011: color_data = Z;
		19'b1001011000011100100: color_data = Z;
		19'b1001011000011100101: color_data = Z;
		19'b1001011000011100110: color_data = Z;
		19'b1001011000011100111: color_data = Z;
		19'b1001011000011101000: color_data = Z;
		19'b1001011000011101001: color_data = Z;
		19'b1001011000100000110: color_data = Z;
		19'b1001011000100110101: color_data = Z;
		19'b1001011000100110110: color_data = Z;
		19'b1001011000100110111: color_data = Z;
		19'b1001011000100111000: color_data = Z;
		19'b1001011000100111001: color_data = Z;
		19'b1001011000100111010: color_data = Z;
		19'b1001011000100111011: color_data = Z;
		19'b1001011000100111100: color_data = Z;
		19'b1001011000100111101: color_data = Z;
		19'b1001011000100111110: color_data = Z;
		19'b1001011000100111111: color_data = Z;
		19'b1001011000101000000: color_data = Z;
		19'b1001011000101000001: color_data = Z;
		19'b1001011000101000010: color_data = Z;
		19'b1001011000101000011: color_data = Z;
		19'b1001011000101000100: color_data = Z;
		19'b1001011000101000101: color_data = Z;
		19'b1001011000101000110: color_data = Z;
		19'b1001011000101000111: color_data = Z;
		19'b1001011000101001000: color_data = Z;
		19'b1001011000101001001: color_data = Z;
		19'b1001011000101110010: color_data = Z;
		19'b1001011000101110011: color_data = Z;
		19'b1001011000101111101: color_data = Z;
		19'b1001011000101111110: color_data = Z;
		19'b1001011000101111111: color_data = Z;
		19'b1001011000110000000: color_data = Z;
		19'b1001011000110000101: color_data = Z;
		19'b1001011000110110001: color_data = Z;
		19'b1001011000110110010: color_data = Z;
		19'b1001011000110110011: color_data = Z;
		19'b1001011000110110110: color_data = Z;
		19'b1001011000110110111: color_data = Z;
		19'b1001011000111001010: color_data = Z;
		19'b1001011000111001011: color_data = Z;
		19'b1001011010011001001: color_data = Z;
		19'b1001011010011010011: color_data = Z;
		19'b1001011010011010100: color_data = Z;
		19'b1001011010011010101: color_data = Z;
		19'b1001011010011010110: color_data = Z;
		19'b1001011010011010111: color_data = Z;
		19'b1001011010011011000: color_data = Z;
		19'b1001011010011011001: color_data = Z;
		19'b1001011010011011010: color_data = Z;
		19'b1001011010011011011: color_data = Z;
		19'b1001011010011011100: color_data = Z;
		19'b1001011010011011101: color_data = Z;
		19'b1001011010011011110: color_data = Z;
		19'b1001011010011011111: color_data = Z;
		19'b1001011010011100000: color_data = Z;
		19'b1001011010011100001: color_data = Z;
		19'b1001011010011100010: color_data = Z;
		19'b1001011010011100011: color_data = Z;
		19'b1001011010011100100: color_data = Z;
		19'b1001011010011100101: color_data = Z;
		19'b1001011010011100110: color_data = Z;
		19'b1001011010011100111: color_data = Z;
		19'b1001011010011101000: color_data = Z;
		19'b1001011010011101001: color_data = Z;
		19'b1001011010100000110: color_data = Z;
		19'b1001011010100000111: color_data = Z;
		19'b1001011010100001000: color_data = Z;
		19'b1001011010100001001: color_data = Z;
		19'b1001011010100001010: color_data = Z;
		19'b1001011010100001011: color_data = Z;
		19'b1001011010100001100: color_data = Z;
		19'b1001011010100110111: color_data = Z;
		19'b1001011010100111000: color_data = Z;
		19'b1001011010100111001: color_data = Z;
		19'b1001011010100111010: color_data = Z;
		19'b1001011010100111011: color_data = Z;
		19'b1001011010100111100: color_data = Z;
		19'b1001011010100111101: color_data = Z;
		19'b1001011010100111110: color_data = Z;
		19'b1001011010100111111: color_data = Z;
		19'b1001011010101000000: color_data = Z;
		19'b1001011010101000001: color_data = Z;
		19'b1001011010101000010: color_data = Z;
		19'b1001011010101000011: color_data = Z;
		19'b1001011010101000100: color_data = Z;
		19'b1001011010101000101: color_data = Z;
		19'b1001011010101000110: color_data = Z;
		19'b1001011010101000111: color_data = Z;
		19'b1001011010101110010: color_data = Z;
		19'b1001011010101111101: color_data = Z;
		19'b1001011010101111110: color_data = Z;
		19'b1001011010101111111: color_data = Z;
		19'b1001011010110000011: color_data = Z;
		19'b1001011010110000100: color_data = Z;
		19'b1001011010110000101: color_data = Z;
		19'b1001011010110000110: color_data = Z;
		19'b1001011010110110001: color_data = Z;
		19'b1001011010110110010: color_data = Z;
		19'b1001011010110110011: color_data = Z;
		19'b1001011010110110110: color_data = Z;
		19'b1001011010110110111: color_data = Z;
		19'b1001011010111001010: color_data = Z;
		19'b1001011010111001011: color_data = Z;
		19'b1001011100011001001: color_data = Z;
		19'b1001011100011001010: color_data = Z;
		19'b1001011100011010011: color_data = Z;
		19'b1001011100011010100: color_data = Z;
		19'b1001011100011010101: color_data = Z;
		19'b1001011100011010110: color_data = Z;
		19'b1001011100011010111: color_data = Z;
		19'b1001011100011011000: color_data = Z;
		19'b1001011100011011001: color_data = Z;
		19'b1001011100011011010: color_data = Z;
		19'b1001011100011011011: color_data = Z;
		19'b1001011100011011100: color_data = Z;
		19'b1001011100011011101: color_data = Z;
		19'b1001011100011011110: color_data = Z;
		19'b1001011100011011111: color_data = Z;
		19'b1001011100011100000: color_data = Z;
		19'b1001011100011100001: color_data = Z;
		19'b1001011100011100010: color_data = Z;
		19'b1001011100011100011: color_data = Z;
		19'b1001011100011100100: color_data = Z;
		19'b1001011100011100101: color_data = Z;
		19'b1001011100011100110: color_data = Z;
		19'b1001011100011100111: color_data = Z;
		19'b1001011100011101000: color_data = Z;
		19'b1001011100011101001: color_data = Z;
		19'b1001011100011101010: color_data = Z;
		19'b1001011100100000110: color_data = Z;
		19'b1001011100100000111: color_data = Z;
		19'b1001011100100001000: color_data = Z;
		19'b1001011100100001001: color_data = Z;
		19'b1001011100100001010: color_data = Z;
		19'b1001011100100001011: color_data = Z;
		19'b1001011100100001100: color_data = Z;
		19'b1001011100100001101: color_data = Z;
		19'b1001011100100001110: color_data = Z;
		19'b1001011100100111011: color_data = Z;
		19'b1001011100100111100: color_data = Z;
		19'b1001011100100111101: color_data = Z;
		19'b1001011100100111110: color_data = Z;
		19'b1001011100100111111: color_data = Z;
		19'b1001011100101000000: color_data = Z;
		19'b1001011100101000001: color_data = Z;
		19'b1001011100101000010: color_data = Z;
		19'b1001011100101011100: color_data = Z;
		19'b1001011100101011101: color_data = Z;
		19'b1001011100101100100: color_data = Z;
		19'b1001011100101111101: color_data = Z;
		19'b1001011100101111110: color_data = Z;
		19'b1001011100101111111: color_data = Z;
		19'b1001011100110000000: color_data = Z;
		19'b1001011100110000001: color_data = Z;
		19'b1001011100110000010: color_data = Z;
		19'b1001011100110000011: color_data = Z;
		19'b1001011100110000100: color_data = Z;
		19'b1001011100110000101: color_data = Z;
		19'b1001011100110000110: color_data = Z;
		19'b1001011100110110000: color_data = Z;
		19'b1001011100110110001: color_data = Z;
		19'b1001011100110110010: color_data = Z;
		19'b1001011100110110011: color_data = Z;
		19'b1001011100110110110: color_data = Z;
		19'b1001011100110110111: color_data = Z;
		19'b1001011100111001010: color_data = Z;
		19'b1001011110011001010: color_data = Z;
		19'b1001011110011010011: color_data = Z;
		19'b1001011110011010100: color_data = Z;
		19'b1001011110011010101: color_data = Z;
		19'b1001011110011010110: color_data = Z;
		19'b1001011110011010111: color_data = Z;
		19'b1001011110011011000: color_data = Z;
		19'b1001011110011011001: color_data = Z;
		19'b1001011110011011010: color_data = Z;
		19'b1001011110011011011: color_data = Z;
		19'b1001011110011011100: color_data = Z;
		19'b1001011110011011101: color_data = Z;
		19'b1001011110011011110: color_data = Z;
		19'b1001011110011011111: color_data = Z;
		19'b1001011110011100000: color_data = Z;
		19'b1001011110011100001: color_data = Z;
		19'b1001011110011100010: color_data = Z;
		19'b1001011110011100011: color_data = Z;
		19'b1001011110011100100: color_data = Z;
		19'b1001011110011100101: color_data = Z;
		19'b1001011110011100110: color_data = Z;
		19'b1001011110011100111: color_data = Z;
		19'b1001011110011101000: color_data = Z;
		19'b1001011110011101001: color_data = Z;
		19'b1001011110011101010: color_data = Z;
		19'b1001011110100000110: color_data = Z;
		19'b1001011110100000111: color_data = Z;
		19'b1001011110100001000: color_data = Z;
		19'b1001011110100001001: color_data = Z;
		19'b1001011110100001010: color_data = Z;
		19'b1001011110100001011: color_data = Z;
		19'b1001011110100001100: color_data = Z;
		19'b1001011110100001101: color_data = Z;
		19'b1001011110100001110: color_data = Z;
		19'b1001011110100001111: color_data = Z;
		19'b1001011110100010000: color_data = Z;
		19'b1001011110101011011: color_data = Z;
		19'b1001011110101011100: color_data = Z;
		19'b1001011110101011101: color_data = Z;
		19'b1001011110101011110: color_data = Z;
		19'b1001011110101100011: color_data = Z;
		19'b1001011110101100100: color_data = Z;
		19'b1001011110101100101: color_data = Z;
		19'b1001011110101111101: color_data = Z;
		19'b1001011110101111110: color_data = Z;
		19'b1001011110101111111: color_data = Z;
		19'b1001011110110000000: color_data = Z;
		19'b1001011110110000001: color_data = Z;
		19'b1001011110110000010: color_data = Z;
		19'b1001011110110000011: color_data = Z;
		19'b1001011110110000100: color_data = Z;
		19'b1001011110110000101: color_data = Z;
		19'b1001011110110110000: color_data = Z;
		19'b1001011110110110001: color_data = Z;
		19'b1001011110110110010: color_data = Z;
		19'b1001011110110110110: color_data = Z;
		19'b1001011110110110111: color_data = Z;
		19'b1001100000011001010: color_data = Z;
		19'b1001100000011001011: color_data = Z;
		19'b1001100000011010100: color_data = Z;
		19'b1001100000011010101: color_data = Z;
		19'b1001100000011010110: color_data = Z;
		19'b1001100000011010111: color_data = Z;
		19'b1001100000011011000: color_data = Z;
		19'b1001100000011011001: color_data = Z;
		19'b1001100000011011010: color_data = Z;
		19'b1001100000011011011: color_data = Z;
		19'b1001100000011011100: color_data = Z;
		19'b1001100000011011101: color_data = Z;
		19'b1001100000011011110: color_data = Z;
		19'b1001100000011011111: color_data = Z;
		19'b1001100000011100000: color_data = Z;
		19'b1001100000011100001: color_data = Z;
		19'b1001100000011100010: color_data = Z;
		19'b1001100000011100011: color_data = Z;
		19'b1001100000011100100: color_data = Z;
		19'b1001100000011100101: color_data = Z;
		19'b1001100000011100110: color_data = Z;
		19'b1001100000011100111: color_data = Z;
		19'b1001100000011101000: color_data = Z;
		19'b1001100000011101001: color_data = Z;
		19'b1001100000011101010: color_data = Z;
		19'b1001100000100000111: color_data = Z;
		19'b1001100000100001000: color_data = Z;
		19'b1001100000100001001: color_data = Z;
		19'b1001100000100001010: color_data = Z;
		19'b1001100000100001011: color_data = Z;
		19'b1001100000100001100: color_data = Z;
		19'b1001100000100001101: color_data = Z;
		19'b1001100000100001110: color_data = Z;
		19'b1001100000100001111: color_data = Z;
		19'b1001100000100010000: color_data = Z;
		19'b1001100000100010001: color_data = Z;
		19'b1001100000100010010: color_data = Z;
		19'b1001100000100010011: color_data = Z;
		19'b1001100000100010100: color_data = Z;
		19'b1001100000101011101: color_data = Z;
		19'b1001100000101011110: color_data = Z;
		19'b1001100000101100010: color_data = Z;
		19'b1001100000101100011: color_data = Z;
		19'b1001100000101100100: color_data = Z;
		19'b1001100000101100101: color_data = Z;
		19'b1001100000101101011: color_data = Z;
		19'b1001100000101101100: color_data = Z;
		19'b1001100000101101110: color_data = Z;
		19'b1001100000101101111: color_data = Z;
		19'b1001100000101111101: color_data = Z;
		19'b1001100000101111110: color_data = Z;
		19'b1001100000101111111: color_data = Z;
		19'b1001100000110000000: color_data = Z;
		19'b1001100000110000001: color_data = Z;
		19'b1001100000110000010: color_data = Z;
		19'b1001100000110000011: color_data = Z;
		19'b1001100000110000100: color_data = Z;
		19'b1001100000110110000: color_data = Z;
		19'b1001100000110110001: color_data = Z;
		19'b1001100000110110010: color_data = Z;
		19'b1001100000110110110: color_data = Z;
		19'b1001100000110110111: color_data = Z;
		19'b1001100000111000110: color_data = Z;
		19'b1001100010011001011: color_data = Z;
		19'b1001100010011010100: color_data = Z;
		19'b1001100010011010101: color_data = Z;
		19'b1001100010011010110: color_data = Z;
		19'b1001100010011010111: color_data = Z;
		19'b1001100010011011000: color_data = Z;
		19'b1001100010011011001: color_data = Z;
		19'b1001100010011011010: color_data = Z;
		19'b1001100010011011011: color_data = Z;
		19'b1001100010011011100: color_data = Z;
		19'b1001100010011011101: color_data = Z;
		19'b1001100010011011110: color_data = Z;
		19'b1001100010011011111: color_data = Z;
		19'b1001100010011100000: color_data = Z;
		19'b1001100010011100001: color_data = Z;
		19'b1001100010011100010: color_data = Z;
		19'b1001100010011100011: color_data = Z;
		19'b1001100010011100100: color_data = Z;
		19'b1001100010011100101: color_data = Z;
		19'b1001100010011100110: color_data = Z;
		19'b1001100010011100111: color_data = Z;
		19'b1001100010011101000: color_data = Z;
		19'b1001100010011101001: color_data = Z;
		19'b1001100010011101010: color_data = Z;
		19'b1001100010100000111: color_data = Z;
		19'b1001100010100001000: color_data = Z;
		19'b1001100010100001001: color_data = Z;
		19'b1001100010100001010: color_data = Z;
		19'b1001100010100001011: color_data = Z;
		19'b1001100010100001100: color_data = Z;
		19'b1001100010100001101: color_data = Z;
		19'b1001100010100001110: color_data = Z;
		19'b1001100010100001111: color_data = Z;
		19'b1001100010100010000: color_data = Z;
		19'b1001100010100010001: color_data = Z;
		19'b1001100010100010010: color_data = Z;
		19'b1001100010100010011: color_data = Z;
		19'b1001100010100010100: color_data = Z;
		19'b1001100010101010001: color_data = Z;
		19'b1001100010101010010: color_data = Z;
		19'b1001100010101010100: color_data = Z;
		19'b1001100010101010101: color_data = Z;
		19'b1001100010101010110: color_data = Z;
		19'b1001100010101011100: color_data = Z;
		19'b1001100010101011101: color_data = Z;
		19'b1001100010101011110: color_data = Z;
		19'b1001100010101100010: color_data = Z;
		19'b1001100010101100011: color_data = Z;
		19'b1001100010101100100: color_data = Z;
		19'b1001100010101100101: color_data = Z;
		19'b1001100010101100110: color_data = Z;
		19'b1001100010101100111: color_data = Z;
		19'b1001100010101101000: color_data = Z;
		19'b1001100010101101001: color_data = Z;
		19'b1001100010101101010: color_data = Z;
		19'b1001100010101101011: color_data = Z;
		19'b1001100010101101100: color_data = Z;
		19'b1001100010101101101: color_data = Z;
		19'b1001100010101101110: color_data = Z;
		19'b1001100010101101111: color_data = Z;
		19'b1001100010101111101: color_data = Z;
		19'b1001100010101111110: color_data = Z;
		19'b1001100010101111111: color_data = Z;
		19'b1001100010110000000: color_data = Z;
		19'b1001100010110000001: color_data = Z;
		19'b1001100010110000010: color_data = Z;
		19'b1001100010110000011: color_data = Z;
		19'b1001100010110000100: color_data = Z;
		19'b1001100010110110000: color_data = Z;
		19'b1001100010110110001: color_data = Z;
		19'b1001100010110110010: color_data = Z;
		19'b1001100010110110110: color_data = Z;
		19'b1001100010110110111: color_data = Z;
		19'b1001100010111000110: color_data = Z;
		19'b1001100010111000111: color_data = Z;
		19'b1001100100011001011: color_data = Z;
		19'b1001100100011001100: color_data = Z;
		19'b1001100100011010100: color_data = Z;
		19'b1001100100011010101: color_data = Z;
		19'b1001100100011010110: color_data = Z;
		19'b1001100100011010111: color_data = Z;
		19'b1001100100011011000: color_data = Z;
		19'b1001100100011011001: color_data = Z;
		19'b1001100100011011010: color_data = Z;
		19'b1001100100011011011: color_data = Z;
		19'b1001100100011011100: color_data = Z;
		19'b1001100100011011101: color_data = Z;
		19'b1001100100011011110: color_data = Z;
		19'b1001100100011011111: color_data = Z;
		19'b1001100100011100000: color_data = Z;
		19'b1001100100011100001: color_data = Z;
		19'b1001100100011100010: color_data = Z;
		19'b1001100100011100100: color_data = Z;
		19'b1001100100011100101: color_data = Z;
		19'b1001100100011100110: color_data = Z;
		19'b1001100100011100111: color_data = Z;
		19'b1001100100011101000: color_data = Z;
		19'b1001100100011101001: color_data = Z;
		19'b1001100100011101010: color_data = Z;
		19'b1001100100100001000: color_data = Z;
		19'b1001100100100001001: color_data = Z;
		19'b1001100100100001010: color_data = Z;
		19'b1001100100100001011: color_data = Z;
		19'b1001100100100001100: color_data = Z;
		19'b1001100100100001101: color_data = Z;
		19'b1001100100100001110: color_data = Z;
		19'b1001100100100001111: color_data = Z;
		19'b1001100100100010000: color_data = Z;
		19'b1001100100100010001: color_data = Z;
		19'b1001100100100010010: color_data = Z;
		19'b1001100100100010011: color_data = Z;
		19'b1001100100100010100: color_data = Z;
		19'b1001100100101010000: color_data = Z;
		19'b1001100100101010001: color_data = Z;
		19'b1001100100101010010: color_data = Z;
		19'b1001100100101010011: color_data = Z;
		19'b1001100100101010100: color_data = Z;
		19'b1001100100101010101: color_data = Z;
		19'b1001100100101010110: color_data = Z;
		19'b1001100100101011001: color_data = Z;
		19'b1001100100101011010: color_data = Z;
		19'b1001100100101011011: color_data = Z;
		19'b1001100100101011100: color_data = Z;
		19'b1001100100101011101: color_data = Z;
		19'b1001100100101011110: color_data = Z;
		19'b1001100100101100010: color_data = Z;
		19'b1001100100101100011: color_data = Z;
		19'b1001100100101100100: color_data = Z;
		19'b1001100100101100101: color_data = Z;
		19'b1001100100101100110: color_data = Z;
		19'b1001100100101100111: color_data = Z;
		19'b1001100100101101000: color_data = Z;
		19'b1001100100101101001: color_data = Z;
		19'b1001100100101101010: color_data = Z;
		19'b1001100100101101011: color_data = Z;
		19'b1001100100101101100: color_data = Z;
		19'b1001100100101101101: color_data = Z;
		19'b1001100100101101110: color_data = Z;
		19'b1001100100101101111: color_data = Z;
		19'b1001100100101110001: color_data = Z;
		19'b1001100100101111101: color_data = Z;
		19'b1001100100101111110: color_data = Z;
		19'b1001100100101111111: color_data = Z;
		19'b1001100100110000000: color_data = Z;
		19'b1001100100110000001: color_data = Z;
		19'b1001100100110000010: color_data = Z;
		19'b1001100100110000011: color_data = Z;
		19'b1001100100110110000: color_data = Z;
		19'b1001100100110110001: color_data = Z;
		19'b1001100100110110110: color_data = Z;
		19'b1001100100110110111: color_data = Z;
		19'b1001100100111000110: color_data = Z;
		19'b1001100100111000111: color_data = Z;
		19'b1001100110011001100: color_data = Z;
		19'b1001100110011010100: color_data = Z;
		19'b1001100110011010101: color_data = Z;
		19'b1001100110011010110: color_data = Z;
		19'b1001100110011010111: color_data = Z;
		19'b1001100110011011000: color_data = Z;
		19'b1001100110011011001: color_data = Z;
		19'b1001100110011011010: color_data = Z;
		19'b1001100110011011011: color_data = Z;
		19'b1001100110011011100: color_data = Z;
		19'b1001100110011011101: color_data = Z;
		19'b1001100110011011110: color_data = Z;
		19'b1001100110011011111: color_data = Z;
		19'b1001100110011100000: color_data = Z;
		19'b1001100110011100001: color_data = Z;
		19'b1001100110011100101: color_data = Z;
		19'b1001100110011100110: color_data = Z;
		19'b1001100110011100111: color_data = Z;
		19'b1001100110011101000: color_data = Z;
		19'b1001100110011101001: color_data = Z;
		19'b1001100110011101010: color_data = Z;
		19'b1001100110100001001: color_data = Z;
		19'b1001100110100001010: color_data = Z;
		19'b1001100110100001011: color_data = Z;
		19'b1001100110100001100: color_data = Z;
		19'b1001100110100001101: color_data = Z;
		19'b1001100110100001110: color_data = Z;
		19'b1001100110100001111: color_data = Z;
		19'b1001100110100010000: color_data = Z;
		19'b1001100110100010001: color_data = Z;
		19'b1001100110100010010: color_data = Z;
		19'b1001100110100010011: color_data = Z;
		19'b1001100110100010100: color_data = Z;
		19'b1001100110101001111: color_data = Z;
		19'b1001100110101010000: color_data = Z;
		19'b1001100110101010001: color_data = Z;
		19'b1001100110101010010: color_data = Z;
		19'b1001100110101010011: color_data = Z;
		19'b1001100110101010100: color_data = Z;
		19'b1001100110101010101: color_data = Z;
		19'b1001100110101010110: color_data = Z;
		19'b1001100110101011000: color_data = Z;
		19'b1001100110101011001: color_data = Z;
		19'b1001100110101011010: color_data = Z;
		19'b1001100110101011011: color_data = Z;
		19'b1001100110101011100: color_data = Z;
		19'b1001100110101011101: color_data = Z;
		19'b1001100110101011110: color_data = Z;
		19'b1001100110101100010: color_data = Z;
		19'b1001100110101100011: color_data = Z;
		19'b1001100110101100100: color_data = Z;
		19'b1001100110101100101: color_data = Z;
		19'b1001100110101100110: color_data = Z;
		19'b1001100110101100111: color_data = Z;
		19'b1001100110101101000: color_data = Z;
		19'b1001100110101101001: color_data = Z;
		19'b1001100110101101010: color_data = Z;
		19'b1001100110101101011: color_data = Z;
		19'b1001100110101101100: color_data = Z;
		19'b1001100110101101101: color_data = Z;
		19'b1001100110101101110: color_data = Z;
		19'b1001100110101101111: color_data = Z;
		19'b1001100110110000000: color_data = Z;
		19'b1001100110110000001: color_data = Z;
		19'b1001100110110101111: color_data = Z;
		19'b1001100110110110000: color_data = Z;
		19'b1001100110110110001: color_data = Z;
		19'b1001100110110110110: color_data = Z;
		19'b1001100110110110111: color_data = Z;
		19'b1001100110111000101: color_data = Z;
		19'b1001100110111000110: color_data = Z;
		19'b1001100110111000111: color_data = Z;
		19'b1001101000011001100: color_data = Z;
		19'b1001101000011010101: color_data = Z;
		19'b1001101000011010110: color_data = Z;
		19'b1001101000011010111: color_data = Z;
		19'b1001101000011011000: color_data = Z;
		19'b1001101000011011001: color_data = Z;
		19'b1001101000011011010: color_data = Z;
		19'b1001101000011011011: color_data = Z;
		19'b1001101000011011100: color_data = Z;
		19'b1001101000011011101: color_data = Z;
		19'b1001101000011011110: color_data = Z;
		19'b1001101000011011111: color_data = Z;
		19'b1001101000011100000: color_data = Z;
		19'b1001101000011100001: color_data = Z;
		19'b1001101000011100101: color_data = Z;
		19'b1001101000011100110: color_data = Z;
		19'b1001101000011100111: color_data = Z;
		19'b1001101000011101000: color_data = Z;
		19'b1001101000011101001: color_data = Z;
		19'b1001101000011101010: color_data = Z;
		19'b1001101000100001101: color_data = Z;
		19'b1001101000100001110: color_data = Z;
		19'b1001101000100001111: color_data = Z;
		19'b1001101000100010000: color_data = Z;
		19'b1001101000100010001: color_data = Z;
		19'b1001101000100010010: color_data = Z;
		19'b1001101000100010011: color_data = Z;
		19'b1001101000100010100: color_data = Z;
		19'b1001101000100110100: color_data = Z;
		19'b1001101000101001111: color_data = Z;
		19'b1001101000101010000: color_data = Z;
		19'b1001101000101010001: color_data = Z;
		19'b1001101000101010010: color_data = Z;
		19'b1001101000101010011: color_data = Z;
		19'b1001101000101010100: color_data = Z;
		19'b1001101000101010101: color_data = Z;
		19'b1001101000101010110: color_data = Z;
		19'b1001101000101010111: color_data = Z;
		19'b1001101000101011000: color_data = Z;
		19'b1001101000101011001: color_data = Z;
		19'b1001101000101011010: color_data = Z;
		19'b1001101000101011011: color_data = Z;
		19'b1001101000101011100: color_data = Z;
		19'b1001101000101011101: color_data = Z;
		19'b1001101000101100010: color_data = Z;
		19'b1001101000101100011: color_data = Z;
		19'b1001101000101100100: color_data = Z;
		19'b1001101000101100101: color_data = Z;
		19'b1001101000101100110: color_data = Z;
		19'b1001101000101100111: color_data = Z;
		19'b1001101000101101000: color_data = Z;
		19'b1001101000101101001: color_data = Z;
		19'b1001101000101101010: color_data = Z;
		19'b1001101000101101011: color_data = Z;
		19'b1001101000101101100: color_data = Z;
		19'b1001101000101101101: color_data = Z;
		19'b1001101000101101110: color_data = Z;
		19'b1001101000101101111: color_data = Z;
		19'b1001101000110101111: color_data = Z;
		19'b1001101000110110000: color_data = Z;
		19'b1001101000110110001: color_data = Z;
		19'b1001101000110110110: color_data = Z;
		19'b1001101000110110111: color_data = Z;
		19'b1001101000111000101: color_data = Z;
		19'b1001101000111000110: color_data = Z;
		19'b1001101010011001100: color_data = Z;
		19'b1001101010011010101: color_data = Z;
		19'b1001101010011010110: color_data = Z;
		19'b1001101010011010111: color_data = Z;
		19'b1001101010011011000: color_data = Z;
		19'b1001101010011011001: color_data = Z;
		19'b1001101010011011010: color_data = Z;
		19'b1001101010011011011: color_data = Z;
		19'b1001101010011011100: color_data = Z;
		19'b1001101010011011101: color_data = Z;
		19'b1001101010011011110: color_data = Z;
		19'b1001101010011011111: color_data = Z;
		19'b1001101010011100000: color_data = Z;
		19'b1001101010011100001: color_data = Z;
		19'b1001101010011100010: color_data = Z;
		19'b1001101010011100110: color_data = Z;
		19'b1001101010011100111: color_data = Z;
		19'b1001101010011101000: color_data = Z;
		19'b1001101010011101001: color_data = Z;
		19'b1001101010100001110: color_data = Z;
		19'b1001101010100001111: color_data = Z;
		19'b1001101010100010000: color_data = Z;
		19'b1001101010100010001: color_data = Z;
		19'b1001101010100010010: color_data = Z;
		19'b1001101010100010011: color_data = Z;
		19'b1001101010100010100: color_data = Z;
		19'b1001101010100100101: color_data = Z;
		19'b1001101010100100110: color_data = Z;
		19'b1001101010100101001: color_data = Z;
		19'b1001101010100111010: color_data = Z;
		19'b1001101010101001001: color_data = Z;
		19'b1001101010101001111: color_data = Z;
		19'b1001101010101010000: color_data = Z;
		19'b1001101010101010001: color_data = Z;
		19'b1001101010101010010: color_data = Z;
		19'b1001101010101010011: color_data = Z;
		19'b1001101010101010100: color_data = Z;
		19'b1001101010101010101: color_data = Z;
		19'b1001101010101010110: color_data = Z;
		19'b1001101010101010111: color_data = Z;
		19'b1001101010101011000: color_data = Z;
		19'b1001101010101011001: color_data = Z;
		19'b1001101010101011010: color_data = Z;
		19'b1001101010101011011: color_data = Z;
		19'b1001101010101011100: color_data = Z;
		19'b1001101010101011101: color_data = Z;
		19'b1001101010101100010: color_data = Z;
		19'b1001101010101100011: color_data = Z;
		19'b1001101010101100100: color_data = Z;
		19'b1001101010101100101: color_data = Z;
		19'b1001101010101100110: color_data = Z;
		19'b1001101010101100111: color_data = Z;
		19'b1001101010101101000: color_data = Z;
		19'b1001101010101101001: color_data = Z;
		19'b1001101010101101010: color_data = Z;
		19'b1001101010101101011: color_data = Z;
		19'b1001101010101101100: color_data = Z;
		19'b1001101010101101101: color_data = Z;
		19'b1001101010101101110: color_data = Z;
		19'b1001101010101101111: color_data = Z;
		19'b1001101010110101111: color_data = Z;
		19'b1001101010110110000: color_data = Z;
		19'b1001101010110110001: color_data = Z;
		19'b1001101010110110101: color_data = Z;
		19'b1001101010110110110: color_data = Z;
		19'b1001101010110110111: color_data = Z;
		19'b1001101010111000101: color_data = Z;
		19'b1001101010111000110: color_data = Z;
		19'b1001101100011001101: color_data = Z;
		19'b1001101100011010101: color_data = Z;
		19'b1001101100011010110: color_data = Z;
		19'b1001101100011010111: color_data = Z;
		19'b1001101100011011000: color_data = Z;
		19'b1001101100011011001: color_data = Z;
		19'b1001101100011011010: color_data = Z;
		19'b1001101100011011011: color_data = Z;
		19'b1001101100011011100: color_data = Z;
		19'b1001101100011011101: color_data = Z;
		19'b1001101100011011110: color_data = Z;
		19'b1001101100011011111: color_data = Z;
		19'b1001101100011100000: color_data = Z;
		19'b1001101100011100001: color_data = Z;
		19'b1001101100011100010: color_data = Z;
		19'b1001101100011100110: color_data = Z;
		19'b1001101100011100111: color_data = Z;
		19'b1001101100011101000: color_data = Z;
		19'b1001101100011101001: color_data = Z;
		19'b1001101100100001111: color_data = Z;
		19'b1001101100100010000: color_data = Z;
		19'b1001101100100010001: color_data = Z;
		19'b1001101100100010010: color_data = Z;
		19'b1001101100100010011: color_data = Z;
		19'b1001101100100100010: color_data = Z;
		19'b1001101100100100100: color_data = Z;
		19'b1001101100100100101: color_data = Z;
		19'b1001101100100100110: color_data = Z;
		19'b1001101100100100111: color_data = Z;
		19'b1001101100100101001: color_data = Z;
		19'b1001101100100101010: color_data = Z;
		19'b1001101100100111010: color_data = Z;
		19'b1001101100101000001: color_data = Z;
		19'b1001101100101000010: color_data = Z;
		19'b1001101100101000011: color_data = Z;
		19'b1001101100101000100: color_data = Z;
		19'b1001101100101001001: color_data = Z;
		19'b1001101100101001110: color_data = Z;
		19'b1001101100101001111: color_data = Z;
		19'b1001101100101010000: color_data = Z;
		19'b1001101100101010001: color_data = Z;
		19'b1001101100101010010: color_data = Z;
		19'b1001101100101010011: color_data = Z;
		19'b1001101100101010100: color_data = Z;
		19'b1001101100101010101: color_data = Z;
		19'b1001101100101010110: color_data = Z;
		19'b1001101100101010111: color_data = Z;
		19'b1001101100101011000: color_data = Z;
		19'b1001101100101011001: color_data = Z;
		19'b1001101100101011010: color_data = Z;
		19'b1001101100101011011: color_data = Z;
		19'b1001101100101011100: color_data = Z;
		19'b1001101100101011101: color_data = Z;
		19'b1001101100101100010: color_data = Z;
		19'b1001101100101100011: color_data = Z;
		19'b1001101100101100100: color_data = Z;
		19'b1001101100101100101: color_data = Z;
		19'b1001101100101100110: color_data = Z;
		19'b1001101100101100111: color_data = Z;
		19'b1001101100101101000: color_data = Z;
		19'b1001101100101101001: color_data = Z;
		19'b1001101100101101010: color_data = Z;
		19'b1001101100101101011: color_data = Z;
		19'b1001101100101101100: color_data = Z;
		19'b1001101100101101101: color_data = Z;
		19'b1001101100101101110: color_data = Z;
		19'b1001101100101101111: color_data = Z;
		19'b1001101100110101111: color_data = Z;
		19'b1001101100110110000: color_data = Z;
		19'b1001101100110110001: color_data = Z;
		19'b1001101100110110101: color_data = Z;
		19'b1001101100110110110: color_data = Z;
		19'b1001101100110110111: color_data = Z;
		19'b1001101100111000101: color_data = Z;
		19'b1001101100111000110: color_data = Z;
		19'b1001101110011001101: color_data = Z;
		19'b1001101110011001110: color_data = Z;
		19'b1001101110011010101: color_data = Z;
		19'b1001101110011010110: color_data = Z;
		19'b1001101110011010111: color_data = Z;
		19'b1001101110011011000: color_data = Z;
		19'b1001101110011011001: color_data = Z;
		19'b1001101110011011010: color_data = Z;
		19'b1001101110011011011: color_data = Z;
		19'b1001101110011011100: color_data = Z;
		19'b1001101110011011101: color_data = Z;
		19'b1001101110011011110: color_data = Z;
		19'b1001101110011011111: color_data = Z;
		19'b1001101110011100000: color_data = Z;
		19'b1001101110011100001: color_data = Z;
		19'b1001101110011100010: color_data = Z;
		19'b1001101110011100110: color_data = Z;
		19'b1001101110011100111: color_data = Z;
		19'b1001101110011101000: color_data = Z;
		19'b1001101110100010000: color_data = Z;
		19'b1001101110100010001: color_data = Z;
		19'b1001101110100010010: color_data = Z;
		19'b1001101110100100010: color_data = Z;
		19'b1001101110100100011: color_data = Z;
		19'b1001101110100100100: color_data = Z;
		19'b1001101110100100101: color_data = Z;
		19'b1001101110100100110: color_data = Z;
		19'b1001101110100100111: color_data = Z;
		19'b1001101110100101010: color_data = Z;
		19'b1001101110100101011: color_data = Z;
		19'b1001101110100111010: color_data = Z;
		19'b1001101110100111011: color_data = Z;
		19'b1001101110101000001: color_data = Z;
		19'b1001101110101000010: color_data = Z;
		19'b1001101110101000011: color_data = Z;
		19'b1001101110101000100: color_data = Z;
		19'b1001101110101000101: color_data = Z;
		19'b1001101110101001111: color_data = Z;
		19'b1001101110101010000: color_data = Z;
		19'b1001101110101010001: color_data = Z;
		19'b1001101110101010010: color_data = Z;
		19'b1001101110101010011: color_data = Z;
		19'b1001101110101010100: color_data = Z;
		19'b1001101110101010101: color_data = Z;
		19'b1001101110101010110: color_data = Z;
		19'b1001101110101010111: color_data = Z;
		19'b1001101110101011000: color_data = Z;
		19'b1001101110101011001: color_data = Z;
		19'b1001101110101011010: color_data = Z;
		19'b1001101110101011011: color_data = Z;
		19'b1001101110101011100: color_data = Z;
		19'b1001101110101100010: color_data = Z;
		19'b1001101110101100011: color_data = Z;
		19'b1001101110101100100: color_data = Z;
		19'b1001101110101100101: color_data = Z;
		19'b1001101110101100110: color_data = Z;
		19'b1001101110101100111: color_data = Z;
		19'b1001101110101101000: color_data = Z;
		19'b1001101110101101001: color_data = Z;
		19'b1001101110101101010: color_data = Z;
		19'b1001101110101101011: color_data = Z;
		19'b1001101110101101100: color_data = Z;
		19'b1001101110101101101: color_data = Z;
		19'b1001101110101101110: color_data = Z;
		19'b1001101110101101111: color_data = Z;
		19'b1001101110110101110: color_data = Z;
		19'b1001101110110101111: color_data = Z;
		19'b1001101110110110000: color_data = Z;
		19'b1001101110110110001: color_data = Z;
		19'b1001101110110110101: color_data = Z;
		19'b1001101110110110110: color_data = Z;
		19'b1001101110110110111: color_data = Z;
		19'b1001101110111000101: color_data = Z;
		19'b1001110000011001110: color_data = Z;
		19'b1001110000011010101: color_data = Z;
		19'b1001110000011010110: color_data = Z;
		19'b1001110000011010111: color_data = Z;
		19'b1001110000011011000: color_data = Z;
		19'b1001110000011011001: color_data = Z;
		19'b1001110000011011010: color_data = Z;
		19'b1001110000011011011: color_data = Z;
		19'b1001110000011011100: color_data = Z;
		19'b1001110000011011101: color_data = Z;
		19'b1001110000011011110: color_data = Z;
		19'b1001110000011011111: color_data = Z;
		19'b1001110000011100000: color_data = Z;
		19'b1001110000011100001: color_data = Z;
		19'b1001110000011100010: color_data = Z;
		19'b1001110000011100111: color_data = Z;
		19'b1001110000011101000: color_data = Z;
		19'b1001110000100100011: color_data = Z;
		19'b1001110000100100100: color_data = Z;
		19'b1001110000100100101: color_data = Z;
		19'b1001110000100100110: color_data = Z;
		19'b1001110000100100111: color_data = Z;
		19'b1001110000100101000: color_data = Z;
		19'b1001110000100101001: color_data = Z;
		19'b1001110000100101010: color_data = Z;
		19'b1001110000100101011: color_data = Z;
		19'b1001110000100101100: color_data = Z;
		19'b1001110000100110101: color_data = Z;
		19'b1001110000100111010: color_data = Z;
		19'b1001110000100111011: color_data = Z;
		19'b1001110000101000001: color_data = Z;
		19'b1001110000101000010: color_data = Z;
		19'b1001110000101000011: color_data = Z;
		19'b1001110000101000100: color_data = Z;
		19'b1001110000101000101: color_data = Z;
		19'b1001110000101010001: color_data = Z;
		19'b1001110000101010010: color_data = Z;
		19'b1001110000101010011: color_data = Z;
		19'b1001110000101010100: color_data = Z;
		19'b1001110000101010101: color_data = Z;
		19'b1001110000101010110: color_data = Z;
		19'b1001110000101010111: color_data = Z;
		19'b1001110000101011000: color_data = Z;
		19'b1001110000101011001: color_data = Z;
		19'b1001110000101011010: color_data = Z;
		19'b1001110000101011011: color_data = Z;
		19'b1001110000101011100: color_data = Z;
		19'b1001110000101100010: color_data = Z;
		19'b1001110000101100011: color_data = Z;
		19'b1001110000101100100: color_data = Z;
		19'b1001110000101100101: color_data = Z;
		19'b1001110000101100110: color_data = Z;
		19'b1001110000101100111: color_data = Z;
		19'b1001110000101101000: color_data = Z;
		19'b1001110000101101001: color_data = Z;
		19'b1001110000101101010: color_data = Z;
		19'b1001110000101101011: color_data = Z;
		19'b1001110000101101100: color_data = Z;
		19'b1001110000101101101: color_data = Z;
		19'b1001110000101101110: color_data = Z;
		19'b1001110000101101111: color_data = Z;
		19'b1001110000110101110: color_data = Z;
		19'b1001110000110101111: color_data = Z;
		19'b1001110000110110000: color_data = Z;
		19'b1001110000110110001: color_data = Z;
		19'b1001110000110110101: color_data = Z;
		19'b1001110000110110110: color_data = Z;
		19'b1001110000110110111: color_data = Z;
		19'b1001110000111000100: color_data = Z;
		19'b1001110000111000101: color_data = Z;
		19'b1001110010011001110: color_data = Z;
		19'b1001110010011010110: color_data = Z;
		19'b1001110010011010111: color_data = Z;
		19'b1001110010011011000: color_data = Z;
		19'b1001110010011011001: color_data = Z;
		19'b1001110010011011010: color_data = Z;
		19'b1001110010011011011: color_data = Z;
		19'b1001110010011011100: color_data = Z;
		19'b1001110010011011101: color_data = Z;
		19'b1001110010011011110: color_data = Z;
		19'b1001110010011011111: color_data = Z;
		19'b1001110010011100000: color_data = Z;
		19'b1001110010011100001: color_data = Z;
		19'b1001110010011100010: color_data = Z;
		19'b1001110010011100111: color_data = Z;
		19'b1001110010011101000: color_data = Z;
		19'b1001110010100100011: color_data = Z;
		19'b1001110010100100100: color_data = Z;
		19'b1001110010100100101: color_data = Z;
		19'b1001110010100100110: color_data = Z;
		19'b1001110010100100111: color_data = Z;
		19'b1001110010100101000: color_data = Z;
		19'b1001110010100101001: color_data = Z;
		19'b1001110010100101010: color_data = Z;
		19'b1001110010100101011: color_data = Z;
		19'b1001110010100101100: color_data = Z;
		19'b1001110010100110101: color_data = Z;
		19'b1001110010100110110: color_data = Z;
		19'b1001110010100110111: color_data = Z;
		19'b1001110010101000000: color_data = Z;
		19'b1001110010101000001: color_data = Z;
		19'b1001110010101000010: color_data = Z;
		19'b1001110010101000011: color_data = Z;
		19'b1001110010101000100: color_data = Z;
		19'b1001110010101000101: color_data = Z;
		19'b1001110010101000110: color_data = Z;
		19'b1001110010101000111: color_data = Z;
		19'b1001110010101010010: color_data = Z;
		19'b1001110010101010011: color_data = Z;
		19'b1001110010101010100: color_data = Z;
		19'b1001110010101010101: color_data = Z;
		19'b1001110010101010110: color_data = Z;
		19'b1001110010101010111: color_data = Z;
		19'b1001110010101011000: color_data = Z;
		19'b1001110010101011001: color_data = Z;
		19'b1001110010101011010: color_data = Z;
		19'b1001110010101011011: color_data = Z;
		19'b1001110010101100001: color_data = Z;
		19'b1001110010101100010: color_data = Z;
		19'b1001110010101100011: color_data = Z;
		19'b1001110010101100100: color_data = Z;
		19'b1001110010101100101: color_data = Z;
		19'b1001110010101100110: color_data = Z;
		19'b1001110010101100111: color_data = Z;
		19'b1001110010101101000: color_data = Z;
		19'b1001110010101101001: color_data = Z;
		19'b1001110010101101010: color_data = Z;
		19'b1001110010101101011: color_data = Z;
		19'b1001110010101101100: color_data = Z;
		19'b1001110010101101101: color_data = Z;
		19'b1001110010101101110: color_data = Z;
		19'b1001110010101101111: color_data = Z;
		19'b1001110010110101110: color_data = Z;
		19'b1001110010110101111: color_data = Z;
		19'b1001110010110110000: color_data = Z;
		19'b1001110010110110001: color_data = Z;
		19'b1001110010110110101: color_data = Z;
		19'b1001110010110110110: color_data = Z;
		19'b1001110010110110111: color_data = Z;
		19'b1001110010111000100: color_data = Z;
		19'b1001110100011001110: color_data = Z;
		19'b1001110100011001111: color_data = Z;
		19'b1001110100011010110: color_data = Z;
		19'b1001110100011010111: color_data = Z;
		19'b1001110100011011000: color_data = Z;
		19'b1001110100011011001: color_data = Z;
		19'b1001110100011011010: color_data = Z;
		19'b1001110100011011011: color_data = Z;
		19'b1001110100011011100: color_data = Z;
		19'b1001110100011011101: color_data = Z;
		19'b1001110100011011110: color_data = Z;
		19'b1001110100011011111: color_data = Z;
		19'b1001110100011100000: color_data = Z;
		19'b1001110100011100001: color_data = Z;
		19'b1001110100011100010: color_data = Z;
		19'b1001110100011100011: color_data = Z;
		19'b1001110100100100100: color_data = Z;
		19'b1001110100100100101: color_data = Z;
		19'b1001110100100100110: color_data = Z;
		19'b1001110100100100111: color_data = Z;
		19'b1001110100100101000: color_data = Z;
		19'b1001110100100101001: color_data = Z;
		19'b1001110100100101010: color_data = Z;
		19'b1001110100100101011: color_data = Z;
		19'b1001110100100101100: color_data = Z;
		19'b1001110100100101101: color_data = Z;
		19'b1001110100100110101: color_data = Z;
		19'b1001110100100110110: color_data = Z;
		19'b1001110100100110111: color_data = Z;
		19'b1001110100101000001: color_data = Z;
		19'b1001110100101000010: color_data = Z;
		19'b1001110100101000011: color_data = Z;
		19'b1001110100101000100: color_data = Z;
		19'b1001110100101000101: color_data = Z;
		19'b1001110100101000110: color_data = Z;
		19'b1001110100101000111: color_data = Z;
		19'b1001110100101001001: color_data = Z;
		19'b1001110100101001010: color_data = Z;
		19'b1001110100101010010: color_data = Z;
		19'b1001110100101010011: color_data = Z;
		19'b1001110100101010100: color_data = Z;
		19'b1001110100101010101: color_data = Z;
		19'b1001110100101010110: color_data = Z;
		19'b1001110100101010111: color_data = Z;
		19'b1001110100101011000: color_data = Z;
		19'b1001110100101011001: color_data = Z;
		19'b1001110100101011010: color_data = Z;
		19'b1001110100101100001: color_data = Z;
		19'b1001110100101100010: color_data = Z;
		19'b1001110100101100011: color_data = Z;
		19'b1001110100101100100: color_data = Z;
		19'b1001110100101100101: color_data = Z;
		19'b1001110100101100110: color_data = Z;
		19'b1001110100101100111: color_data = Z;
		19'b1001110100101101000: color_data = Z;
		19'b1001110100101101001: color_data = Z;
		19'b1001110100101101010: color_data = Z;
		19'b1001110100101101011: color_data = Z;
		19'b1001110100101101100: color_data = Z;
		19'b1001110100101101101: color_data = Z;
		19'b1001110100110101101: color_data = Z;
		19'b1001110100110101110: color_data = Z;
		19'b1001110100110101111: color_data = Z;
		19'b1001110100110110000: color_data = Z;
		19'b1001110100110110001: color_data = Z;
		19'b1001110100110110101: color_data = Z;
		19'b1001110100110110110: color_data = Z;
		19'b1001110100110110111: color_data = Z;
		19'b1001110100111000011: color_data = Z;
		19'b1001110110011010110: color_data = Z;
		19'b1001110110011010111: color_data = Z;
		19'b1001110110011011000: color_data = Z;
		19'b1001110110011011001: color_data = Z;
		19'b1001110110011011010: color_data = Z;
		19'b1001110110011011011: color_data = Z;
		19'b1001110110011011100: color_data = Z;
		19'b1001110110011011101: color_data = Z;
		19'b1001110110011011110: color_data = Z;
		19'b1001110110011011111: color_data = Z;
		19'b1001110110011100000: color_data = Z;
		19'b1001110110011100001: color_data = Z;
		19'b1001110110011100010: color_data = Z;
		19'b1001110110011100011: color_data = Z;
		19'b1001110110100100101: color_data = Z;
		19'b1001110110100100110: color_data = Z;
		19'b1001110110100100111: color_data = Z;
		19'b1001110110100101000: color_data = Z;
		19'b1001110110100101001: color_data = Z;
		19'b1001110110100101010: color_data = Z;
		19'b1001110110100101011: color_data = Z;
		19'b1001110110100101100: color_data = Z;
		19'b1001110110100101101: color_data = Z;
		19'b1001110110100101110: color_data = Z;
		19'b1001110110100101111: color_data = Z;
		19'b1001110110100110000: color_data = Z;
		19'b1001110110100110101: color_data = Z;
		19'b1001110110100110110: color_data = Z;
		19'b1001110110100110111: color_data = Z;
		19'b1001110110100111000: color_data = Z;
		19'b1001110110101000001: color_data = Z;
		19'b1001110110101000010: color_data = Z;
		19'b1001110110101000011: color_data = Z;
		19'b1001110110101000100: color_data = Z;
		19'b1001110110101000101: color_data = Z;
		19'b1001110110101000110: color_data = Z;
		19'b1001110110101000111: color_data = Z;
		19'b1001110110101001000: color_data = Z;
		19'b1001110110101001001: color_data = Z;
		19'b1001110110101001010: color_data = Z;
		19'b1001110110101010010: color_data = Z;
		19'b1001110110101010011: color_data = Z;
		19'b1001110110101010100: color_data = Z;
		19'b1001110110101010101: color_data = Z;
		19'b1001110110101010110: color_data = Z;
		19'b1001110110101010111: color_data = Z;
		19'b1001110110101011000: color_data = Z;
		19'b1001110110101011001: color_data = Z;
		19'b1001110110101011010: color_data = Z;
		19'b1001110110101100001: color_data = Z;
		19'b1001110110101100010: color_data = Z;
		19'b1001110110101100011: color_data = Z;
		19'b1001110110101100100: color_data = Z;
		19'b1001110110101100101: color_data = Z;
		19'b1001110110101100110: color_data = Z;
		19'b1001110110101100111: color_data = Z;
		19'b1001110110101101000: color_data = Z;
		19'b1001110110101101001: color_data = Z;
		19'b1001110110101101010: color_data = Z;
		19'b1001110110101101011: color_data = Z;
		19'b1001110110101101100: color_data = Z;
		19'b1001110110110101101: color_data = Z;
		19'b1001110110110101110: color_data = Z;
		19'b1001110110110101111: color_data = Z;
		19'b1001110110110110000: color_data = Z;
		19'b1001110110110110001: color_data = Z;
		19'b1001110110110110100: color_data = Z;
		19'b1001110110110110101: color_data = Z;
		19'b1001110110110110110: color_data = Z;
		19'b1001110110111000011: color_data = Z;
		19'b1001111000011010110: color_data = Z;
		19'b1001111000011010111: color_data = Z;
		19'b1001111000011011000: color_data = Z;
		19'b1001111000011011001: color_data = Z;
		19'b1001111000011011010: color_data = Z;
		19'b1001111000011011011: color_data = Z;
		19'b1001111000011011100: color_data = Z;
		19'b1001111000011011101: color_data = Z;
		19'b1001111000011011110: color_data = Z;
		19'b1001111000011011111: color_data = Z;
		19'b1001111000011100000: color_data = Z;
		19'b1001111000011100001: color_data = Z;
		19'b1001111000011100010: color_data = Z;
		19'b1001111000011100011: color_data = Z;
		19'b1001111000100100110: color_data = Z;
		19'b1001111000100100111: color_data = Z;
		19'b1001111000100101000: color_data = Z;
		19'b1001111000100101001: color_data = Z;
		19'b1001111000100101010: color_data = Z;
		19'b1001111000100101011: color_data = Z;
		19'b1001111000100101100: color_data = Z;
		19'b1001111000100101101: color_data = Z;
		19'b1001111000100101110: color_data = Z;
		19'b1001111000100101111: color_data = Z;
		19'b1001111000100110000: color_data = Z;
		19'b1001111000100110101: color_data = Z;
		19'b1001111000100110110: color_data = Z;
		19'b1001111000100110111: color_data = Z;
		19'b1001111000100111000: color_data = Z;
		19'b1001111000100111001: color_data = Z;
		19'b1001111000100111011: color_data = Z;
		19'b1001111000101000001: color_data = Z;
		19'b1001111000101000010: color_data = Z;
		19'b1001111000101000011: color_data = Z;
		19'b1001111000101000100: color_data = Z;
		19'b1001111000101000101: color_data = Z;
		19'b1001111000101000110: color_data = Z;
		19'b1001111000101000111: color_data = Z;
		19'b1001111000101001000: color_data = Z;
		19'b1001111000101001001: color_data = Z;
		19'b1001111000101001010: color_data = Z;
		19'b1001111000101001011: color_data = Z;
		19'b1001111000101010010: color_data = Z;
		19'b1001111000101010011: color_data = Z;
		19'b1001111000101010100: color_data = Z;
		19'b1001111000101010101: color_data = Z;
		19'b1001111000101010110: color_data = Z;
		19'b1001111000101010111: color_data = Z;
		19'b1001111000101011000: color_data = Z;
		19'b1001111000101011001: color_data = Z;
		19'b1001111000101100001: color_data = Z;
		19'b1001111000101100010: color_data = Z;
		19'b1001111000101100011: color_data = Z;
		19'b1001111000101100100: color_data = Z;
		19'b1001111000101100101: color_data = Z;
		19'b1001111000101100110: color_data = Z;
		19'b1001111000101100111: color_data = Z;
		19'b1001111000101101001: color_data = Z;
		19'b1001111000101101010: color_data = Z;
		19'b1001111000101101011: color_data = Z;
		19'b1001111000110101100: color_data = Z;
		19'b1001111000110101101: color_data = Z;
		19'b1001111000110101110: color_data = Z;
		19'b1001111000110101111: color_data = Z;
		19'b1001111000110110000: color_data = Z;
		19'b1001111000110110100: color_data = Z;
		19'b1001111000110110101: color_data = Z;
		19'b1001111000110110110: color_data = Z;
		19'b1001111000110111100: color_data = Z;
		19'b1001111010011010110: color_data = Z;
		19'b1001111010011010111: color_data = Z;
		19'b1001111010011011000: color_data = Z;
		19'b1001111010011011001: color_data = Z;
		19'b1001111010011011010: color_data = Z;
		19'b1001111010011011011: color_data = Z;
		19'b1001111010011011100: color_data = Z;
		19'b1001111010011011101: color_data = Z;
		19'b1001111010011011110: color_data = Z;
		19'b1001111010011011111: color_data = Z;
		19'b1001111010011100000: color_data = Z;
		19'b1001111010011100001: color_data = Z;
		19'b1001111010011100010: color_data = Z;
		19'b1001111010011100011: color_data = Z;
		19'b1001111010100101000: color_data = Z;
		19'b1001111010100101001: color_data = Z;
		19'b1001111010100101010: color_data = Z;
		19'b1001111010100101011: color_data = Z;
		19'b1001111010100101100: color_data = Z;
		19'b1001111010100101101: color_data = Z;
		19'b1001111010100101110: color_data = Z;
		19'b1001111010100101111: color_data = Z;
		19'b1001111010100110101: color_data = Z;
		19'b1001111010100110110: color_data = Z;
		19'b1001111010100110111: color_data = Z;
		19'b1001111010100111000: color_data = Z;
		19'b1001111010100111001: color_data = Z;
		19'b1001111010100111010: color_data = Z;
		19'b1001111010100111011: color_data = Z;
		19'b1001111010101000001: color_data = Z;
		19'b1001111010101000010: color_data = Z;
		19'b1001111010101000011: color_data = Z;
		19'b1001111010101000100: color_data = Z;
		19'b1001111010101000101: color_data = Z;
		19'b1001111010101000110: color_data = Z;
		19'b1001111010101000111: color_data = Z;
		19'b1001111010101001000: color_data = Z;
		19'b1001111010101001001: color_data = Z;
		19'b1001111010101001010: color_data = Z;
		19'b1001111010101001011: color_data = Z;
		19'b1001111010101010010: color_data = Z;
		19'b1001111010101010011: color_data = Z;
		19'b1001111010101010100: color_data = Z;
		19'b1001111010101010101: color_data = Z;
		19'b1001111010101010110: color_data = Z;
		19'b1001111010101010111: color_data = Z;
		19'b1001111010101011000: color_data = Z;
		19'b1001111010101100001: color_data = Z;
		19'b1001111010101100010: color_data = Z;
		19'b1001111010101100011: color_data = Z;
		19'b1001111010101100100: color_data = Z;
		19'b1001111010101100101: color_data = Z;
		19'b1001111010110101100: color_data = Z;
		19'b1001111010110101101: color_data = Z;
		19'b1001111010110101110: color_data = Z;
		19'b1001111010110101111: color_data = Z;
		19'b1001111010110110000: color_data = Z;
		19'b1001111010110110100: color_data = Z;
		19'b1001111010110110101: color_data = Z;
		19'b1001111010110110110: color_data = Z;
		19'b1001111010110111100: color_data = Z;
		19'b1001111100011000101: color_data = Z;
		19'b1001111100011010111: color_data = Z;
		19'b1001111100011011000: color_data = Z;
		19'b1001111100011011001: color_data = Z;
		19'b1001111100011011010: color_data = Z;
		19'b1001111100011011011: color_data = Z;
		19'b1001111100011011100: color_data = Z;
		19'b1001111100011011101: color_data = Z;
		19'b1001111100011011110: color_data = Z;
		19'b1001111100011011111: color_data = Z;
		19'b1001111100011100000: color_data = Z;
		19'b1001111100011100001: color_data = Z;
		19'b1001111100011100010: color_data = Z;
		19'b1001111100011100011: color_data = Z;
		19'b1001111100100101100: color_data = Z;
		19'b1001111100100101101: color_data = Z;
		19'b1001111100100101110: color_data = Z;
		19'b1001111100100110101: color_data = Z;
		19'b1001111100100110110: color_data = Z;
		19'b1001111100100110111: color_data = Z;
		19'b1001111100100111000: color_data = Z;
		19'b1001111100100111001: color_data = Z;
		19'b1001111100100111010: color_data = Z;
		19'b1001111100100111011: color_data = Z;
		19'b1001111100100111100: color_data = Z;
		19'b1001111100101000001: color_data = Z;
		19'b1001111100101000010: color_data = Z;
		19'b1001111100101000011: color_data = Z;
		19'b1001111100101000100: color_data = Z;
		19'b1001111100101000101: color_data = Z;
		19'b1001111100101000110: color_data = Z;
		19'b1001111100101000111: color_data = Z;
		19'b1001111100101001000: color_data = Z;
		19'b1001111100101001001: color_data = Z;
		19'b1001111100101001010: color_data = Z;
		19'b1001111100101010010: color_data = Z;
		19'b1001111100101010011: color_data = Z;
		19'b1001111100101010100: color_data = Z;
		19'b1001111100101010101: color_data = Z;
		19'b1001111100101010110: color_data = Z;
		19'b1001111100101010111: color_data = Z;
		19'b1001111100101011000: color_data = Z;
		19'b1001111100101100010: color_data = Z;
		19'b1001111100101100011: color_data = Z;
		19'b1001111100101100100: color_data = Z;
		19'b1001111100101100101: color_data = Z;
		19'b1001111100110101011: color_data = Z;
		19'b1001111100110101100: color_data = Z;
		19'b1001111100110101101: color_data = Z;
		19'b1001111100110101110: color_data = Z;
		19'b1001111100110101111: color_data = Z;
		19'b1001111100110110000: color_data = Z;
		19'b1001111100110110100: color_data = Z;
		19'b1001111100110110101: color_data = Z;
		19'b1001111100110110110: color_data = Z;
		19'b1001111100110111011: color_data = Z;
		19'b1001111110011000110: color_data = Z;
		19'b1001111110011010111: color_data = Z;
		19'b1001111110011011000: color_data = Z;
		19'b1001111110011011001: color_data = Z;
		19'b1001111110011011010: color_data = Z;
		19'b1001111110011011011: color_data = Z;
		19'b1001111110011011100: color_data = Z;
		19'b1001111110011011101: color_data = Z;
		19'b1001111110011011110: color_data = Z;
		19'b1001111110011011111: color_data = Z;
		19'b1001111110011100000: color_data = Z;
		19'b1001111110011100001: color_data = Z;
		19'b1001111110011100010: color_data = Z;
		19'b1001111110011100011: color_data = Z;
		19'b1001111110100110101: color_data = Z;
		19'b1001111110100110110: color_data = Z;
		19'b1001111110100110111: color_data = Z;
		19'b1001111110100111000: color_data = Z;
		19'b1001111110100111001: color_data = Z;
		19'b1001111110100111010: color_data = Z;
		19'b1001111110100111011: color_data = Z;
		19'b1001111110100111100: color_data = Z;
		19'b1001111110101000001: color_data = Z;
		19'b1001111110101000010: color_data = Z;
		19'b1001111110101000011: color_data = Z;
		19'b1001111110101000100: color_data = Z;
		19'b1001111110101000101: color_data = Z;
		19'b1001111110101000110: color_data = Z;
		19'b1001111110101000111: color_data = Z;
		19'b1001111110101010010: color_data = Z;
		19'b1001111110101010011: color_data = Z;
		19'b1001111110101010100: color_data = Z;
		19'b1001111110101010101: color_data = Z;
		19'b1001111110101010110: color_data = Z;
		19'b1001111110101010111: color_data = Z;
		19'b1001111110101100010: color_data = Z;
		19'b1001111110101100011: color_data = Z;
		19'b1001111110101100100: color_data = Z;
		19'b1001111110110101011: color_data = Z;
		19'b1001111110110101100: color_data = Z;
		19'b1001111110110101101: color_data = Z;
		19'b1001111110110101110: color_data = Z;
		19'b1001111110110101111: color_data = Z;
		19'b1001111110110110000: color_data = Z;
		19'b1001111110110110011: color_data = Z;
		19'b1001111110110110100: color_data = Z;
		19'b1001111110110110101: color_data = Z;
		19'b1001111110110110110: color_data = Z;
		19'b1001111110110111011: color_data = Z;
		19'b1010000000011000110: color_data = Z;
		19'b1010000000011010111: color_data = Z;
		19'b1010000000011011000: color_data = Z;
		19'b1010000000011011001: color_data = Z;
		19'b1010000000011011010: color_data = Z;
		19'b1010000000011011011: color_data = Z;
		19'b1010000000011011100: color_data = Z;
		19'b1010000000011011101: color_data = Z;
		19'b1010000000011011110: color_data = Z;
		19'b1010000000011011111: color_data = Z;
		19'b1010000000011100000: color_data = Z;
		19'b1010000000011100001: color_data = Z;
		19'b1010000000011100010: color_data = Z;
		19'b1010000000011100011: color_data = Z;
		19'b1010000000100110101: color_data = Z;
		19'b1010000000100110110: color_data = Z;
		19'b1010000000100110111: color_data = Z;
		19'b1010000000100111000: color_data = Z;
		19'b1010000000100111001: color_data = Z;
		19'b1010000000100111010: color_data = Z;
		19'b1010000000100111011: color_data = Z;
		19'b1010000000100111100: color_data = Z;
		19'b1010000000101000001: color_data = Z;
		19'b1010000000101000010: color_data = Z;
		19'b1010000000101000011: color_data = Z;
		19'b1010000000101000100: color_data = Z;
		19'b1010000000101010011: color_data = Z;
		19'b1010000000101010100: color_data = Z;
		19'b1010000000101010101: color_data = Z;
		19'b1010000000101010110: color_data = Z;
		19'b1010000000101100011: color_data = Z;
		19'b1010000000110101011: color_data = Z;
		19'b1010000000110101100: color_data = Z;
		19'b1010000000110101101: color_data = Z;
		19'b1010000000110101110: color_data = Z;
		19'b1010000000110101111: color_data = Z;
		19'b1010000000110110000: color_data = Z;
		19'b1010000000110110011: color_data = Z;
		19'b1010000000110110100: color_data = Z;
		19'b1010000000110110101: color_data = Z;
		19'b1010000010011010111: color_data = Z;
		19'b1010000010011011000: color_data = Z;
		19'b1010000010011011001: color_data = Z;
		19'b1010000010011011010: color_data = Z;
		19'b1010000010011011011: color_data = Z;
		19'b1010000010011011100: color_data = Z;
		19'b1010000010011011101: color_data = Z;
		19'b1010000010011011110: color_data = Z;
		19'b1010000010011011111: color_data = Z;
		19'b1010000010011100000: color_data = Z;
		19'b1010000010011100001: color_data = Z;
		19'b1010000010011100010: color_data = Z;
		19'b1010000010011100011: color_data = Z;
		19'b1010000010100110101: color_data = Z;
		19'b1010000010100110110: color_data = Z;
		19'b1010000010100110111: color_data = Z;
		19'b1010000010100111000: color_data = Z;
		19'b1010000010100111001: color_data = Z;
		19'b1010000010100111010: color_data = Z;
		19'b1010000010100111011: color_data = Z;
		19'b1010000010100111100: color_data = Z;
		19'b1010000010100111101: color_data = Z;
		19'b1010000010110101010: color_data = Z;
		19'b1010000010110101011: color_data = Z;
		19'b1010000010110101100: color_data = Z;
		19'b1010000010110101101: color_data = Z;
		19'b1010000010110101110: color_data = Z;
		19'b1010000010110101111: color_data = Z;
		19'b1010000010110110000: color_data = Z;
		19'b1010000010110110011: color_data = Z;
		19'b1010000010110110100: color_data = Z;
		19'b1010000010110110101: color_data = Z;
		19'b1010000100011000111: color_data = Z;
		19'b1010000100011011000: color_data = Z;
		19'b1010000100011011001: color_data = Z;
		19'b1010000100011011010: color_data = Z;
		19'b1010000100011011011: color_data = Z;
		19'b1010000100011011100: color_data = Z;
		19'b1010000100011011101: color_data = Z;
		19'b1010000100011011110: color_data = Z;
		19'b1010000100011011111: color_data = Z;
		19'b1010000100011100000: color_data = Z;
		19'b1010000100011100001: color_data = Z;
		19'b1010000100011100010: color_data = Z;
		19'b1010000100011100011: color_data = Z;
		19'b1010000100011100100: color_data = Z;
		19'b1010000100100110101: color_data = Z;
		19'b1010000100100110110: color_data = Z;
		19'b1010000100100110111: color_data = Z;
		19'b1010000100100111000: color_data = Z;
		19'b1010000100100111001: color_data = Z;
		19'b1010000100100111010: color_data = Z;
		19'b1010000100100111011: color_data = Z;
		19'b1010000100100111100: color_data = Z;
		19'b1010000100110101010: color_data = Z;
		19'b1010000100110101011: color_data = Z;
		19'b1010000100110101100: color_data = Z;
		19'b1010000100110101101: color_data = Z;
		19'b1010000100110101110: color_data = Z;
		19'b1010000100110101111: color_data = Z;
		19'b1010000100110110000: color_data = Z;
		19'b1010000100110110010: color_data = Z;
		19'b1010000100110110011: color_data = Z;
		19'b1010000100110110100: color_data = Z;
		19'b1010000100110110101: color_data = Z;
		19'b1010000110011011000: color_data = Z;
		19'b1010000110011011001: color_data = Z;
		19'b1010000110011011010: color_data = Z;
		19'b1010000110011011011: color_data = Z;
		19'b1010000110011011100: color_data = Z;
		19'b1010000110011011101: color_data = Z;
		19'b1010000110011011110: color_data = Z;
		19'b1010000110011011111: color_data = Z;
		19'b1010000110011100000: color_data = Z;
		19'b1010000110011100001: color_data = Z;
		19'b1010000110011100010: color_data = Z;
		19'b1010000110011100011: color_data = Z;
		19'b1010000110011100100: color_data = Z;
		19'b1010000110100110110: color_data = Z;
		19'b1010000110100110111: color_data = Z;
		19'b1010000110100111000: color_data = Z;
		19'b1010000110100111001: color_data = Z;
		19'b1010000110100111010: color_data = Z;
		19'b1010000110100111011: color_data = Z;
		19'b1010000110100111100: color_data = Z;
		19'b1010000110110101001: color_data = Z;
		19'b1010000110110101010: color_data = Z;
		19'b1010000110110101011: color_data = Z;
		19'b1010000110110101100: color_data = Z;
		19'b1010000110110101101: color_data = Z;
		19'b1010000110110101110: color_data = Z;
		19'b1010000110110101111: color_data = Z;
		19'b1010000110110110010: color_data = Z;
		19'b1010000110110110011: color_data = Z;
		19'b1010000110110110100: color_data = Z;
		19'b1010000110110110101: color_data = Z;
		19'b1010001000011001000: color_data = Z;
		19'b1010001000011011001: color_data = Z;
		19'b1010001000011011010: color_data = Z;
		19'b1010001000011011011: color_data = Z;
		19'b1010001000011011100: color_data = Z;
		19'b1010001000011011101: color_data = Z;
		19'b1010001000011011110: color_data = Z;
		19'b1010001000011011111: color_data = Z;
		19'b1010001000011100000: color_data = Z;
		19'b1010001000011100001: color_data = Z;
		19'b1010001000011100010: color_data = Z;
		19'b1010001000011100011: color_data = Z;
		19'b1010001000011100100: color_data = Z;
		19'b1010001000100110110: color_data = Z;
		19'b1010001000100110111: color_data = Z;
		19'b1010001000100111000: color_data = Z;
		19'b1010001000100111001: color_data = Z;
		19'b1010001000100111010: color_data = Z;
		19'b1010001000100111011: color_data = Z;
		19'b1010001000110101001: color_data = Z;
		19'b1010001000110101010: color_data = Z;
		19'b1010001000110101011: color_data = Z;
		19'b1010001000110101100: color_data = Z;
		19'b1010001000110101101: color_data = Z;
		19'b1010001000110101110: color_data = Z;
		19'b1010001000110101111: color_data = Z;
		19'b1010001000110110001: color_data = Z;
		19'b1010001000110110010: color_data = Z;
		19'b1010001000110110011: color_data = Z;
		19'b1010001000110110100: color_data = Z;
		19'b1010001000110110101: color_data = Z;
		19'b1010001010011001000: color_data = Z;
		19'b1010001010011011001: color_data = Z;
		19'b1010001010011011010: color_data = Z;
		19'b1010001010011011011: color_data = Z;
		19'b1010001010011011100: color_data = Z;
		19'b1010001010011011101: color_data = Z;
		19'b1010001010011011110: color_data = Z;
		19'b1010001010011011111: color_data = Z;
		19'b1010001010011100000: color_data = Z;
		19'b1010001010011100001: color_data = Z;
		19'b1010001010011100010: color_data = Z;
		19'b1010001010011100011: color_data = Z;
		19'b1010001010011100100: color_data = Z;
		19'b1010001010011100101: color_data = Z;
		19'b1010001010100111001: color_data = Z;
		19'b1010001010100111010: color_data = Z;
		19'b1010001010100111011: color_data = Z;
		19'b1010001010110101000: color_data = Z;
		19'b1010001010110101001: color_data = Z;
		19'b1010001010110101010: color_data = Z;
		19'b1010001010110101011: color_data = Z;
		19'b1010001010110101100: color_data = Z;
		19'b1010001010110101101: color_data = Z;
		19'b1010001010110101110: color_data = Z;
		19'b1010001010110101111: color_data = Z;
		19'b1010001010110110000: color_data = Z;
		19'b1010001010110110001: color_data = Z;
		19'b1010001010110110010: color_data = Z;
		19'b1010001010110110011: color_data = Z;
		19'b1010001010110110100: color_data = Z;
		19'b1010001010110110101: color_data = Z;
		19'b1010001100011001001: color_data = Z;
		19'b1010001100011011010: color_data = Z;
		19'b1010001100011011011: color_data = Z;
		19'b1010001100011011100: color_data = Z;
		19'b1010001100011011101: color_data = Z;
		19'b1010001100011011110: color_data = Z;
		19'b1010001100011011111: color_data = Z;
		19'b1010001100011100000: color_data = Z;
		19'b1010001100011100001: color_data = Z;
		19'b1010001100011100010: color_data = Z;
		19'b1010001100011100011: color_data = Z;
		19'b1010001100011100100: color_data = Z;
		19'b1010001100011100101: color_data = Z;
		19'b1010001100110101000: color_data = Z;
		19'b1010001100110101001: color_data = Z;
		19'b1010001100110101010: color_data = Z;
		19'b1010001100110101011: color_data = Z;
		19'b1010001100110101100: color_data = Z;
		19'b1010001100110101101: color_data = Z;
		19'b1010001100110101110: color_data = Z;
		19'b1010001100110101111: color_data = Z;
		19'b1010001100110110000: color_data = Z;
		19'b1010001100110110001: color_data = Z;
		19'b1010001100110110010: color_data = Z;
		19'b1010001100110110011: color_data = Z;
		19'b1010001100110110100: color_data = Z;
		19'b1010001110011001001: color_data = Z;
		19'b1010001110011001010: color_data = Z;
		19'b1010001110011011010: color_data = Z;
		19'b1010001110011011011: color_data = Z;
		19'b1010001110011011100: color_data = Z;
		19'b1010001110011011101: color_data = Z;
		19'b1010001110011011110: color_data = Z;
		19'b1010001110011011111: color_data = Z;
		19'b1010001110011100000: color_data = Z;
		19'b1010001110011100001: color_data = Z;
		19'b1010001110011100010: color_data = Z;
		19'b1010001110011100011: color_data = Z;
		19'b1010001110011100100: color_data = Z;
		19'b1010001110011100101: color_data = Z;
		19'b1010001110011100110: color_data = Z;
		19'b1010001110110100111: color_data = Z;
		19'b1010001110110101000: color_data = Z;
		19'b1010001110110101010: color_data = Z;
		19'b1010001110110101011: color_data = Z;
		19'b1010001110110101100: color_data = Z;
		19'b1010001110110101101: color_data = Z;
		19'b1010001110110101110: color_data = Z;
		19'b1010001110110101111: color_data = Z;
		19'b1010001110110110000: color_data = Z;
		19'b1010001110110110001: color_data = Z;
		19'b1010001110110110010: color_data = Z;
		19'b1010001110110110011: color_data = Z;
		19'b1010001110110110100: color_data = Z;
		19'b1010010000011001010: color_data = Z;
		19'b1010010000011001011: color_data = Z;
		19'b1010010000011011010: color_data = Z;
		19'b1010010000011011011: color_data = Z;
		19'b1010010000011011100: color_data = Z;
		19'b1010010000011011101: color_data = Z;
		19'b1010010000011011110: color_data = Z;
		19'b1010010000011011111: color_data = Z;
		19'b1010010000011100000: color_data = Z;
		19'b1010010000011100001: color_data = Z;
		19'b1010010000011100010: color_data = Z;
		19'b1010010000011100011: color_data = Z;
		19'b1010010000011100100: color_data = Z;
		19'b1010010000011100101: color_data = Z;
		19'b1010010000011100110: color_data = Z;
		19'b1010010000110100111: color_data = Z;
		19'b1010010000110101000: color_data = Z;
		19'b1010010000110101010: color_data = Z;
		19'b1010010000110101011: color_data = Z;
		19'b1010010000110101100: color_data = Z;
		19'b1010010000110101101: color_data = Z;
		19'b1010010000110101110: color_data = Z;
		19'b1010010000110101111: color_data = Z;
		19'b1010010000110110000: color_data = Z;
		19'b1010010000110110001: color_data = Z;
		19'b1010010000110110010: color_data = Z;
		19'b1010010000110110011: color_data = Z;
		19'b1010010000110110100: color_data = Z;
		19'b1010010010011001010: color_data = Z;
		19'b1010010010011001011: color_data = Z;
		19'b1010010010011011011: color_data = Z;
		19'b1010010010011011100: color_data = Z;
		19'b1010010010011011101: color_data = Z;
		19'b1010010010011011110: color_data = Z;
		19'b1010010010011011111: color_data = Z;
		19'b1010010010011100000: color_data = Z;
		19'b1010010010011100001: color_data = Z;
		19'b1010010010011100010: color_data = Z;
		19'b1010010010011100011: color_data = Z;
		19'b1010010010011100100: color_data = Z;
		19'b1010010010011100101: color_data = Z;
		19'b1010010010011100110: color_data = Z;
		19'b1010010010110100110: color_data = Z;
		19'b1010010010110100111: color_data = Z;
		19'b1010010010110101000: color_data = Z;
		19'b1010010010110101001: color_data = Z;
		19'b1010010010110101010: color_data = Z;
		19'b1010010010110101011: color_data = Z;
		19'b1010010010110101100: color_data = Z;
		19'b1010010010110101101: color_data = Z;
		19'b1010010010110101110: color_data = Z;
		19'b1010010010110101111: color_data = Z;
		19'b1010010010110110000: color_data = Z;
		19'b1010010010110110001: color_data = Z;
		19'b1010010010110110010: color_data = Z;
		19'b1010010010110110011: color_data = Z;
		19'b1010010010110110100: color_data = Z;
		19'b1010010100011001010: color_data = Z;
		19'b1010010100011001011: color_data = Z;
		19'b1010010100011001100: color_data = Z;
		19'b1010010100011011011: color_data = Z;
		19'b1010010100011011100: color_data = Z;
		19'b1010010100011011101: color_data = Z;
		19'b1010010100011011110: color_data = Z;
		19'b1010010100011011111: color_data = Z;
		19'b1010010100011100000: color_data = Z;
		19'b1010010100011100001: color_data = Z;
		19'b1010010100011100010: color_data = Z;
		19'b1010010100011100011: color_data = Z;
		19'b1010010100011100100: color_data = Z;
		19'b1010010100011100101: color_data = Z;
		19'b1010010100011100110: color_data = Z;
		19'b1010010100011100111: color_data = Z;
		19'b1010010100110001101: color_data = Z;
		19'b1010010100110001110: color_data = Z;
		19'b1010010100110100101: color_data = Z;
		19'b1010010100110100110: color_data = Z;
		19'b1010010100110100111: color_data = Z;
		19'b1010010100110101000: color_data = Z;
		19'b1010010100110101001: color_data = Z;
		19'b1010010100110101010: color_data = Z;
		19'b1010010100110101011: color_data = Z;
		19'b1010010100110101100: color_data = Z;
		19'b1010010100110101101: color_data = Z;
		19'b1010010100110101110: color_data = Z;
		19'b1010010100110101111: color_data = Z;
		19'b1010010100110110000: color_data = Z;
		19'b1010010100110110001: color_data = Z;
		19'b1010010110011001011: color_data = Z;
		19'b1010010110011001100: color_data = Z;
		19'b1010010110011011101: color_data = Z;
		19'b1010010110011011110: color_data = Z;
		19'b1010010110011011111: color_data = Z;
		19'b1010010110011100000: color_data = Z;
		19'b1010010110011100001: color_data = Z;
		19'b1010010110011100010: color_data = Z;
		19'b1010010110011100011: color_data = Z;
		19'b1010010110011100100: color_data = Z;
		19'b1010010110011100101: color_data = Z;
		19'b1010010110011100110: color_data = Z;
		19'b1010010110011100111: color_data = Z;
		19'b1010010110110001100: color_data = Z;
		19'b1010010110110001101: color_data = Z;
		19'b1010010110110001110: color_data = Z;
		19'b1010010110110001111: color_data = Z;
		19'b1010010110110100101: color_data = Z;
		19'b1010010110110100110: color_data = Z;
		19'b1010010110110100111: color_data = Z;
		19'b1010010110110101000: color_data = Z;
		19'b1010010110110101001: color_data = Z;
		19'b1010010110110101010: color_data = Z;
		19'b1010010110110101011: color_data = Z;
		19'b1010010110110101100: color_data = Z;
		19'b1010010110110101101: color_data = Z;
		19'b1010010110110101110: color_data = Z;
		19'b1010010110110110000: color_data = Z;
		19'b1010010110110110001: color_data = Z;
		19'b1010011000011001011: color_data = Z;
		19'b1010011000011001100: color_data = Z;
		19'b1010011000011001101: color_data = Z;
		19'b1010011000011011101: color_data = Z;
		19'b1010011000011011110: color_data = Z;
		19'b1010011000011011111: color_data = Z;
		19'b1010011000011100000: color_data = Z;
		19'b1010011000011100001: color_data = Z;
		19'b1010011000011100010: color_data = Z;
		19'b1010011000011100011: color_data = Z;
		19'b1010011000011100100: color_data = Z;
		19'b1010011000011100101: color_data = Z;
		19'b1010011000011100110: color_data = Z;
		19'b1010011000011100111: color_data = Z;
		19'b1010011000011101000: color_data = Z;
		19'b1010011000011101001: color_data = Z;
		19'b1010011000011101010: color_data = Z;
		19'b1010011000011101011: color_data = Z;
		19'b1010011000110001001: color_data = Z;
		19'b1010011000110001010: color_data = Z;
		19'b1010011000110001011: color_data = Z;
		19'b1010011000110001100: color_data = Z;
		19'b1010011000110001101: color_data = Z;
		19'b1010011000110001110: color_data = Z;
		19'b1010011000110001111: color_data = Z;
		19'b1010011000110100100: color_data = Z;
		19'b1010011000110100101: color_data = Z;
		19'b1010011000110100110: color_data = Z;
		19'b1010011000110100111: color_data = Z;
		19'b1010011000110101000: color_data = Z;
		19'b1010011000110101001: color_data = Z;
		19'b1010011000110101010: color_data = Z;
		19'b1010011000110101011: color_data = Z;
		19'b1010011000110101100: color_data = Z;
		19'b1010011000110101101: color_data = Z;
		19'b1010011000110101110: color_data = Z;
		19'b1010011000110110000: color_data = Z;
		19'b1010011010011001100: color_data = Z;
		19'b1010011010011001101: color_data = Z;
		19'b1010011010011001110: color_data = Z;
		19'b1010011010011011101: color_data = Z;
		19'b1010011010011011110: color_data = Z;
		19'b1010011010011011111: color_data = Z;
		19'b1010011010011100000: color_data = Z;
		19'b1010011010011100001: color_data = Z;
		19'b1010011010011100010: color_data = Z;
		19'b1010011010011100011: color_data = Z;
		19'b1010011010011100100: color_data = Z;
		19'b1010011010011100101: color_data = Z;
		19'b1010011010011100110: color_data = Z;
		19'b1010011010011100111: color_data = Z;
		19'b1010011010011101000: color_data = Z;
		19'b1010011010011101001: color_data = Z;
		19'b1010011010011101010: color_data = Z;
		19'b1010011010011101011: color_data = Z;
		19'b1010011010011101100: color_data = Z;
		19'b1010011010011101101: color_data = Z;
		19'b1010011010101111011: color_data = Z;
		19'b1010011010101111100: color_data = Z;
		19'b1010011010110001000: color_data = Z;
		19'b1010011010110001001: color_data = Z;
		19'b1010011010110001010: color_data = Z;
		19'b1010011010110001011: color_data = Z;
		19'b1010011010110001100: color_data = Z;
		19'b1010011010110001101: color_data = Z;
		19'b1010011010110001110: color_data = Z;
		19'b1010011010110001111: color_data = Z;
		19'b1010011010110100100: color_data = Z;
		19'b1010011010110100101: color_data = Z;
		19'b1010011010110100110: color_data = Z;
		19'b1010011010110100111: color_data = Z;
		19'b1010011010110101000: color_data = Z;
		19'b1010011010110101001: color_data = Z;
		19'b1010011010110101010: color_data = Z;
		19'b1010011010110101011: color_data = Z;
		19'b1010011010110101100: color_data = Z;
		19'b1010011010110101101: color_data = Z;
		19'b1010011010110101110: color_data = Z;
		19'b1010011010110101111: color_data = Z;
		19'b1010011100011001101: color_data = Z;
		19'b1010011100011001110: color_data = Z;
		19'b1010011100011001111: color_data = Z;
		19'b1010011100011011110: color_data = Z;
		19'b1010011100011011111: color_data = Z;
		19'b1010011100011100000: color_data = Z;
		19'b1010011100011100001: color_data = Z;
		19'b1010011100011100010: color_data = Z;
		19'b1010011100011100011: color_data = Z;
		19'b1010011100011100100: color_data = Z;
		19'b1010011100011100101: color_data = Z;
		19'b1010011100011100110: color_data = Z;
		19'b1010011100011100111: color_data = Z;
		19'b1010011100011101000: color_data = Z;
		19'b1010011100011101001: color_data = Z;
		19'b1010011100011101010: color_data = Z;
		19'b1010011100011101011: color_data = Z;
		19'b1010011100011101100: color_data = Z;
		19'b1010011100011101101: color_data = Z;
		19'b1010011100011101110: color_data = Z;
		19'b1010011100101111010: color_data = Z;
		19'b1010011100101111011: color_data = Z;
		19'b1010011100101111100: color_data = Z;
		19'b1010011100110001000: color_data = Z;
		19'b1010011100110001001: color_data = Z;
		19'b1010011100110001010: color_data = Z;
		19'b1010011100110001011: color_data = Z;
		19'b1010011100110001100: color_data = Z;
		19'b1010011100110001101: color_data = Z;
		19'b1010011100110001110: color_data = Z;
		19'b1010011100110001111: color_data = Z;
		19'b1010011100110100011: color_data = Z;
		19'b1010011100110100100: color_data = Z;
		19'b1010011100110100101: color_data = Z;
		19'b1010011100110100110: color_data = Z;
		19'b1010011100110100111: color_data = Z;
		19'b1010011100110101000: color_data = Z;
		19'b1010011100110101001: color_data = Z;
		19'b1010011100110101010: color_data = Z;
		19'b1010011100110101011: color_data = Z;
		19'b1010011100110101100: color_data = Z;
		19'b1010011100110101101: color_data = Z;
		19'b1010011100110101110: color_data = Z;
		19'b1010011100110101111: color_data = Z;
		19'b1010011110011001101: color_data = Z;
		19'b1010011110011001110: color_data = Z;
		19'b1010011110011001111: color_data = Z;
		19'b1010011110011011110: color_data = Z;
		19'b1010011110011011111: color_data = Z;
		19'b1010011110011100000: color_data = Z;
		19'b1010011110011100001: color_data = Z;
		19'b1010011110011100010: color_data = Z;
		19'b1010011110011100011: color_data = Z;
		19'b1010011110011100100: color_data = Z;
		19'b1010011110011100101: color_data = Z;
		19'b1010011110011100110: color_data = Z;
		19'b1010011110011100111: color_data = Z;
		19'b1010011110011101000: color_data = Z;
		19'b1010011110011101001: color_data = Z;
		19'b1010011110011101010: color_data = Z;
		19'b1010011110011101011: color_data = Z;
		19'b1010011110011101100: color_data = Z;
		19'b1010011110011101101: color_data = Z;
		19'b1010011110011101110: color_data = Z;
		19'b1010011110011101111: color_data = Z;
		19'b1010011110101111010: color_data = Z;
		19'b1010011110101111011: color_data = Z;
		19'b1010011110101111100: color_data = Z;
		19'b1010011110110000111: color_data = Z;
		19'b1010011110110001000: color_data = Z;
		19'b1010011110110001001: color_data = Z;
		19'b1010011110110001010: color_data = Z;
		19'b1010011110110001011: color_data = Z;
		19'b1010011110110001100: color_data = Z;
		19'b1010011110110001101: color_data = Z;
		19'b1010011110110001110: color_data = Z;
		19'b1010011110110001111: color_data = Z;
		19'b1010011110110100011: color_data = Z;
		19'b1010011110110100100: color_data = Z;
		19'b1010011110110100101: color_data = Z;
		19'b1010011110110100110: color_data = Z;
		19'b1010011110110100111: color_data = Z;
		19'b1010011110110101000: color_data = Z;
		19'b1010011110110101001: color_data = Z;
		19'b1010011110110101010: color_data = Z;
		19'b1010011110110101011: color_data = Z;
		19'b1010011110110101100: color_data = Z;
		19'b1010011110110101101: color_data = Z;
		19'b1010011110110101110: color_data = Z;
		19'b1010011110110101111: color_data = Z;
		19'b1010100000011001110: color_data = Z;
		19'b1010100000011001111: color_data = Z;
		19'b1010100000011010000: color_data = Z;
		19'b1010100000011011111: color_data = Z;
		19'b1010100000011100000: color_data = Z;
		19'b1010100000011100001: color_data = Z;
		19'b1010100000011100010: color_data = Z;
		19'b1010100000011100011: color_data = Z;
		19'b1010100000011100100: color_data = Z;
		19'b1010100000011100101: color_data = Z;
		19'b1010100000011100110: color_data = Z;
		19'b1010100000011100111: color_data = Z;
		19'b1010100000011101000: color_data = Z;
		19'b1010100000011101001: color_data = Z;
		19'b1010100000011101010: color_data = Z;
		19'b1010100000011101011: color_data = Z;
		19'b1010100000011101100: color_data = Z;
		19'b1010100000011101101: color_data = Z;
		19'b1010100000011101110: color_data = Z;
		19'b1010100000011101111: color_data = Z;
		19'b1010100000011110000: color_data = Z;
		19'b1010100000011110001: color_data = Z;
		19'b1010100000101110111: color_data = Z;
		19'b1010100000101111000: color_data = Z;
		19'b1010100000101111001: color_data = Z;
		19'b1010100000101111010: color_data = Z;
		19'b1010100000101111011: color_data = Z;
		19'b1010100000101111100: color_data = Z;
		19'b1010100000110000111: color_data = Z;
		19'b1010100000110001000: color_data = Z;
		19'b1010100000110001001: color_data = Z;
		19'b1010100000110001010: color_data = Z;
		19'b1010100000110001011: color_data = Z;
		19'b1010100000110001100: color_data = Z;
		19'b1010100000110001101: color_data = Z;
		19'b1010100000110001110: color_data = Z;
		19'b1010100000110001111: color_data = Z;
		19'b1010100000110100010: color_data = Z;
		19'b1010100000110100011: color_data = Z;
		19'b1010100000110100100: color_data = Z;
		19'b1010100000110100101: color_data = Z;
		19'b1010100000110100110: color_data = Z;
		19'b1010100000110100111: color_data = Z;
		19'b1010100000110101000: color_data = Z;
		19'b1010100000110101001: color_data = Z;
		19'b1010100000110101010: color_data = Z;
		19'b1010100000110101011: color_data = Z;
		19'b1010100000110101100: color_data = Z;
		19'b1010100000110101101: color_data = Z;
		19'b1010100000110101110: color_data = Z;
		19'b1010100000110101111: color_data = Z;
		19'b1010100010011001111: color_data = Z;
		19'b1010100010011010000: color_data = Z;
		19'b1010100010011010001: color_data = Z;
		19'b1010100010011011111: color_data = Z;
		19'b1010100010011100000: color_data = Z;
		19'b1010100010011100001: color_data = Z;
		19'b1010100010011100010: color_data = Z;
		19'b1010100010011100011: color_data = Z;
		19'b1010100010011100100: color_data = Z;
		19'b1010100010011100101: color_data = Z;
		19'b1010100010011100110: color_data = Z;
		19'b1010100010011100111: color_data = Z;
		19'b1010100010011101000: color_data = Z;
		19'b1010100010011101001: color_data = Z;
		19'b1010100010011101010: color_data = Z;
		19'b1010100010011101011: color_data = Z;
		19'b1010100010011101100: color_data = Z;
		19'b1010100010011101101: color_data = Z;
		19'b1010100010011101110: color_data = Z;
		19'b1010100010011101111: color_data = Z;
		19'b1010100010011110000: color_data = Z;
		19'b1010100010011110001: color_data = Z;
		19'b1010100010011110010: color_data = Z;
		19'b1010100010101110110: color_data = Z;
		19'b1010100010101110111: color_data = Z;
		19'b1010100010101111000: color_data = Z;
		19'b1010100010101111001: color_data = Z;
		19'b1010100010101111010: color_data = Z;
		19'b1010100010101111011: color_data = Z;
		19'b1010100010101111100: color_data = Z;
		19'b1010100010110000111: color_data = Z;
		19'b1010100010110001000: color_data = Z;
		19'b1010100010110001001: color_data = Z;
		19'b1010100010110001010: color_data = Z;
		19'b1010100010110001011: color_data = Z;
		19'b1010100010110001100: color_data = Z;
		19'b1010100010110001101: color_data = Z;
		19'b1010100010110001110: color_data = Z;
		19'b1010100010110001111: color_data = Z;
		19'b1010100010110100010: color_data = Z;
		19'b1010100010110100011: color_data = Z;
		19'b1010100010110100100: color_data = Z;
		19'b1010100010110100101: color_data = Z;
		19'b1010100010110100110: color_data = Z;
		19'b1010100010110100111: color_data = Z;
		19'b1010100010110101000: color_data = Z;
		19'b1010100010110101001: color_data = Z;
		19'b1010100010110101010: color_data = Z;
		19'b1010100010110101011: color_data = Z;
		19'b1010100010110101100: color_data = Z;
		19'b1010100010110101101: color_data = Z;
		19'b1010100100011010000: color_data = Z;
		19'b1010100100011010001: color_data = Z;
		19'b1010100100011010010: color_data = Z;
		19'b1010100100011100000: color_data = Z;
		19'b1010100100011100001: color_data = Z;
		19'b1010100100011100010: color_data = Z;
		19'b1010100100011100011: color_data = Z;
		19'b1010100100011100100: color_data = Z;
		19'b1010100100011100101: color_data = Z;
		19'b1010100100011100110: color_data = Z;
		19'b1010100100011100111: color_data = Z;
		19'b1010100100011101000: color_data = Z;
		19'b1010100100011101001: color_data = Z;
		19'b1010100100011101010: color_data = Z;
		19'b1010100100011101011: color_data = Z;
		19'b1010100100011101100: color_data = Z;
		19'b1010100100011101101: color_data = Z;
		19'b1010100100011101110: color_data = Z;
		19'b1010100100011101111: color_data = Z;
		19'b1010100100011110000: color_data = Z;
		19'b1010100100011110001: color_data = Z;
		19'b1010100100011110010: color_data = Z;
		19'b1010100100011110011: color_data = Z;
		19'b1010100100011110100: color_data = Z;
		19'b1010100100101110101: color_data = Z;
		19'b1010100100101110110: color_data = Z;
		19'b1010100100101110111: color_data = Z;
		19'b1010100100101111000: color_data = Z;
		19'b1010100100101111001: color_data = Z;
		19'b1010100100101111010: color_data = Z;
		19'b1010100100101111011: color_data = Z;
		19'b1010100100101111100: color_data = Z;
		19'b1010100100101111101: color_data = Z;
		19'b1010100100110000111: color_data = Z;
		19'b1010100100110001000: color_data = Z;
		19'b1010100100110001001: color_data = Z;
		19'b1010100100110001011: color_data = Z;
		19'b1010100100110001100: color_data = Z;
		19'b1010100100110001101: color_data = Z;
		19'b1010100100110001110: color_data = Z;
		19'b1010100100110001111: color_data = Z;
		19'b1010100100110100010: color_data = Z;
		19'b1010100100110100011: color_data = Z;
		19'b1010100100110100100: color_data = Z;
		19'b1010100100110100101: color_data = Z;
		19'b1010100100110100110: color_data = Z;
		19'b1010100100110100111: color_data = Z;
		19'b1010100100110101000: color_data = Z;
		19'b1010100100110101001: color_data = Z;
		19'b1010100100110101010: color_data = Z;
		19'b1010100100110101011: color_data = Z;
		19'b1010100100110101100: color_data = Z;
		19'b1010100110011010001: color_data = Z;
		19'b1010100110011010010: color_data = Z;
		19'b1010100110011010011: color_data = Z;
		19'b1010100110011100001: color_data = Z;
		19'b1010100110011100010: color_data = Z;
		19'b1010100110011100011: color_data = Z;
		19'b1010100110011100100: color_data = Z;
		19'b1010100110011100101: color_data = Z;
		19'b1010100110011100110: color_data = Z;
		19'b1010100110011100111: color_data = Z;
		19'b1010100110011101000: color_data = Z;
		19'b1010100110011101001: color_data = Z;
		19'b1010100110011101010: color_data = Z;
		19'b1010100110011101011: color_data = Z;
		19'b1010100110011101100: color_data = Z;
		19'b1010100110011101101: color_data = Z;
		19'b1010100110011101110: color_data = Z;
		19'b1010100110011101111: color_data = Z;
		19'b1010100110011110000: color_data = Z;
		19'b1010100110011110001: color_data = Z;
		19'b1010100110011110010: color_data = Z;
		19'b1010100110011110011: color_data = Z;
		19'b1010100110011110100: color_data = Z;
		19'b1010100110011110101: color_data = Z;
		19'b1010100110011110110: color_data = Z;
		19'b1010100110101110101: color_data = Z;
		19'b1010100110101110110: color_data = Z;
		19'b1010100110101110111: color_data = Z;
		19'b1010100110101111000: color_data = Z;
		19'b1010100110101111001: color_data = Z;
		19'b1010100110101111010: color_data = Z;
		19'b1010100110101111011: color_data = Z;
		19'b1010100110101111100: color_data = Z;
		19'b1010100110101111101: color_data = Z;
		19'b1010100110110000110: color_data = Z;
		19'b1010100110110000111: color_data = Z;
		19'b1010100110110001000: color_data = Z;
		19'b1010100110110001001: color_data = Z;
		19'b1010100110110001100: color_data = Z;
		19'b1010100110110001101: color_data = Z;
		19'b1010100110110001110: color_data = Z;
		19'b1010100110110001111: color_data = Z;
		19'b1010100110110100001: color_data = Z;
		19'b1010100110110100010: color_data = Z;
		19'b1010100110110100011: color_data = Z;
		19'b1010100110110100100: color_data = Z;
		19'b1010100110110100101: color_data = Z;
		19'b1010100110110100110: color_data = Z;
		19'b1010100110110100111: color_data = Z;
		19'b1010100110110101000: color_data = Z;
		19'b1010100110110101001: color_data = Z;
		19'b1010100110110101010: color_data = Z;
		19'b1010100110110101011: color_data = Z;
		19'b1010101000011010011: color_data = Z;
		19'b1010101000011010100: color_data = Z;
		19'b1010101000011100010: color_data = Z;
		19'b1010101000011100011: color_data = Z;
		19'b1010101000011100100: color_data = Z;
		19'b1010101000011100101: color_data = Z;
		19'b1010101000011100110: color_data = Z;
		19'b1010101000011100111: color_data = Z;
		19'b1010101000011101000: color_data = Z;
		19'b1010101000011101001: color_data = Z;
		19'b1010101000011101010: color_data = Z;
		19'b1010101000011101011: color_data = Z;
		19'b1010101000011101100: color_data = Z;
		19'b1010101000011101101: color_data = Z;
		19'b1010101000011101110: color_data = Z;
		19'b1010101000011101111: color_data = Z;
		19'b1010101000011110000: color_data = Z;
		19'b1010101000011110001: color_data = Z;
		19'b1010101000011110010: color_data = Z;
		19'b1010101000011110011: color_data = Z;
		19'b1010101000011110100: color_data = Z;
		19'b1010101000011110101: color_data = Z;
		19'b1010101000011110110: color_data = Z;
		19'b1010101000011110111: color_data = Z;
		19'b1010101000101110101: color_data = Z;
		19'b1010101000101110110: color_data = Z;
		19'b1010101000101110111: color_data = Z;
		19'b1010101000101111000: color_data = Z;
		19'b1010101000101111001: color_data = Z;
		19'b1010101000101111010: color_data = Z;
		19'b1010101000101111011: color_data = Z;
		19'b1010101000101111100: color_data = Z;
		19'b1010101000101111101: color_data = Z;
		19'b1010101000110000110: color_data = Z;
		19'b1010101000110000111: color_data = Z;
		19'b1010101000110001000: color_data = Z;
		19'b1010101000110001001: color_data = Z;
		19'b1010101000110001100: color_data = Z;
		19'b1010101000110001101: color_data = Z;
		19'b1010101000110001110: color_data = Z;
		19'b1010101000110001111: color_data = Z;
		19'b1010101000110100001: color_data = Z;
		19'b1010101000110100010: color_data = Z;
		19'b1010101000110100011: color_data = Z;
		19'b1010101000110100100: color_data = Z;
		19'b1010101000110100101: color_data = Z;
		19'b1010101000110100110: color_data = Z;
		19'b1010101000110100111: color_data = Z;
		19'b1010101000110101000: color_data = Z;
		19'b1010101000110101001: color_data = Z;
		19'b1010101000110101010: color_data = Z;
		19'b1010101000110101011: color_data = Z;
		19'b1010101010011010011: color_data = Z;
		19'b1010101010011010100: color_data = Z;
		19'b1010101010011010101: color_data = Z;
		19'b1010101010011100010: color_data = Z;
		19'b1010101010011100011: color_data = Z;
		19'b1010101010011100100: color_data = Z;
		19'b1010101010011100101: color_data = Z;
		19'b1010101010011100110: color_data = Z;
		19'b1010101010011100111: color_data = Z;
		19'b1010101010011101000: color_data = Z;
		19'b1010101010011101001: color_data = Z;
		19'b1010101010011101010: color_data = Z;
		19'b1010101010011101011: color_data = Z;
		19'b1010101010011101100: color_data = Z;
		19'b1010101010011101101: color_data = Z;
		19'b1010101010011101110: color_data = Z;
		19'b1010101010011101111: color_data = Z;
		19'b1010101010011110000: color_data = Z;
		19'b1010101010011110001: color_data = Z;
		19'b1010101010011110010: color_data = Z;
		19'b1010101010011110011: color_data = Z;
		19'b1010101010011110100: color_data = Z;
		19'b1010101010011110101: color_data = Z;
		19'b1010101010011110110: color_data = Z;
		19'b1010101010011110111: color_data = Z;
		19'b1010101010011111000: color_data = Z;
		19'b1010101010011111001: color_data = Z;
		19'b1010101010101110101: color_data = Z;
		19'b1010101010101110110: color_data = Z;
		19'b1010101010101110111: color_data = Z;
		19'b1010101010101111000: color_data = Z;
		19'b1010101010101111001: color_data = Z;
		19'b1010101010101111010: color_data = Z;
		19'b1010101010101111011: color_data = Z;
		19'b1010101010101111100: color_data = Z;
		19'b1010101010101111101: color_data = Z;
		19'b1010101010110000110: color_data = Z;
		19'b1010101010110000111: color_data = Z;
		19'b1010101010110001000: color_data = Z;
		19'b1010101010110001001: color_data = Z;
		19'b1010101010110001100: color_data = Z;
		19'b1010101010110001101: color_data = Z;
		19'b1010101010110001110: color_data = Z;
		19'b1010101010110001111: color_data = Z;
		19'b1010101010110010000: color_data = Z;
		19'b1010101010110100000: color_data = Z;
		19'b1010101010110100001: color_data = Z;
		19'b1010101010110100010: color_data = Z;
		19'b1010101010110100011: color_data = Z;
		19'b1010101010110100100: color_data = Z;
		19'b1010101010110100101: color_data = Z;
		19'b1010101010110100110: color_data = Z;
		19'b1010101010110100111: color_data = Z;
		19'b1010101010110101000: color_data = Z;
		19'b1010101010110101001: color_data = Z;
		19'b1010101010110101010: color_data = Z;
		19'b1010101100011010100: color_data = Z;
		19'b1010101100011010101: color_data = Z;
		19'b1010101100011010110: color_data = Z;
		19'b1010101100011100011: color_data = Z;
		19'b1010101100011100100: color_data = Z;
		19'b1010101100011100101: color_data = Z;
		19'b1010101100011100110: color_data = Z;
		19'b1010101100011100111: color_data = Z;
		19'b1010101100011101000: color_data = Z;
		19'b1010101100011101001: color_data = Z;
		19'b1010101100011101010: color_data = Z;
		19'b1010101100011101011: color_data = Z;
		19'b1010101100011101100: color_data = Z;
		19'b1010101100011101101: color_data = Z;
		19'b1010101100011101110: color_data = Z;
		19'b1010101100011101111: color_data = Z;
		19'b1010101100011110000: color_data = Z;
		19'b1010101100011110001: color_data = Z;
		19'b1010101100011110010: color_data = Z;
		19'b1010101100011110011: color_data = Z;
		19'b1010101100011110100: color_data = Z;
		19'b1010101100011110101: color_data = Z;
		19'b1010101100011110110: color_data = Z;
		19'b1010101100011110111: color_data = Z;
		19'b1010101100011111000: color_data = Z;
		19'b1010101100011111001: color_data = Z;
		19'b1010101100011111010: color_data = Z;
		19'b1010101100101110100: color_data = Z;
		19'b1010101100101110101: color_data = Z;
		19'b1010101100101110110: color_data = Z;
		19'b1010101100101110111: color_data = Z;
		19'b1010101100101111000: color_data = Z;
		19'b1010101100101111001: color_data = Z;
		19'b1010101100101111010: color_data = Z;
		19'b1010101100101111011: color_data = Z;
		19'b1010101100101111100: color_data = Z;
		19'b1010101100110000111: color_data = Z;
		19'b1010101100110001000: color_data = Z;
		19'b1010101100110001001: color_data = Z;
		19'b1010101100110001011: color_data = Z;
		19'b1010101100110001100: color_data = Z;
		19'b1010101100110001101: color_data = Z;
		19'b1010101100110001110: color_data = Z;
		19'b1010101100110001111: color_data = Z;
		19'b1010101100110100000: color_data = Z;
		19'b1010101100110100001: color_data = Z;
		19'b1010101100110100010: color_data = Z;
		19'b1010101100110100011: color_data = Z;
		19'b1010101100110100100: color_data = Z;
		19'b1010101100110100101: color_data = Z;
		19'b1010101100110100110: color_data = Z;
		19'b1010101100110100111: color_data = Z;
		19'b1010101100110101000: color_data = Z;
		19'b1010101100110101001: color_data = Z;
		19'b1010101100110101010: color_data = Z;
		19'b1010101110011010101: color_data = Z;
		19'b1010101110011010110: color_data = Z;
		19'b1010101110011010111: color_data = Z;
		19'b1010101110011100011: color_data = Z;
		19'b1010101110011100100: color_data = Z;
		19'b1010101110011100101: color_data = Z;
		19'b1010101110011100110: color_data = Z;
		19'b1010101110011100111: color_data = Z;
		19'b1010101110011101000: color_data = Z;
		19'b1010101110011101001: color_data = Z;
		19'b1010101110011101010: color_data = Z;
		19'b1010101110011101011: color_data = Z;
		19'b1010101110011101100: color_data = Z;
		19'b1010101110011101101: color_data = Z;
		19'b1010101110011101110: color_data = Z;
		19'b1010101110011101111: color_data = Z;
		19'b1010101110011110000: color_data = Z;
		19'b1010101110011110001: color_data = Z;
		19'b1010101110011110010: color_data = Z;
		19'b1010101110011110011: color_data = Z;
		19'b1010101110011110100: color_data = Z;
		19'b1010101110011110101: color_data = Z;
		19'b1010101110011110110: color_data = Z;
		19'b1010101110011110111: color_data = Z;
		19'b1010101110011111000: color_data = Z;
		19'b1010101110011111001: color_data = Z;
		19'b1010101110011111010: color_data = Z;
		19'b1010101110011111011: color_data = Z;
		19'b1010101110011111100: color_data = Z;
		19'b1010101110101110100: color_data = Z;
		19'b1010101110101110101: color_data = Z;
		19'b1010101110101110110: color_data = Z;
		19'b1010101110101110111: color_data = Z;
		19'b1010101110101111000: color_data = Z;
		19'b1010101110101111001: color_data = Z;
		19'b1010101110101111010: color_data = Z;
		19'b1010101110101111011: color_data = Z;
		19'b1010101110101111100: color_data = Z;
		19'b1010101110110000111: color_data = Z;
		19'b1010101110110001000: color_data = Z;
		19'b1010101110110001001: color_data = Z;
		19'b1010101110110001010: color_data = Z;
		19'b1010101110110001100: color_data = Z;
		19'b1010101110110001101: color_data = Z;
		19'b1010101110110001110: color_data = Z;
		19'b1010101110110001111: color_data = Z;
		19'b1010101110110011111: color_data = Z;
		19'b1010101110110100000: color_data = Z;
		19'b1010101110110100001: color_data = Z;
		19'b1010101110110100010: color_data = Z;
		19'b1010101110110100011: color_data = Z;
		19'b1010101110110100100: color_data = Z;
		19'b1010101110110100101: color_data = Z;
		19'b1010101110110100110: color_data = Z;
		19'b1010101110110100111: color_data = Z;
		19'b1010101110110101000: color_data = Z;
		19'b1010101110110101001: color_data = Z;
		19'b1010110000011010110: color_data = Z;
		19'b1010110000011010111: color_data = Z;
		19'b1010110000011011000: color_data = Z;
		19'b1010110000011100100: color_data = Z;
		19'b1010110000011100101: color_data = Z;
		19'b1010110000011100110: color_data = Z;
		19'b1010110000011100111: color_data = Z;
		19'b1010110000011101000: color_data = Z;
		19'b1010110000011101001: color_data = Z;
		19'b1010110000011101010: color_data = Z;
		19'b1010110000011101011: color_data = Z;
		19'b1010110000011101100: color_data = Z;
		19'b1010110000011101101: color_data = Z;
		19'b1010110000011101110: color_data = Z;
		19'b1010110000011101111: color_data = Z;
		19'b1010110000011110000: color_data = Z;
		19'b1010110000011110001: color_data = Z;
		19'b1010110000011110010: color_data = Z;
		19'b1010110000011110011: color_data = Z;
		19'b1010110000011110100: color_data = Z;
		19'b1010110000011110101: color_data = Z;
		19'b1010110000011110110: color_data = Z;
		19'b1010110000011110111: color_data = Z;
		19'b1010110000011111000: color_data = Z;
		19'b1010110000011111001: color_data = Z;
		19'b1010110000011111010: color_data = Z;
		19'b1010110000011111011: color_data = Z;
		19'b1010110000011111100: color_data = Z;
		19'b1010110000011111101: color_data = Z;
		19'b1010110000101110100: color_data = Z;
		19'b1010110000101110101: color_data = Z;
		19'b1010110000101110110: color_data = Z;
		19'b1010110000101110111: color_data = Z;
		19'b1010110000101111000: color_data = Z;
		19'b1010110000101111001: color_data = Z;
		19'b1010110000101111010: color_data = Z;
		19'b1010110000101111011: color_data = Z;
		19'b1010110000101111100: color_data = Z;
		19'b1010110000110000111: color_data = Z;
		19'b1010110000110001000: color_data = Z;
		19'b1010110000110001001: color_data = Z;
		19'b1010110000110001010: color_data = Z;
		19'b1010110000110011111: color_data = Z;
		19'b1010110000110100000: color_data = Z;
		19'b1010110000110100001: color_data = Z;
		19'b1010110000110100010: color_data = Z;
		19'b1010110000110100011: color_data = Z;
		19'b1010110000110100100: color_data = Z;
		19'b1010110000110100101: color_data = Z;
		19'b1010110000110100110: color_data = Z;
		19'b1010110000110100111: color_data = Z;
		19'b1010110000110101000: color_data = Z;
		19'b1010110010011010111: color_data = Z;
		19'b1010110010011011000: color_data = Z;
		19'b1010110010011011001: color_data = Z;
		19'b1010110010011100100: color_data = Z;
		19'b1010110010011100101: color_data = Z;
		19'b1010110010011100110: color_data = Z;
		19'b1010110010011100111: color_data = Z;
		19'b1010110010011101000: color_data = Z;
		19'b1010110010011101001: color_data = Z;
		19'b1010110010011101010: color_data = Z;
		19'b1010110010011101011: color_data = Z;
		19'b1010110010011101100: color_data = Z;
		19'b1010110010011101101: color_data = Z;
		19'b1010110010011101110: color_data = Z;
		19'b1010110010011101111: color_data = Z;
		19'b1010110010011110000: color_data = Z;
		19'b1010110010011110001: color_data = Z;
		19'b1010110010011110010: color_data = Z;
		19'b1010110010011110011: color_data = Z;
		19'b1010110010011110100: color_data = Z;
		19'b1010110010011110101: color_data = Z;
		19'b1010110010011110110: color_data = Z;
		19'b1010110010011110111: color_data = Z;
		19'b1010110010011111000: color_data = Z;
		19'b1010110010011111001: color_data = Z;
		19'b1010110010011111010: color_data = Z;
		19'b1010110010011111011: color_data = Z;
		19'b1010110010011111100: color_data = Z;
		19'b1010110010011111101: color_data = Z;
		19'b1010110010011111110: color_data = Z;
		19'b1010110010101110100: color_data = Z;
		19'b1010110010101110101: color_data = Z;
		19'b1010110010101110110: color_data = Z;
		19'b1010110010101110111: color_data = Z;
		19'b1010110010101111000: color_data = Z;
		19'b1010110010101111001: color_data = Z;
		19'b1010110010101111010: color_data = Z;
		19'b1010110010110000111: color_data = Z;
		19'b1010110010110001000: color_data = Z;
		19'b1010110010110001001: color_data = Z;
		19'b1010110010110011111: color_data = Z;
		19'b1010110010110100000: color_data = Z;
		19'b1010110010110100001: color_data = Z;
		19'b1010110010110100010: color_data = Z;
		19'b1010110010110100011: color_data = Z;
		19'b1010110010110100100: color_data = Z;
		19'b1010110010110100101: color_data = Z;
		19'b1010110010110100110: color_data = Z;
		19'b1010110010110100111: color_data = Z;
		19'b1010110010110101000: color_data = Z;
		19'b1010110100011011000: color_data = Z;
		19'b1010110100011011001: color_data = Z;
		19'b1010110100011011010: color_data = Z;
		19'b1010110100011100100: color_data = Z;
		19'b1010110100011100101: color_data = Z;
		19'b1010110100011100110: color_data = Z;
		19'b1010110100011100111: color_data = Z;
		19'b1010110100011101000: color_data = Z;
		19'b1010110100011101001: color_data = Z;
		19'b1010110100011101010: color_data = Z;
		19'b1010110100011101011: color_data = Z;
		19'b1010110100011101100: color_data = Z;
		19'b1010110100011101101: color_data = Z;
		19'b1010110100011101110: color_data = Z;
		19'b1010110100011101111: color_data = Z;
		19'b1010110100011110000: color_data = Z;
		19'b1010110100011110001: color_data = Z;
		19'b1010110100011110010: color_data = Z;
		19'b1010110100011110011: color_data = Z;
		19'b1010110100011110100: color_data = Z;
		19'b1010110100011110101: color_data = Z;
		19'b1010110100011110110: color_data = Z;
		19'b1010110100011110111: color_data = Z;
		19'b1010110100011111000: color_data = Z;
		19'b1010110100011111001: color_data = Z;
		19'b1010110100011111010: color_data = Z;
		19'b1010110100011111011: color_data = Z;
		19'b1010110100011111100: color_data = Z;
		19'b1010110100011111101: color_data = Z;
		19'b1010110100011111110: color_data = Z;
		19'b1010110100011111111: color_data = Z;
		19'b1010110100100110101: color_data = Z;
		19'b1010110100100110110: color_data = Z;
		19'b1010110100100110111: color_data = Z;
		19'b1010110100100111000: color_data = Z;
		19'b1010110100101110011: color_data = Z;
		19'b1010110100101110100: color_data = Z;
		19'b1010110100101110101: color_data = Z;
		19'b1010110100101110110: color_data = Z;
		19'b1010110100101110111: color_data = Z;
		19'b1010110100101111000: color_data = Z;
		19'b1010110100101111001: color_data = Z;
		19'b1010110100110000111: color_data = Z;
		19'b1010110100110001000: color_data = Z;
		19'b1010110100110001001: color_data = Z;
		19'b1010110100110011110: color_data = Z;
		19'b1010110100110011111: color_data = Z;
		19'b1010110100110100000: color_data = Z;
		19'b1010110100110100001: color_data = Z;
		19'b1010110100110100010: color_data = Z;
		19'b1010110100110100011: color_data = Z;
		19'b1010110100110100100: color_data = Z;
		19'b1010110100110100101: color_data = Z;
		19'b1010110100110100110: color_data = Z;
		19'b1010110100110100111: color_data = Z;
		19'b1010110110011011001: color_data = Z;
		19'b1010110110011011010: color_data = Z;
		19'b1010110110011011011: color_data = Z;
		19'b1010110110011100101: color_data = Z;
		19'b1010110110011100110: color_data = Z;
		19'b1010110110011100111: color_data = Z;
		19'b1010110110011101000: color_data = Z;
		19'b1010110110011101001: color_data = Z;
		19'b1010110110011101010: color_data = Z;
		19'b1010110110011101011: color_data = Z;
		19'b1010110110011101100: color_data = Z;
		19'b1010110110011101101: color_data = Z;
		19'b1010110110011101110: color_data = Z;
		19'b1010110110011101111: color_data = Z;
		19'b1010110110011110000: color_data = Z;
		19'b1010110110011110001: color_data = Z;
		19'b1010110110011110010: color_data = Z;
		19'b1010110110011110011: color_data = Z;
		19'b1010110110011110100: color_data = Z;
		19'b1010110110011110101: color_data = Z;
		19'b1010110110011110110: color_data = Z;
		19'b1010110110011110111: color_data = Z;
		19'b1010110110011111000: color_data = Z;
		19'b1010110110011111001: color_data = Z;
		19'b1010110110011111010: color_data = Z;
		19'b1010110110011111011: color_data = Z;
		19'b1010110110011111100: color_data = Z;
		19'b1010110110011111101: color_data = Z;
		19'b1010110110011111110: color_data = Z;
		19'b1010110110011111111: color_data = Z;
		19'b1010110110100000000: color_data = Z;
		19'b1010110110100000001: color_data = Z;
		19'b1010110110100000010: color_data = Z;
		19'b1010110110100110100: color_data = Z;
		19'b1010110110100110101: color_data = Z;
		19'b1010110110100110110: color_data = Z;
		19'b1010110110100110111: color_data = Z;
		19'b1010110110100111000: color_data = Z;
		19'b1010110110100111001: color_data = Z;
		19'b1010110110101101011: color_data = Z;
		19'b1010110110101110011: color_data = Z;
		19'b1010110110101110100: color_data = Z;
		19'b1010110110101110101: color_data = Z;
		19'b1010110110101110110: color_data = Z;
		19'b1010110110101110111: color_data = Z;
		19'b1010110110101111000: color_data = Z;
		19'b1010110110110000111: color_data = Z;
		19'b1010110110110001000: color_data = Z;
		19'b1010110110110011110: color_data = Z;
		19'b1010110110110011111: color_data = Z;
		19'b1010110110110100000: color_data = Z;
		19'b1010110110110100001: color_data = Z;
		19'b1010110110110100010: color_data = Z;
		19'b1010110110110100011: color_data = Z;
		19'b1010110110110100100: color_data = Z;
		19'b1010110110110100101: color_data = Z;
		19'b1010110110110100110: color_data = Z;
		19'b1010110110110100111: color_data = Z;
		19'b1010111000011011010: color_data = Z;
		19'b1010111000011011011: color_data = Z;
		19'b1010111000011011100: color_data = Z;
		19'b1010111000011100101: color_data = Z;
		19'b1010111000011100110: color_data = Z;
		19'b1010111000011100111: color_data = Z;
		19'b1010111000011101000: color_data = Z;
		19'b1010111000011101001: color_data = Z;
		19'b1010111000011101010: color_data = Z;
		19'b1010111000011101011: color_data = Z;
		19'b1010111000011101100: color_data = Z;
		19'b1010111000011101101: color_data = Z;
		19'b1010111000011101110: color_data = Z;
		19'b1010111000011101111: color_data = Z;
		19'b1010111000011110000: color_data = Z;
		19'b1010111000011110001: color_data = Z;
		19'b1010111000011110010: color_data = Z;
		19'b1010111000011110011: color_data = Z;
		19'b1010111000011110100: color_data = Z;
		19'b1010111000011110101: color_data = Z;
		19'b1010111000011110110: color_data = Z;
		19'b1010111000011110111: color_data = Z;
		19'b1010111000011111000: color_data = Z;
		19'b1010111000011111001: color_data = Z;
		19'b1010111000011111010: color_data = Z;
		19'b1010111000011111011: color_data = Z;
		19'b1010111000011111100: color_data = Z;
		19'b1010111000011111101: color_data = Z;
		19'b1010111000011111110: color_data = Z;
		19'b1010111000011111111: color_data = Z;
		19'b1010111000100000000: color_data = Z;
		19'b1010111000100000001: color_data = Z;
		19'b1010111000100000010: color_data = Z;
		19'b1010111000100000011: color_data = Z;
		19'b1010111000100000100: color_data = Z;
		19'b1010111000100000101: color_data = Z;
		19'b1010111000100110100: color_data = Z;
		19'b1010111000100110101: color_data = Z;
		19'b1010111000100110110: color_data = Z;
		19'b1010111000100110111: color_data = Z;
		19'b1010111000100111000: color_data = Z;
		19'b1010111000100111001: color_data = Z;
		19'b1010111000100111010: color_data = Z;
		19'b1010111000101100110: color_data = Z;
		19'b1010111000101100111: color_data = Z;
		19'b1010111000101101000: color_data = Z;
		19'b1010111000101101001: color_data = Z;
		19'b1010111000101101010: color_data = Z;
		19'b1010111000101101011: color_data = Z;
		19'b1010111000101101100: color_data = Z;
		19'b1010111000101110011: color_data = Z;
		19'b1010111000101110100: color_data = Z;
		19'b1010111000101110101: color_data = Z;
		19'b1010111000101110110: color_data = Z;
		19'b1010111000101110111: color_data = Z;
		19'b1010111000101111000: color_data = Z;
		19'b1010111000110011101: color_data = Z;
		19'b1010111000110011110: color_data = Z;
		19'b1010111000110011111: color_data = Z;
		19'b1010111000110100000: color_data = Z;
		19'b1010111000110100001: color_data = Z;
		19'b1010111000110100010: color_data = Z;
		19'b1010111000110100011: color_data = Z;
		19'b1010111000110100100: color_data = Z;
		19'b1010111000110100101: color_data = Z;
		19'b1010111000110100110: color_data = Z;
		19'b1010111010011011011: color_data = Z;
		19'b1010111010011011100: color_data = Z;
		19'b1010111010011011111: color_data = Z;
		19'b1010111010011100000: color_data = Z;
		19'b1010111010011100101: color_data = Z;
		19'b1010111010011100110: color_data = Z;
		19'b1010111010011100111: color_data = Z;
		19'b1010111010011101000: color_data = Z;
		19'b1010111010011101001: color_data = Z;
		19'b1010111010011101010: color_data = Z;
		19'b1010111010011101011: color_data = Z;
		19'b1010111010011101100: color_data = Z;
		19'b1010111010011101101: color_data = Z;
		19'b1010111010011101110: color_data = Z;
		19'b1010111010011101111: color_data = Z;
		19'b1010111010011110000: color_data = Z;
		19'b1010111010011110001: color_data = Z;
		19'b1010111010011110010: color_data = Z;
		19'b1010111010011110011: color_data = Z;
		19'b1010111010011110100: color_data = Z;
		19'b1010111010011110101: color_data = Z;
		19'b1010111010011110110: color_data = Z;
		19'b1010111010011110111: color_data = Z;
		19'b1010111010011111000: color_data = Z;
		19'b1010111010011111001: color_data = Z;
		19'b1010111010011111010: color_data = Z;
		19'b1010111010011111011: color_data = Z;
		19'b1010111010011111100: color_data = Z;
		19'b1010111010011111101: color_data = Z;
		19'b1010111010011111110: color_data = Z;
		19'b1010111010011111111: color_data = Z;
		19'b1010111010100000000: color_data = Z;
		19'b1010111010100000001: color_data = Z;
		19'b1010111010100000010: color_data = Z;
		19'b1010111010100000011: color_data = Z;
		19'b1010111010100000100: color_data = Z;
		19'b1010111010100000101: color_data = Z;
		19'b1010111010100000110: color_data = Z;
		19'b1010111010100110100: color_data = Z;
		19'b1010111010100110101: color_data = Z;
		19'b1010111010100110110: color_data = Z;
		19'b1010111010100110111: color_data = Z;
		19'b1010111010100111000: color_data = Z;
		19'b1010111010100111001: color_data = Z;
		19'b1010111010100111010: color_data = Z;
		19'b1010111010100111011: color_data = Z;
		19'b1010111010101011011: color_data = Z;
		19'b1010111010101100101: color_data = Z;
		19'b1010111010101100110: color_data = Z;
		19'b1010111010101100111: color_data = Z;
		19'b1010111010101101000: color_data = Z;
		19'b1010111010101101001: color_data = Z;
		19'b1010111010101101010: color_data = Z;
		19'b1010111010101101011: color_data = Z;
		19'b1010111010101101100: color_data = Z;
		19'b1010111010101110010: color_data = Z;
		19'b1010111010101110011: color_data = Z;
		19'b1010111010101110100: color_data = Z;
		19'b1010111010101110101: color_data = Z;
		19'b1010111010101110110: color_data = Z;
		19'b1010111010101110111: color_data = Z;
		19'b1010111010110011101: color_data = Z;
		19'b1010111010110011110: color_data = Z;
		19'b1010111010110011111: color_data = Z;
		19'b1010111010110100000: color_data = Z;
		19'b1010111010110100001: color_data = Z;
		19'b1010111010110100010: color_data = Z;
		19'b1010111010110100011: color_data = Z;
		19'b1010111010110100100: color_data = Z;
		19'b1010111010110100101: color_data = Z;
		19'b1010111010110100110: color_data = Z;
		19'b1010111100011011100: color_data = Z;
		19'b1010111100011011101: color_data = Z;
		19'b1010111100011011111: color_data = Z;
		19'b1010111100011100000: color_data = Z;
		19'b1010111100011100001: color_data = Z;
		19'b1010111100011100010: color_data = Z;
		19'b1010111100011100101: color_data = Z;
		19'b1010111100011100110: color_data = Z;
		19'b1010111100011100111: color_data = Z;
		19'b1010111100011101000: color_data = Z;
		19'b1010111100011101001: color_data = Z;
		19'b1010111100011101010: color_data = Z;
		19'b1010111100011101011: color_data = Z;
		19'b1010111100011101100: color_data = Z;
		19'b1010111100011101101: color_data = Z;
		19'b1010111100011101110: color_data = Z;
		19'b1010111100011101111: color_data = Z;
		19'b1010111100011110000: color_data = Z;
		19'b1010111100011110001: color_data = Z;
		19'b1010111100011110010: color_data = Z;
		19'b1010111100011110011: color_data = Z;
		19'b1010111100011110100: color_data = Z;
		19'b1010111100011110101: color_data = Z;
		19'b1010111100011110110: color_data = Z;
		19'b1010111100011110111: color_data = Z;
		19'b1010111100011111000: color_data = Z;
		19'b1010111100011111001: color_data = Z;
		19'b1010111100011111010: color_data = Z;
		19'b1010111100011111011: color_data = Z;
		19'b1010111100011111100: color_data = Z;
		19'b1010111100011111101: color_data = Z;
		19'b1010111100011111110: color_data = Z;
		19'b1010111100011111111: color_data = Z;
		19'b1010111100100000000: color_data = Z;
		19'b1010111100100000001: color_data = Z;
		19'b1010111100100000010: color_data = Z;
		19'b1010111100100000011: color_data = Z;
		19'b1010111100100000100: color_data = Z;
		19'b1010111100100000101: color_data = Z;
		19'b1010111100100000110: color_data = Z;
		19'b1010111100100000111: color_data = Z;
		19'b1010111100100001000: color_data = Z;
		19'b1010111100100110100: color_data = Z;
		19'b1010111100100110101: color_data = Z;
		19'b1010111100100110110: color_data = Z;
		19'b1010111100100110111: color_data = Z;
		19'b1010111100100111000: color_data = Z;
		19'b1010111100100111001: color_data = Z;
		19'b1010111100100111010: color_data = Z;
		19'b1010111100100111011: color_data = Z;
		19'b1010111100101011010: color_data = Z;
		19'b1010111100101011011: color_data = Z;
		19'b1010111100101011100: color_data = Z;
		19'b1010111100101100101: color_data = Z;
		19'b1010111100101100110: color_data = Z;
		19'b1010111100101100111: color_data = Z;
		19'b1010111100101101000: color_data = Z;
		19'b1010111100101101001: color_data = Z;
		19'b1010111100101101010: color_data = Z;
		19'b1010111100101101011: color_data = Z;
		19'b1010111100101101100: color_data = Z;
		19'b1010111100101110010: color_data = Z;
		19'b1010111100101110011: color_data = Z;
		19'b1010111100101110100: color_data = Z;
		19'b1010111100101110101: color_data = Z;
		19'b1010111100101110110: color_data = Z;
		19'b1010111100110011101: color_data = Z;
		19'b1010111100110011110: color_data = Z;
		19'b1010111100110011111: color_data = Z;
		19'b1010111100110100000: color_data = Z;
		19'b1010111100110100001: color_data = Z;
		19'b1010111100110100010: color_data = Z;
		19'b1010111100110100011: color_data = Z;
		19'b1010111100110100100: color_data = Z;
		19'b1010111100110100101: color_data = Z;
		19'b1010111110011011101: color_data = Z;
		19'b1010111110011011110: color_data = Z;
		19'b1010111110011011111: color_data = Z;
		19'b1010111110011100000: color_data = Z;
		19'b1010111110011100001: color_data = Z;
		19'b1010111110011100010: color_data = Z;
		19'b1010111110011100011: color_data = Z;
		19'b1010111110011100101: color_data = Z;
		19'b1010111110011100110: color_data = Z;
		19'b1010111110011100111: color_data = Z;
		19'b1010111110011101000: color_data = Z;
		19'b1010111110011101001: color_data = Z;
		19'b1010111110011101010: color_data = Z;
		19'b1010111110011101011: color_data = Z;
		19'b1010111110011101100: color_data = Z;
		19'b1010111110011101101: color_data = Z;
		19'b1010111110011101110: color_data = Z;
		19'b1010111110011101111: color_data = Z;
		19'b1010111110011110000: color_data = Z;
		19'b1010111110011110001: color_data = Z;
		19'b1010111110011110010: color_data = Z;
		19'b1010111110011110011: color_data = Z;
		19'b1010111110011110100: color_data = Z;
		19'b1010111110011110101: color_data = Z;
		19'b1010111110011110110: color_data = Z;
		19'b1010111110011110111: color_data = Z;
		19'b1010111110011111000: color_data = Z;
		19'b1010111110011111001: color_data = Z;
		19'b1010111110011111010: color_data = Z;
		19'b1010111110011111011: color_data = Z;
		19'b1010111110011111100: color_data = Z;
		19'b1010111110011111101: color_data = Z;
		19'b1010111110011111110: color_data = Z;
		19'b1010111110011111111: color_data = Z;
		19'b1010111110100000000: color_data = Z;
		19'b1010111110100000001: color_data = Z;
		19'b1010111110100000010: color_data = Z;
		19'b1010111110100000011: color_data = Z;
		19'b1010111110100000100: color_data = Z;
		19'b1010111110100000101: color_data = Z;
		19'b1010111110100000110: color_data = Z;
		19'b1010111110100000111: color_data = Z;
		19'b1010111110100001000: color_data = Z;
		19'b1010111110100001001: color_data = Z;
		19'b1010111110100001010: color_data = Z;
		19'b1010111110100110011: color_data = Z;
		19'b1010111110100110100: color_data = Z;
		19'b1010111110100110101: color_data = Z;
		19'b1010111110100110110: color_data = Z;
		19'b1010111110100110111: color_data = Z;
		19'b1010111110100111000: color_data = Z;
		19'b1010111110100111001: color_data = Z;
		19'b1010111110100111010: color_data = Z;
		19'b1010111110100111011: color_data = Z;
		19'b1010111110101010100: color_data = Z;
		19'b1010111110101010101: color_data = Z;
		19'b1010111110101010110: color_data = Z;
		19'b1010111110101010111: color_data = Z;
		19'b1010111110101011001: color_data = Z;
		19'b1010111110101011010: color_data = Z;
		19'b1010111110101011011: color_data = Z;
		19'b1010111110101011100: color_data = Z;
		19'b1010111110101100100: color_data = Z;
		19'b1010111110101100101: color_data = Z;
		19'b1010111110101100110: color_data = Z;
		19'b1010111110101100111: color_data = Z;
		19'b1010111110101101000: color_data = Z;
		19'b1010111110101101001: color_data = Z;
		19'b1010111110101101010: color_data = Z;
		19'b1010111110101101011: color_data = Z;
		19'b1010111110101101100: color_data = Z;
		19'b1010111110101110010: color_data = Z;
		19'b1010111110101110011: color_data = Z;
		19'b1010111110101110100: color_data = Z;
		19'b1010111110101110101: color_data = Z;
		19'b1010111110101110110: color_data = Z;
		19'b1010111110110011101: color_data = Z;
		19'b1010111110110011110: color_data = Z;
		19'b1010111110110011111: color_data = Z;
		19'b1010111110110100000: color_data = Z;
		19'b1010111110110100001: color_data = Z;
		19'b1010111110110100010: color_data = Z;
		19'b1010111110110100011: color_data = Z;
		19'b1010111110110100100: color_data = Z;
		19'b1010111110110100101: color_data = Z;
		19'b1011000000011011111: color_data = Z;
		19'b1011000000011100000: color_data = Z;
		19'b1011000000011100001: color_data = Z;
		19'b1011000000011100010: color_data = Z;
		19'b1011000000011100011: color_data = Z;
		19'b1011000000011100100: color_data = Z;
		19'b1011000000011100101: color_data = Z;
		19'b1011000000011100110: color_data = Z;
		19'b1011000000011100111: color_data = Z;
		19'b1011000000011101000: color_data = Z;
		19'b1011000000011101001: color_data = Z;
		19'b1011000000011101010: color_data = Z;
		19'b1011000000011101011: color_data = Z;
		19'b1011000000011101100: color_data = Z;
		19'b1011000000011101101: color_data = Z;
		19'b1011000000011101110: color_data = Z;
		19'b1011000000011101111: color_data = Z;
		19'b1011000000011110000: color_data = Z;
		19'b1011000000011110001: color_data = Z;
		19'b1011000000011110010: color_data = Z;
		19'b1011000000011110011: color_data = Z;
		19'b1011000000011110100: color_data = Z;
		19'b1011000000011110101: color_data = Z;
		19'b1011000000011110110: color_data = Z;
		19'b1011000000011110111: color_data = Z;
		19'b1011000000011111000: color_data = Z;
		19'b1011000000011111001: color_data = Z;
		19'b1011000000011111010: color_data = Z;
		19'b1011000000011111011: color_data = Z;
		19'b1011000000011111100: color_data = Z;
		19'b1011000000011111101: color_data = Z;
		19'b1011000000011111110: color_data = Z;
		19'b1011000000011111111: color_data = Z;
		19'b1011000000100000000: color_data = Z;
		19'b1011000000100000001: color_data = Z;
		19'b1011000000100000010: color_data = Z;
		19'b1011000000100000011: color_data = Z;
		19'b1011000000100000100: color_data = Z;
		19'b1011000000100000101: color_data = Z;
		19'b1011000000100000110: color_data = Z;
		19'b1011000000100000111: color_data = Z;
		19'b1011000000100001000: color_data = Z;
		19'b1011000000100001001: color_data = Z;
		19'b1011000000100001010: color_data = Z;
		19'b1011000000100001011: color_data = Z;
		19'b1011000000100110011: color_data = Z;
		19'b1011000000100110100: color_data = Z;
		19'b1011000000100110101: color_data = Z;
		19'b1011000000100110110: color_data = Z;
		19'b1011000000100110111: color_data = Z;
		19'b1011000000100111000: color_data = Z;
		19'b1011000000100111001: color_data = Z;
		19'b1011000000100111010: color_data = Z;
		19'b1011000000100111011: color_data = Z;
		19'b1011000000101010000: color_data = Z;
		19'b1011000000101010001: color_data = Z;
		19'b1011000000101010010: color_data = Z;
		19'b1011000000101010011: color_data = Z;
		19'b1011000000101010100: color_data = Z;
		19'b1011000000101010101: color_data = Z;
		19'b1011000000101010110: color_data = Z;
		19'b1011000000101010111: color_data = Z;
		19'b1011000000101011000: color_data = Z;
		19'b1011000000101011001: color_data = Z;
		19'b1011000000101011010: color_data = Z;
		19'b1011000000101011011: color_data = Z;
		19'b1011000000101011100: color_data = Z;
		19'b1011000000101100100: color_data = Z;
		19'b1011000000101100101: color_data = Z;
		19'b1011000000101100110: color_data = Z;
		19'b1011000000101100111: color_data = Z;
		19'b1011000000101101000: color_data = Z;
		19'b1011000000101101001: color_data = Z;
		19'b1011000000101101010: color_data = Z;
		19'b1011000000101101011: color_data = Z;
		19'b1011000000101101100: color_data = Z;
		19'b1011000000101110001: color_data = Z;
		19'b1011000000101110010: color_data = Z;
		19'b1011000000101110011: color_data = Z;
		19'b1011000000101110100: color_data = Z;
		19'b1011000000101110101: color_data = Z;
		19'b1011000000110011100: color_data = Z;
		19'b1011000000110011101: color_data = Z;
		19'b1011000000110011110: color_data = Z;
		19'b1011000000110011111: color_data = Z;
		19'b1011000000110100000: color_data = Z;
		19'b1011000000110100001: color_data = Z;
		19'b1011000000110100010: color_data = Z;
		19'b1011000000110100011: color_data = Z;
		19'b1011000000110100100: color_data = Z;
		19'b1011000010011100000: color_data = Z;
		19'b1011000010011100001: color_data = Z;
		19'b1011000010011100010: color_data = Z;
		19'b1011000010011100011: color_data = Z;
		19'b1011000010011100100: color_data = Z;
		19'b1011000010011100101: color_data = Z;
		19'b1011000010011100110: color_data = Z;
		19'b1011000010011100111: color_data = Z;
		19'b1011000010011101000: color_data = Z;
		19'b1011000010011101001: color_data = Z;
		19'b1011000010011101010: color_data = Z;
		19'b1011000010011101011: color_data = Z;
		19'b1011000010011101100: color_data = Z;
		19'b1011000010011101101: color_data = Z;
		19'b1011000010011101110: color_data = Z;
		19'b1011000010011101111: color_data = Z;
		19'b1011000010011110000: color_data = Z;
		19'b1011000010011110001: color_data = Z;
		19'b1011000010011110010: color_data = Z;
		19'b1011000010011110011: color_data = Z;
		19'b1011000010011110100: color_data = Z;
		19'b1011000010011110101: color_data = Z;
		19'b1011000010011110110: color_data = Z;
		19'b1011000010011110111: color_data = Z;
		19'b1011000010011111000: color_data = Z;
		19'b1011000010011111001: color_data = Z;
		19'b1011000010011111010: color_data = Z;
		19'b1011000010011111011: color_data = Z;
		19'b1011000010011111100: color_data = Z;
		19'b1011000010011111101: color_data = Z;
		19'b1011000010011111110: color_data = Z;
		19'b1011000010011111111: color_data = Z;
		19'b1011000010100000000: color_data = Z;
		19'b1011000010100000001: color_data = Z;
		19'b1011000010100000010: color_data = Z;
		19'b1011000010100000011: color_data = Z;
		19'b1011000010100000100: color_data = Z;
		19'b1011000010100000101: color_data = Z;
		19'b1011000010100000110: color_data = Z;
		19'b1011000010100000111: color_data = Z;
		19'b1011000010100001000: color_data = Z;
		19'b1011000010100001001: color_data = Z;
		19'b1011000010100001010: color_data = Z;
		19'b1011000010100001011: color_data = Z;
		19'b1011000010100001100: color_data = Z;
		19'b1011000010100110011: color_data = Z;
		19'b1011000010100110100: color_data = Z;
		19'b1011000010100110101: color_data = Z;
		19'b1011000010100110110: color_data = Z;
		19'b1011000010100110111: color_data = Z;
		19'b1011000010100111000: color_data = Z;
		19'b1011000010100111001: color_data = Z;
		19'b1011000010100111010: color_data = Z;
		19'b1011000010100111011: color_data = Z;
		19'b1011000010101001111: color_data = Z;
		19'b1011000010101010000: color_data = Z;
		19'b1011000010101010001: color_data = Z;
		19'b1011000010101010010: color_data = Z;
		19'b1011000010101010011: color_data = Z;
		19'b1011000010101010100: color_data = Z;
		19'b1011000010101010101: color_data = Z;
		19'b1011000010101010110: color_data = Z;
		19'b1011000010101010111: color_data = Z;
		19'b1011000010101011000: color_data = Z;
		19'b1011000010101011001: color_data = Z;
		19'b1011000010101011010: color_data = Z;
		19'b1011000010101011011: color_data = Z;
		19'b1011000010101011100: color_data = Z;
		19'b1011000010101100100: color_data = Z;
		19'b1011000010101100101: color_data = Z;
		19'b1011000010101100110: color_data = Z;
		19'b1011000010101100111: color_data = Z;
		19'b1011000010101101000: color_data = Z;
		19'b1011000010101101001: color_data = Z;
		19'b1011000010101101010: color_data = Z;
		19'b1011000010101101011: color_data = Z;
		19'b1011000010101101100: color_data = Z;
		19'b1011000010101110001: color_data = Z;
		19'b1011000010101110010: color_data = Z;
		19'b1011000010101110011: color_data = Z;
		19'b1011000010110011100: color_data = Z;
		19'b1011000010110011101: color_data = Z;
		19'b1011000010110011110: color_data = Z;
		19'b1011000010110011111: color_data = Z;
		19'b1011000010110100000: color_data = Z;
		19'b1011000010110100001: color_data = Z;
		19'b1011000010110100010: color_data = Z;
		19'b1011000010110100011: color_data = Z;
		19'b1011000010110100100: color_data = Z;
		19'b1011000100011100010: color_data = Z;
		19'b1011000100011100011: color_data = Z;
		19'b1011000100011100100: color_data = Z;
		19'b1011000100011100101: color_data = Z;
		19'b1011000100011100110: color_data = Z;
		19'b1011000100011100111: color_data = Z;
		19'b1011000100011101000: color_data = Z;
		19'b1011000100011101001: color_data = Z;
		19'b1011000100011101010: color_data = Z;
		19'b1011000100011101011: color_data = Z;
		19'b1011000100011101100: color_data = Z;
		19'b1011000100011101101: color_data = Z;
		19'b1011000100011101110: color_data = Z;
		19'b1011000100011101111: color_data = Z;
		19'b1011000100011110000: color_data = Z;
		19'b1011000100011110001: color_data = Z;
		19'b1011000100011110010: color_data = Z;
		19'b1011000100011110011: color_data = Z;
		19'b1011000100011110100: color_data = Z;
		19'b1011000100011110101: color_data = Z;
		19'b1011000100011110110: color_data = Z;
		19'b1011000100011110111: color_data = Z;
		19'b1011000100011111000: color_data = Z;
		19'b1011000100011111001: color_data = Z;
		19'b1011000100011111010: color_data = Z;
		19'b1011000100011111011: color_data = Z;
		19'b1011000100011111100: color_data = Z;
		19'b1011000100011111101: color_data = Z;
		19'b1011000100011111110: color_data = Z;
		19'b1011000100011111111: color_data = Z;
		19'b1011000100100000000: color_data = Z;
		19'b1011000100100000001: color_data = Z;
		19'b1011000100100000010: color_data = Z;
		19'b1011000100100000011: color_data = Z;
		19'b1011000100100000100: color_data = Z;
		19'b1011000100100000101: color_data = Z;
		19'b1011000100100000110: color_data = Z;
		19'b1011000100100000111: color_data = Z;
		19'b1011000100100001000: color_data = Z;
		19'b1011000100100001001: color_data = Z;
		19'b1011000100100001010: color_data = Z;
		19'b1011000100100001011: color_data = Z;
		19'b1011000100100001100: color_data = Z;
		19'b1011000100100001101: color_data = Z;
		19'b1011000100100110010: color_data = Z;
		19'b1011000100100110011: color_data = Z;
		19'b1011000100100110100: color_data = Z;
		19'b1011000100100110101: color_data = Z;
		19'b1011000100100110110: color_data = Z;
		19'b1011000100100110111: color_data = Z;
		19'b1011000100100111000: color_data = Z;
		19'b1011000100100111001: color_data = Z;
		19'b1011000100100111010: color_data = Z;
		19'b1011000100100111011: color_data = Z;
		19'b1011000100101000000: color_data = Z;
		19'b1011000100101000001: color_data = Z;
		19'b1011000100101001111: color_data = Z;
		19'b1011000100101010000: color_data = Z;
		19'b1011000100101010001: color_data = Z;
		19'b1011000100101010010: color_data = Z;
		19'b1011000100101010011: color_data = Z;
		19'b1011000100101010100: color_data = Z;
		19'b1011000100101010101: color_data = Z;
		19'b1011000100101010110: color_data = Z;
		19'b1011000100101010111: color_data = Z;
		19'b1011000100101011000: color_data = Z;
		19'b1011000100101011001: color_data = Z;
		19'b1011000100101011010: color_data = Z;
		19'b1011000100101011011: color_data = Z;
		19'b1011000100101100011: color_data = Z;
		19'b1011000100101100100: color_data = Z;
		19'b1011000100101100101: color_data = Z;
		19'b1011000100101100110: color_data = Z;
		19'b1011000100101100111: color_data = Z;
		19'b1011000100101101000: color_data = Z;
		19'b1011000100101101001: color_data = Z;
		19'b1011000100101101010: color_data = Z;
		19'b1011000100101101011: color_data = Z;
		19'b1011000100101110010: color_data = Z;
		19'b1011000100110011011: color_data = Z;
		19'b1011000100110011100: color_data = Z;
		19'b1011000100110011101: color_data = Z;
		19'b1011000100110011110: color_data = Z;
		19'b1011000100110011111: color_data = Z;
		19'b1011000100110100000: color_data = Z;
		19'b1011000100110100001: color_data = Z;
		19'b1011000100110100010: color_data = Z;
		19'b1011000100110100011: color_data = Z;
		19'b1011000110011100011: color_data = Z;
		19'b1011000110011100100: color_data = Z;
		19'b1011000110011100101: color_data = Z;
		19'b1011000110011100110: color_data = Z;
		19'b1011000110011100111: color_data = Z;
		19'b1011000110011101000: color_data = Z;
		19'b1011000110011101001: color_data = Z;
		19'b1011000110011101010: color_data = Z;
		19'b1011000110011101011: color_data = Z;
		19'b1011000110011101100: color_data = Z;
		19'b1011000110011101101: color_data = Z;
		19'b1011000110011101110: color_data = Z;
		19'b1011000110011101111: color_data = Z;
		19'b1011000110011110000: color_data = Z;
		19'b1011000110011110001: color_data = Z;
		19'b1011000110011110010: color_data = Z;
		19'b1011000110011110011: color_data = Z;
		19'b1011000110011110100: color_data = Z;
		19'b1011000110011110101: color_data = Z;
		19'b1011000110011110110: color_data = Z;
		19'b1011000110011110111: color_data = Z;
		19'b1011000110011111000: color_data = Z;
		19'b1011000110011111001: color_data = Z;
		19'b1011000110011111010: color_data = Z;
		19'b1011000110011111011: color_data = Z;
		19'b1011000110011111100: color_data = Z;
		19'b1011000110011111101: color_data = Z;
		19'b1011000110011111110: color_data = Z;
		19'b1011000110011111111: color_data = Z;
		19'b1011000110100000000: color_data = Z;
		19'b1011000110100000001: color_data = Z;
		19'b1011000110100000010: color_data = Z;
		19'b1011000110100000011: color_data = Z;
		19'b1011000110100000100: color_data = Z;
		19'b1011000110100000101: color_data = Z;
		19'b1011000110100000110: color_data = Z;
		19'b1011000110100000111: color_data = Z;
		19'b1011000110100001000: color_data = Z;
		19'b1011000110100001001: color_data = Z;
		19'b1011000110100001010: color_data = Z;
		19'b1011000110100001011: color_data = Z;
		19'b1011000110100001100: color_data = Z;
		19'b1011000110100001101: color_data = Z;
		19'b1011000110100001110: color_data = Z;
		19'b1011000110100001111: color_data = Z;
		19'b1011000110100101010: color_data = Z;
		19'b1011000110100110010: color_data = Z;
		19'b1011000110100110011: color_data = Z;
		19'b1011000110100110100: color_data = Z;
		19'b1011000110100110101: color_data = Z;
		19'b1011000110100110110: color_data = Z;
		19'b1011000110100110111: color_data = Z;
		19'b1011000110100111000: color_data = Z;
		19'b1011000110100111001: color_data = Z;
		19'b1011000110100111010: color_data = Z;
		19'b1011000110100111011: color_data = Z;
		19'b1011000110101000000: color_data = Z;
		19'b1011000110101000001: color_data = Z;
		19'b1011000110101000010: color_data = Z;
		19'b1011000110101000011: color_data = Z;
		19'b1011000110101001111: color_data = Z;
		19'b1011000110101010000: color_data = Z;
		19'b1011000110101010001: color_data = Z;
		19'b1011000110101010010: color_data = Z;
		19'b1011000110101010011: color_data = Z;
		19'b1011000110101010100: color_data = Z;
		19'b1011000110101010101: color_data = Z;
		19'b1011000110101010110: color_data = Z;
		19'b1011000110101010111: color_data = Z;
		19'b1011000110101011000: color_data = Z;
		19'b1011000110101011001: color_data = Z;
		19'b1011000110101011010: color_data = Z;
		19'b1011000110101011011: color_data = Z;
		19'b1011000110101100011: color_data = Z;
		19'b1011000110101100100: color_data = Z;
		19'b1011000110101100101: color_data = Z;
		19'b1011000110101100110: color_data = Z;
		19'b1011000110101100111: color_data = Z;
		19'b1011000110101101000: color_data = Z;
		19'b1011000110101101001: color_data = Z;
		19'b1011000110101101010: color_data = Z;
		19'b1011000110101101011: color_data = Z;
		19'b1011000110110011010: color_data = Z;
		19'b1011000110110011011: color_data = Z;
		19'b1011000110110011100: color_data = Z;
		19'b1011000110110011101: color_data = Z;
		19'b1011000110110011110: color_data = Z;
		19'b1011000110110011111: color_data = Z;
		19'b1011000110110100000: color_data = Z;
		19'b1011000110110100001: color_data = Z;
		19'b1011000110110100010: color_data = Z;
		19'b1011001000011100100: color_data = Z;
		19'b1011001000011100101: color_data = Z;
		19'b1011001000011100110: color_data = Z;
		19'b1011001000011100111: color_data = Z;
		19'b1011001000011101000: color_data = Z;
		19'b1011001000011101001: color_data = Z;
		19'b1011001000011101010: color_data = Z;
		19'b1011001000011101011: color_data = Z;
		19'b1011001000011101100: color_data = Z;
		19'b1011001000011101101: color_data = Z;
		19'b1011001000011101110: color_data = Z;
		19'b1011001000011101111: color_data = Z;
		19'b1011001000011110000: color_data = Z;
		19'b1011001000011110001: color_data = Z;
		19'b1011001000011110010: color_data = Z;
		19'b1011001000011110011: color_data = Z;
		19'b1011001000011110100: color_data = Z;
		19'b1011001000011110101: color_data = Z;
		19'b1011001000011110110: color_data = Z;
		19'b1011001000011110111: color_data = Z;
		19'b1011001000011111000: color_data = Z;
		19'b1011001000011111001: color_data = Z;
		19'b1011001000011111010: color_data = Z;
		19'b1011001000011111011: color_data = Z;
		19'b1011001000011111100: color_data = Z;
		19'b1011001000011111101: color_data = Z;
		19'b1011001000011111110: color_data = Z;
		19'b1011001000011111111: color_data = Z;
		19'b1011001000100000000: color_data = Z;
		19'b1011001000100000001: color_data = Z;
		19'b1011001000100000010: color_data = Z;
		19'b1011001000100000011: color_data = Z;
		19'b1011001000100000100: color_data = Z;
		19'b1011001000100000101: color_data = Z;
		19'b1011001000100000110: color_data = Z;
		19'b1011001000100000111: color_data = Z;
		19'b1011001000100001000: color_data = Z;
		19'b1011001000100001001: color_data = Z;
		19'b1011001000100001010: color_data = Z;
		19'b1011001000100001011: color_data = Z;
		19'b1011001000100001100: color_data = Z;
		19'b1011001000100001101: color_data = Z;
		19'b1011001000100001110: color_data = Z;
		19'b1011001000100001111: color_data = Z;
		19'b1011001000100010000: color_data = Z;
		19'b1011001000100010001: color_data = Z;
		19'b1011001000100010010: color_data = Z;
		19'b1011001000100101010: color_data = Z;
		19'b1011001000100110010: color_data = Z;
		19'b1011001000100110011: color_data = Z;
		19'b1011001000100110100: color_data = Z;
		19'b1011001000100110101: color_data = Z;
		19'b1011001000100110110: color_data = Z;
		19'b1011001000100110111: color_data = Z;
		19'b1011001000100111000: color_data = Z;
		19'b1011001000100111001: color_data = Z;
		19'b1011001000100111010: color_data = Z;
		19'b1011001000100111011: color_data = Z;
		19'b1011001000101000000: color_data = Z;
		19'b1011001000101000001: color_data = Z;
		19'b1011001000101000010: color_data = Z;
		19'b1011001000101000011: color_data = Z;
		19'b1011001000101000100: color_data = Z;
		19'b1011001000101000101: color_data = Z;
		19'b1011001000101000110: color_data = Z;
		19'b1011001000101001110: color_data = Z;
		19'b1011001000101001111: color_data = Z;
		19'b1011001000101010000: color_data = Z;
		19'b1011001000101010001: color_data = Z;
		19'b1011001000101010010: color_data = Z;
		19'b1011001000101010011: color_data = Z;
		19'b1011001000101010100: color_data = Z;
		19'b1011001000101010101: color_data = Z;
		19'b1011001000101010110: color_data = Z;
		19'b1011001000101010111: color_data = Z;
		19'b1011001000101011000: color_data = Z;
		19'b1011001000101011001: color_data = Z;
		19'b1011001000101011010: color_data = Z;
		19'b1011001000101011011: color_data = Z;
		19'b1011001000101100011: color_data = Z;
		19'b1011001000101100100: color_data = Z;
		19'b1011001000101100101: color_data = Z;
		19'b1011001000101100110: color_data = Z;
		19'b1011001000101100111: color_data = Z;
		19'b1011001000101101000: color_data = Z;
		19'b1011001000101101001: color_data = Z;
		19'b1011001000101101010: color_data = Z;
		19'b1011001000101101011: color_data = Z;
		19'b1011001000101101100: color_data = Z;
		19'b1011001000110011000: color_data = Z;
		19'b1011001000110011001: color_data = Z;
		19'b1011001000110011010: color_data = Z;
		19'b1011001000110011011: color_data = Z;
		19'b1011001000110011100: color_data = Z;
		19'b1011001000110011101: color_data = Z;
		19'b1011001000110011110: color_data = Z;
		19'b1011001000110011111: color_data = Z;
		19'b1011001000110100000: color_data = Z;
		19'b1011001000110100001: color_data = Z;
		19'b1011001010011100101: color_data = Z;
		19'b1011001010011100110: color_data = Z;
		19'b1011001010011100111: color_data = Z;
		19'b1011001010011101000: color_data = Z;
		19'b1011001010011101001: color_data = Z;
		19'b1011001010011101010: color_data = Z;
		19'b1011001010011101011: color_data = Z;
		19'b1011001010011101100: color_data = Z;
		19'b1011001010011101101: color_data = Z;
		19'b1011001010011101110: color_data = Z;
		19'b1011001010011101111: color_data = Z;
		19'b1011001010011110000: color_data = Z;
		19'b1011001010011110001: color_data = Z;
		19'b1011001010011110010: color_data = Z;
		19'b1011001010011110011: color_data = Z;
		19'b1011001010011110100: color_data = Z;
		19'b1011001010011110101: color_data = Z;
		19'b1011001010011110110: color_data = Z;
		19'b1011001010011110111: color_data = Z;
		19'b1011001010011111000: color_data = Z;
		19'b1011001010011111001: color_data = Z;
		19'b1011001010011111010: color_data = Z;
		19'b1011001010011111011: color_data = Z;
		19'b1011001010011111100: color_data = Z;
		19'b1011001010011111101: color_data = Z;
		19'b1011001010011111110: color_data = Z;
		19'b1011001010011111111: color_data = Z;
		19'b1011001010100000000: color_data = Z;
		19'b1011001010100000001: color_data = Z;
		19'b1011001010100000010: color_data = Z;
		19'b1011001010100000011: color_data = Z;
		19'b1011001010100000100: color_data = Z;
		19'b1011001010100000101: color_data = Z;
		19'b1011001010100000110: color_data = Z;
		19'b1011001010100000111: color_data = Z;
		19'b1011001010100001000: color_data = Z;
		19'b1011001010100001001: color_data = Z;
		19'b1011001010100001010: color_data = Z;
		19'b1011001010100001011: color_data = Z;
		19'b1011001010100001100: color_data = Z;
		19'b1011001010100001101: color_data = Z;
		19'b1011001010100001110: color_data = Z;
		19'b1011001010100001111: color_data = Z;
		19'b1011001010100010000: color_data = Z;
		19'b1011001010100010001: color_data = Z;
		19'b1011001010100010010: color_data = Z;
		19'b1011001010100010011: color_data = Z;
		19'b1011001010100010100: color_data = Z;
		19'b1011001010100110010: color_data = Z;
		19'b1011001010100110011: color_data = Z;
		19'b1011001010100110100: color_data = Z;
		19'b1011001010100110110: color_data = Z;
		19'b1011001010100110111: color_data = Z;
		19'b1011001010100111000: color_data = Z;
		19'b1011001010100111001: color_data = Z;
		19'b1011001010100111010: color_data = Z;
		19'b1011001010100111011: color_data = Z;
		19'b1011001010101000000: color_data = Z;
		19'b1011001010101000001: color_data = Z;
		19'b1011001010101000010: color_data = Z;
		19'b1011001010101000011: color_data = Z;
		19'b1011001010101000100: color_data = Z;
		19'b1011001010101000101: color_data = Z;
		19'b1011001010101000110: color_data = Z;
		19'b1011001010101001110: color_data = Z;
		19'b1011001010101001111: color_data = Z;
		19'b1011001010101010000: color_data = Z;
		19'b1011001010101010001: color_data = Z;
		19'b1011001010101010010: color_data = Z;
		19'b1011001010101010011: color_data = Z;
		19'b1011001010101010100: color_data = Z;
		19'b1011001010101010101: color_data = Z;
		19'b1011001010101010110: color_data = Z;
		19'b1011001010101010111: color_data = Z;
		19'b1011001010101011000: color_data = Z;
		19'b1011001010101011001: color_data = Z;
		19'b1011001010101011010: color_data = Z;
		19'b1011001010101011011: color_data = Z;
		19'b1011001010101100011: color_data = Z;
		19'b1011001010101100100: color_data = Z;
		19'b1011001010101100101: color_data = Z;
		19'b1011001010101100110: color_data = Z;
		19'b1011001010101100111: color_data = Z;
		19'b1011001010101101000: color_data = Z;
		19'b1011001010101101001: color_data = Z;
		19'b1011001010101101010: color_data = Z;
		19'b1011001010101101011: color_data = Z;
		19'b1011001010110010110: color_data = Z;
		19'b1011001010110010111: color_data = Z;
		19'b1011001010110011000: color_data = Z;
		19'b1011001010110011001: color_data = Z;
		19'b1011001010110011010: color_data = Z;
		19'b1011001010110011011: color_data = Z;
		19'b1011001010110011100: color_data = Z;
		19'b1011001010110011101: color_data = Z;
		19'b1011001010110011110: color_data = Z;
		19'b1011001010110011111: color_data = Z;
		19'b1011001010110100000: color_data = Z;
		19'b1011001100011100111: color_data = Z;
		19'b1011001100011101000: color_data = Z;
		19'b1011001100011101001: color_data = Z;
		19'b1011001100011101010: color_data = Z;
		19'b1011001100011101011: color_data = Z;
		19'b1011001100011101100: color_data = Z;
		19'b1011001100011101101: color_data = Z;
		19'b1011001100011101110: color_data = Z;
		19'b1011001100011101111: color_data = Z;
		19'b1011001100011110000: color_data = Z;
		19'b1011001100011110001: color_data = Z;
		19'b1011001100011110010: color_data = Z;
		19'b1011001100011110011: color_data = Z;
		19'b1011001100011110100: color_data = Z;
		19'b1011001100011110101: color_data = Z;
		19'b1011001100011110110: color_data = Z;
		19'b1011001100011110111: color_data = Z;
		19'b1011001100011111000: color_data = Z;
		19'b1011001100011111001: color_data = Z;
		19'b1011001100011111010: color_data = Z;
		19'b1011001100011111011: color_data = Z;
		19'b1011001100011111100: color_data = Z;
		19'b1011001100011111101: color_data = Z;
		19'b1011001100011111110: color_data = Z;
		19'b1011001100011111111: color_data = Z;
		19'b1011001100100000000: color_data = Z;
		19'b1011001100100000001: color_data = Z;
		19'b1011001100100000010: color_data = Z;
		19'b1011001100100000011: color_data = Z;
		19'b1011001100100000100: color_data = Z;
		19'b1011001100100000101: color_data = Z;
		19'b1011001100100000110: color_data = Z;
		19'b1011001100100000111: color_data = Z;
		19'b1011001100100001000: color_data = Z;
		19'b1011001100100001001: color_data = Z;
		19'b1011001100100001010: color_data = Z;
		19'b1011001100100001011: color_data = Z;
		19'b1011001100100001100: color_data = Z;
		19'b1011001100100001101: color_data = Z;
		19'b1011001100100001110: color_data = Z;
		19'b1011001100100001111: color_data = Z;
		19'b1011001100100010000: color_data = Z;
		19'b1011001100100010001: color_data = Z;
		19'b1011001100100010010: color_data = Z;
		19'b1011001100100010011: color_data = Z;
		19'b1011001100100010100: color_data = Z;
		19'b1011001100100010101: color_data = Z;
		19'b1011001100100010110: color_data = Z;
		19'b1011001100100010111: color_data = Z;
		19'b1011001100100011000: color_data = Z;
		19'b1011001100100110111: color_data = Z;
		19'b1011001100100111000: color_data = Z;
		19'b1011001100100111001: color_data = Z;
		19'b1011001100100111010: color_data = Z;
		19'b1011001100100111011: color_data = Z;
		19'b1011001100101000000: color_data = Z;
		19'b1011001100101000001: color_data = Z;
		19'b1011001100101000010: color_data = Z;
		19'b1011001100101000011: color_data = Z;
		19'b1011001100101000100: color_data = Z;
		19'b1011001100101000101: color_data = Z;
		19'b1011001100101000110: color_data = Z;
		19'b1011001100101001110: color_data = Z;
		19'b1011001100101001111: color_data = Z;
		19'b1011001100101010000: color_data = Z;
		19'b1011001100101010001: color_data = Z;
		19'b1011001100101010010: color_data = Z;
		19'b1011001100101010011: color_data = Z;
		19'b1011001100101010101: color_data = Z;
		19'b1011001100101010110: color_data = Z;
		19'b1011001100101010111: color_data = Z;
		19'b1011001100101011000: color_data = Z;
		19'b1011001100101011001: color_data = Z;
		19'b1011001100101011010: color_data = Z;
		19'b1011001100101011011: color_data = Z;
		19'b1011001100101100011: color_data = Z;
		19'b1011001100101100100: color_data = Z;
		19'b1011001100101100101: color_data = Z;
		19'b1011001100101100110: color_data = Z;
		19'b1011001100101100111: color_data = Z;
		19'b1011001100101101000: color_data = Z;
		19'b1011001100101101001: color_data = Z;
		19'b1011001100110010010: color_data = Z;
		19'b1011001100110010011: color_data = Z;
		19'b1011001100110010100: color_data = Z;
		19'b1011001100110010101: color_data = Z;
		19'b1011001100110010110: color_data = Z;
		19'b1011001100110010111: color_data = Z;
		19'b1011001100110011000: color_data = Z;
		19'b1011001100110011001: color_data = Z;
		19'b1011001100110011010: color_data = Z;
		19'b1011001100110011011: color_data = Z;
		19'b1011001100110011100: color_data = Z;
		19'b1011001100110011101: color_data = Z;
		19'b1011001100110011110: color_data = Z;
		19'b1011001100110011111: color_data = Z;
		19'b1011001110011101000: color_data = Z;
		19'b1011001110011101001: color_data = Z;
		19'b1011001110011101010: color_data = Z;
		19'b1011001110011101011: color_data = Z;
		19'b1011001110011101100: color_data = Z;
		19'b1011001110011101101: color_data = Z;
		19'b1011001110011101110: color_data = Z;
		19'b1011001110011101111: color_data = Z;
		19'b1011001110011110000: color_data = Z;
		19'b1011001110011110001: color_data = Z;
		19'b1011001110011110010: color_data = Z;
		19'b1011001110011110011: color_data = Z;
		19'b1011001110011110100: color_data = Z;
		19'b1011001110011110101: color_data = Z;
		19'b1011001110011110110: color_data = Z;
		19'b1011001110011110111: color_data = Z;
		19'b1011001110011111000: color_data = Z;
		19'b1011001110011111001: color_data = Z;
		19'b1011001110011111010: color_data = Z;
		19'b1011001110011111011: color_data = Z;
		19'b1011001110011111100: color_data = Z;
		19'b1011001110011111101: color_data = Z;
		19'b1011001110011111110: color_data = Z;
		19'b1011001110011111111: color_data = Z;
		19'b1011001110100000000: color_data = Z;
		19'b1011001110100000001: color_data = Z;
		19'b1011001110100000010: color_data = Z;
		19'b1011001110100000011: color_data = Z;
		19'b1011001110100000100: color_data = Z;
		19'b1011001110100000101: color_data = Z;
		19'b1011001110100000110: color_data = Z;
		19'b1011001110100000111: color_data = Z;
		19'b1011001110100001000: color_data = Z;
		19'b1011001110100001001: color_data = Z;
		19'b1011001110100001010: color_data = Z;
		19'b1011001110100001011: color_data = Z;
		19'b1011001110100001100: color_data = Z;
		19'b1011001110100001101: color_data = Z;
		19'b1011001110100001110: color_data = Z;
		19'b1011001110100001111: color_data = Z;
		19'b1011001110100010000: color_data = Z;
		19'b1011001110100010001: color_data = Z;
		19'b1011001110100010010: color_data = Z;
		19'b1011001110100010011: color_data = Z;
		19'b1011001110100010100: color_data = Z;
		19'b1011001110100010101: color_data = Z;
		19'b1011001110100010110: color_data = Z;
		19'b1011001110100010111: color_data = Z;
		19'b1011001110100011000: color_data = Z;
		19'b1011001110100011001: color_data = Z;
		19'b1011001110100011010: color_data = Z;
		19'b1011001110100111000: color_data = Z;
		19'b1011001110100111001: color_data = Z;
		19'b1011001110100111010: color_data = Z;
		19'b1011001110100111011: color_data = Z;
		19'b1011001110101000000: color_data = Z;
		19'b1011001110101000001: color_data = Z;
		19'b1011001110101000010: color_data = Z;
		19'b1011001110101000011: color_data = Z;
		19'b1011001110101000100: color_data = Z;
		19'b1011001110101000101: color_data = Z;
		19'b1011001110101001110: color_data = Z;
		19'b1011001110101001111: color_data = Z;
		19'b1011001110101010000: color_data = Z;
		19'b1011001110101010001: color_data = Z;
		19'b1011001110101010010: color_data = Z;
		19'b1011001110101010011: color_data = Z;
		19'b1011001110101010101: color_data = Z;
		19'b1011001110101010110: color_data = Z;
		19'b1011001110101010111: color_data = Z;
		19'b1011001110101011000: color_data = Z;
		19'b1011001110101011001: color_data = Z;
		19'b1011001110101011010: color_data = Z;
		19'b1011001110101011011: color_data = Z;
		19'b1011001110101100011: color_data = Z;
		19'b1011001110101100101: color_data = Z;
		19'b1011001110101100110: color_data = Z;
		19'b1011001110101100111: color_data = Z;
		19'b1011001110101101000: color_data = Z;
		19'b1011001110110001100: color_data = Z;
		19'b1011001110110001101: color_data = Z;
		19'b1011001110110001110: color_data = Z;
		19'b1011001110110001111: color_data = Z;
		19'b1011001110110010000: color_data = Z;
		19'b1011001110110010001: color_data = Z;
		19'b1011001110110010010: color_data = Z;
		19'b1011001110110010011: color_data = Z;
		19'b1011001110110010100: color_data = Z;
		19'b1011001110110010101: color_data = Z;
		19'b1011001110110010110: color_data = Z;
		19'b1011001110110010111: color_data = Z;
		19'b1011001110110011000: color_data = Z;
		19'b1011001110110011001: color_data = Z;
		19'b1011001110110011010: color_data = Z;
		19'b1011001110110011011: color_data = Z;
		19'b1011001110110011100: color_data = Z;
		19'b1011001110110011101: color_data = Z;
		19'b1011001110110011110: color_data = Z;
		19'b1011010000011101001: color_data = Z;
		19'b1011010000011101010: color_data = Z;
		19'b1011010000011101011: color_data = Z;
		19'b1011010000011101100: color_data = Z;
		19'b1011010000011101101: color_data = Z;
		19'b1011010000011101110: color_data = Z;
		19'b1011010000011101111: color_data = Z;
		19'b1011010000011110000: color_data = Z;
		19'b1011010000011110001: color_data = Z;
		19'b1011010000011110010: color_data = Z;
		19'b1011010000011110011: color_data = Z;
		19'b1011010000011110100: color_data = Z;
		19'b1011010000011110101: color_data = Z;
		19'b1011010000011110110: color_data = Z;
		19'b1011010000011110111: color_data = Z;
		19'b1011010000011111000: color_data = Z;
		19'b1011010000011111001: color_data = Z;
		19'b1011010000011111010: color_data = Z;
		19'b1011010000011111011: color_data = Z;
		19'b1011010000011111100: color_data = Z;
		19'b1011010000011111101: color_data = Z;
		19'b1011010000011111110: color_data = Z;
		19'b1011010000011111111: color_data = Z;
		19'b1011010000100000000: color_data = Z;
		19'b1011010000100000001: color_data = Z;
		19'b1011010000100000010: color_data = Z;
		19'b1011010000100000011: color_data = Z;
		19'b1011010000100000100: color_data = Z;
		19'b1011010000100000101: color_data = Z;
		19'b1011010000100000110: color_data = Z;
		19'b1011010000100000111: color_data = Z;
		19'b1011010000100001000: color_data = Z;
		19'b1011010000100001001: color_data = Z;
		19'b1011010000100001010: color_data = Z;
		19'b1011010000100001011: color_data = Z;
		19'b1011010000100001100: color_data = Z;
		19'b1011010000100001101: color_data = Z;
		19'b1011010000100001110: color_data = Z;
		19'b1011010000100001111: color_data = Z;
		19'b1011010000100010000: color_data = Z;
		19'b1011010000100010001: color_data = Z;
		19'b1011010000100010010: color_data = Z;
		19'b1011010000100010011: color_data = Z;
		19'b1011010000100010100: color_data = Z;
		19'b1011010000100010101: color_data = Z;
		19'b1011010000100010110: color_data = Z;
		19'b1011010000100010111: color_data = Z;
		19'b1011010000100011000: color_data = Z;
		19'b1011010000100011001: color_data = Z;
		19'b1011010000100011010: color_data = Z;
		19'b1011010000100011011: color_data = Z;
		19'b1011010000100011100: color_data = Z;
		19'b1011010000100111000: color_data = Z;
		19'b1011010000100111001: color_data = Z;
		19'b1011010000100111010: color_data = Z;
		19'b1011010000100111011: color_data = Z;
		19'b1011010000101000000: color_data = Z;
		19'b1011010000101000011: color_data = Z;
		19'b1011010000101000100: color_data = Z;
		19'b1011010000101000101: color_data = Z;
		19'b1011010000101001110: color_data = Z;
		19'b1011010000101001111: color_data = Z;
		19'b1011010000101010000: color_data = Z;
		19'b1011010000101010001: color_data = Z;
		19'b1011010000101010010: color_data = Z;
		19'b1011010000101010110: color_data = Z;
		19'b1011010000101010111: color_data = Z;
		19'b1011010000101011001: color_data = Z;
		19'b1011010000101011010: color_data = Z;
		19'b1011010000101011011: color_data = Z;
		19'b1011010000101100100: color_data = Z;
		19'b1011010000110000110: color_data = Z;
		19'b1011010000110000111: color_data = Z;
		19'b1011010000110001000: color_data = Z;
		19'b1011010000110001001: color_data = Z;
		19'b1011010000110001010: color_data = Z;
		19'b1011010000110001011: color_data = Z;
		19'b1011010000110001100: color_data = Z;
		19'b1011010000110001101: color_data = Z;
		19'b1011010000110001110: color_data = Z;
		19'b1011010000110001111: color_data = Z;
		19'b1011010000110010000: color_data = Z;
		19'b1011010000110010001: color_data = Z;
		19'b1011010000110010010: color_data = Z;
		19'b1011010000110010011: color_data = Z;
		19'b1011010000110010100: color_data = Z;
		19'b1011010000110010101: color_data = Z;
		19'b1011010000110010110: color_data = Z;
		19'b1011010000110010111: color_data = Z;
		19'b1011010000110011000: color_data = Z;
		19'b1011010000110011001: color_data = Z;
		19'b1011010000110011010: color_data = Z;
		19'b1011010000110011011: color_data = Z;
		19'b1011010000110011100: color_data = Z;
		19'b1011010000110011101: color_data = Z;
		19'b1011010010011101010: color_data = Z;
		19'b1011010010011101011: color_data = Z;
		19'b1011010010011101100: color_data = Z;
		19'b1011010010011101101: color_data = Z;
		19'b1011010010011101110: color_data = Z;
		19'b1011010010011101111: color_data = Z;
		19'b1011010010011110000: color_data = Z;
		19'b1011010010011110001: color_data = Z;
		19'b1011010010011110010: color_data = Z;
		19'b1011010010011110011: color_data = Z;
		19'b1011010010011110100: color_data = Z;
		19'b1011010010011110101: color_data = Z;
		19'b1011010010011110110: color_data = Z;
		19'b1011010010011110111: color_data = Z;
		19'b1011010010011111000: color_data = Z;
		19'b1011010010011111001: color_data = Z;
		19'b1011010010011111010: color_data = Z;
		19'b1011010010011111011: color_data = Z;
		19'b1011010010011111100: color_data = Z;
		19'b1011010010011111101: color_data = Z;
		19'b1011010010011111110: color_data = Z;
		19'b1011010010011111111: color_data = Z;
		19'b1011010010100000000: color_data = Z;
		19'b1011010010100000001: color_data = Z;
		19'b1011010010100000010: color_data = Z;
		19'b1011010010100000011: color_data = Z;
		19'b1011010010100000100: color_data = Z;
		19'b1011010010100000101: color_data = Z;
		19'b1011010010100000110: color_data = Z;
		19'b1011010010100000111: color_data = Z;
		19'b1011010010100001000: color_data = Z;
		19'b1011010010100001001: color_data = Z;
		19'b1011010010100001010: color_data = Z;
		19'b1011010010100001011: color_data = Z;
		19'b1011010010100001100: color_data = Z;
		19'b1011010010100001101: color_data = Z;
		19'b1011010010100001110: color_data = Z;
		19'b1011010010100001111: color_data = Z;
		19'b1011010010100010000: color_data = Z;
		19'b1011010010100010001: color_data = Z;
		19'b1011010010100010010: color_data = Z;
		19'b1011010010100010011: color_data = Z;
		19'b1011010010100010100: color_data = Z;
		19'b1011010010100010101: color_data = Z;
		19'b1011010010100010110: color_data = Z;
		19'b1011010010100010111: color_data = Z;
		19'b1011010010100011000: color_data = Z;
		19'b1011010010100011001: color_data = Z;
		19'b1011010010100011010: color_data = Z;
		19'b1011010010100011011: color_data = Z;
		19'b1011010010100011100: color_data = Z;
		19'b1011010010100011101: color_data = Z;
		19'b1011010010100011110: color_data = Z;
		19'b1011010010100011111: color_data = Z;
		19'b1011010010100111010: color_data = Z;
		19'b1011010010100111011: color_data = Z;
		19'b1011010010101000000: color_data = Z;
		19'b1011010010101000100: color_data = Z;
		19'b1011010010101000101: color_data = Z;
		19'b1011010010101001110: color_data = Z;
		19'b1011010010101001111: color_data = Z;
		19'b1011010010101010000: color_data = Z;
		19'b1011010010101010001: color_data = Z;
		19'b1011010010101010010: color_data = Z;
		19'b1011010010101011001: color_data = Z;
		19'b1011010010101011010: color_data = Z;
		19'b1011010010101011011: color_data = Z;
		19'b1011010010110000011: color_data = Z;
		19'b1011010010110000100: color_data = Z;
		19'b1011010010110000101: color_data = Z;
		19'b1011010010110000110: color_data = Z;
		19'b1011010010110000111: color_data = Z;
		19'b1011010010110001000: color_data = Z;
		19'b1011010010110001001: color_data = Z;
		19'b1011010010110001010: color_data = Z;
		19'b1011010010110001011: color_data = Z;
		19'b1011010010110001100: color_data = Z;
		19'b1011010010110001101: color_data = Z;
		19'b1011010010110001110: color_data = Z;
		19'b1011010010110001111: color_data = Z;
		19'b1011010010110010000: color_data = Z;
		19'b1011010010110010001: color_data = Z;
		19'b1011010010110010010: color_data = Z;
		19'b1011010010110010011: color_data = Z;
		19'b1011010010110010100: color_data = Z;
		19'b1011010010110010101: color_data = Z;
		19'b1011010010110010110: color_data = Z;
		19'b1011010010110010111: color_data = Z;
		19'b1011010010110011000: color_data = Z;
		19'b1011010010110011001: color_data = Z;
		19'b1011010010110011010: color_data = Z;
		19'b1011010010110011011: color_data = Z;
		19'b1011010010110011100: color_data = Z;
		19'b1011010100011101011: color_data = Z;
		19'b1011010100011101100: color_data = Z;
		19'b1011010100011101101: color_data = Z;
		19'b1011010100011101110: color_data = Z;
		19'b1011010100011101111: color_data = Z;
		19'b1011010100011110000: color_data = Z;
		19'b1011010100011110001: color_data = Z;
		19'b1011010100011110010: color_data = Z;
		19'b1011010100011110011: color_data = Z;
		19'b1011010100011110100: color_data = Z;
		19'b1011010100011110101: color_data = Z;
		19'b1011010100011110110: color_data = Z;
		19'b1011010100011110111: color_data = Z;
		19'b1011010100011111000: color_data = Z;
		19'b1011010100011111001: color_data = Z;
		19'b1011010100011111010: color_data = Z;
		19'b1011010100011111011: color_data = Z;
		19'b1011010100011111100: color_data = Z;
		19'b1011010100011111101: color_data = Z;
		19'b1011010100011111110: color_data = Z;
		19'b1011010100011111111: color_data = Z;
		19'b1011010100100000000: color_data = Z;
		19'b1011010100100000001: color_data = Z;
		19'b1011010100100000010: color_data = Z;
		19'b1011010100100000011: color_data = Z;
		19'b1011010100100000100: color_data = Z;
		19'b1011010100100000101: color_data = Z;
		19'b1011010100100000110: color_data = Z;
		19'b1011010100100000111: color_data = Z;
		19'b1011010100100001000: color_data = Z;
		19'b1011010100100001001: color_data = Z;
		19'b1011010100100001010: color_data = Z;
		19'b1011010100100001011: color_data = Z;
		19'b1011010100100001100: color_data = Z;
		19'b1011010100100001101: color_data = Z;
		19'b1011010100100001110: color_data = Z;
		19'b1011010100100001111: color_data = Z;
		19'b1011010100100010000: color_data = Z;
		19'b1011010100100010001: color_data = Z;
		19'b1011010100100010010: color_data = Z;
		19'b1011010100100010011: color_data = Z;
		19'b1011010100100010100: color_data = Z;
		19'b1011010100100010101: color_data = Z;
		19'b1011010100100010110: color_data = Z;
		19'b1011010100100010111: color_data = Z;
		19'b1011010100100011000: color_data = Z;
		19'b1011010100100011001: color_data = Z;
		19'b1011010100100011010: color_data = Z;
		19'b1011010100100011011: color_data = Z;
		19'b1011010100100011100: color_data = Z;
		19'b1011010100100011101: color_data = Z;
		19'b1011010100100011110: color_data = Z;
		19'b1011010100100011111: color_data = Z;
		19'b1011010100100100000: color_data = Z;
		19'b1011010100100100001: color_data = Z;
		19'b1011010100100100010: color_data = Z;
		19'b1011010100100100011: color_data = Z;
		19'b1011010100100111011: color_data = Z;
		19'b1011010100100111111: color_data = Z;
		19'b1011010100101000000: color_data = Z;
		19'b1011010100101000101: color_data = Z;
		19'b1011010100101001110: color_data = Z;
		19'b1011010100101001111: color_data = Z;
		19'b1011010100101010000: color_data = Z;
		19'b1011010100101010001: color_data = Z;
		19'b1011010100101010010: color_data = Z;
		19'b1011010100101011001: color_data = Z;
		19'b1011010100101011010: color_data = Z;
		19'b1011010100101011011: color_data = Z;
		19'b1011010100101011100: color_data = Z;
		19'b1011010100110000000: color_data = Z;
		19'b1011010100110000001: color_data = Z;
		19'b1011010100110000010: color_data = Z;
		19'b1011010100110000011: color_data = Z;
		19'b1011010100110000100: color_data = Z;
		19'b1011010100110000101: color_data = Z;
		19'b1011010100110000110: color_data = Z;
		19'b1011010100110000111: color_data = Z;
		19'b1011010100110001000: color_data = Z;
		19'b1011010100110001001: color_data = Z;
		19'b1011010100110001010: color_data = Z;
		19'b1011010100110001011: color_data = Z;
		19'b1011010100110001100: color_data = Z;
		19'b1011010100110001101: color_data = Z;
		19'b1011010100110001110: color_data = Z;
		19'b1011010100110001111: color_data = Z;
		19'b1011010100110010000: color_data = Z;
		19'b1011010100110010001: color_data = Z;
		19'b1011010100110010010: color_data = Z;
		19'b1011010100110010011: color_data = Z;
		19'b1011010100110010100: color_data = Z;
		19'b1011010100110010101: color_data = Z;
		19'b1011010100110010110: color_data = Z;
		19'b1011010100110010111: color_data = Z;
		19'b1011010100110011000: color_data = Z;
		19'b1011010100110011001: color_data = Z;
		19'b1011010100110011010: color_data = Z;
		19'b1011010100110011011: color_data = Z;
		19'b1011010110011101101: color_data = Z;
		19'b1011010110011101110: color_data = Z;
		19'b1011010110011101111: color_data = Z;
		19'b1011010110011110000: color_data = Z;
		19'b1011010110011110001: color_data = Z;
		19'b1011010110011110010: color_data = Z;
		19'b1011010110011110011: color_data = Z;
		19'b1011010110011110100: color_data = Z;
		19'b1011010110011110101: color_data = Z;
		19'b1011010110011110110: color_data = Z;
		19'b1011010110011110111: color_data = Z;
		19'b1011010110011111000: color_data = Z;
		19'b1011010110011111001: color_data = Z;
		19'b1011010110011111010: color_data = Z;
		19'b1011010110011111011: color_data = Z;
		19'b1011010110011111100: color_data = Z;
		19'b1011010110011111101: color_data = Z;
		19'b1011010110011111110: color_data = Z;
		19'b1011010110011111111: color_data = Z;
		19'b1011010110100000000: color_data = Z;
		19'b1011010110100000001: color_data = Z;
		19'b1011010110100000010: color_data = Z;
		19'b1011010110100000011: color_data = Z;
		19'b1011010110100000100: color_data = Z;
		19'b1011010110100000101: color_data = Z;
		19'b1011010110100000110: color_data = Z;
		19'b1011010110100000111: color_data = Z;
		19'b1011010110100001000: color_data = Z;
		19'b1011010110100001001: color_data = Z;
		19'b1011010110100001010: color_data = Z;
		19'b1011010110100001011: color_data = Z;
		19'b1011010110100001100: color_data = Z;
		19'b1011010110100001101: color_data = Z;
		19'b1011010110100001110: color_data = Z;
		19'b1011010110100001111: color_data = Z;
		19'b1011010110100010000: color_data = Z;
		19'b1011010110100010001: color_data = Z;
		19'b1011010110100010010: color_data = Z;
		19'b1011010110100010011: color_data = Z;
		19'b1011010110100010100: color_data = Z;
		19'b1011010110100010101: color_data = Z;
		19'b1011010110100010110: color_data = Z;
		19'b1011010110100010111: color_data = Z;
		19'b1011010110100011000: color_data = Z;
		19'b1011010110100011001: color_data = Z;
		19'b1011010110100011010: color_data = Z;
		19'b1011010110100011011: color_data = Z;
		19'b1011010110100011100: color_data = Z;
		19'b1011010110100011101: color_data = Z;
		19'b1011010110100011110: color_data = Z;
		19'b1011010110100011111: color_data = Z;
		19'b1011010110100100000: color_data = Z;
		19'b1011010110100100001: color_data = Z;
		19'b1011010110100100010: color_data = Z;
		19'b1011010110100100011: color_data = Z;
		19'b1011010110100100100: color_data = Z;
		19'b1011010110100100101: color_data = Z;
		19'b1011010110100100110: color_data = Z;
		19'b1011010110101000100: color_data = Z;
		19'b1011010110101000101: color_data = Z;
		19'b1011010110101001110: color_data = Z;
		19'b1011010110101001111: color_data = Z;
		19'b1011010110101010000: color_data = Z;
		19'b1011010110101010001: color_data = Z;
		19'b1011010110101011001: color_data = Z;
		19'b1011010110101011010: color_data = Z;
		19'b1011010110101011011: color_data = Z;
		19'b1011010110101011100: color_data = Z;
		19'b1011010110101111101: color_data = Z;
		19'b1011010110101111110: color_data = Z;
		19'b1011010110101111111: color_data = Z;
		19'b1011010110110000000: color_data = Z;
		19'b1011010110110000001: color_data = Z;
		19'b1011010110110000010: color_data = Z;
		19'b1011010110110000011: color_data = Z;
		19'b1011010110110000100: color_data = Z;
		19'b1011010110110000101: color_data = Z;
		19'b1011010110110000110: color_data = Z;
		19'b1011010110110000111: color_data = Z;
		19'b1011010110110001000: color_data = Z;
		19'b1011010110110001001: color_data = Z;
		19'b1011010110110001010: color_data = Z;
		19'b1011010110110001011: color_data = Z;
		19'b1011010110110001100: color_data = Z;
		19'b1011010110110001101: color_data = Z;
		19'b1011010110110001110: color_data = Z;
		19'b1011010110110001111: color_data = Z;
		19'b1011010110110010000: color_data = Z;
		19'b1011010110110010001: color_data = Z;
		19'b1011010110110010010: color_data = Z;
		19'b1011010110110010011: color_data = Z;
		19'b1011010110110010100: color_data = Z;
		19'b1011010110110010101: color_data = Z;
		19'b1011010110110010110: color_data = Z;
		19'b1011010110110010111: color_data = Z;
		19'b1011010110110011000: color_data = Z;
		19'b1011010110110011001: color_data = Z;
		19'b1011010110110011010: color_data = Z;
		19'b1011011000011101110: color_data = Z;
		19'b1011011000011101111: color_data = Z;
		19'b1011011000011110000: color_data = Z;
		19'b1011011000011110001: color_data = Z;
		19'b1011011000011110010: color_data = Z;
		19'b1011011000011110011: color_data = Z;
		19'b1011011000011110100: color_data = Z;
		19'b1011011000011110101: color_data = Z;
		19'b1011011000011110110: color_data = Z;
		19'b1011011000011110111: color_data = Z;
		19'b1011011000011111000: color_data = Z;
		19'b1011011000011111001: color_data = Z;
		19'b1011011000011111010: color_data = Z;
		19'b1011011000011111011: color_data = Z;
		19'b1011011000011111100: color_data = Z;
		19'b1011011000011111101: color_data = Z;
		19'b1011011000011111110: color_data = Z;
		19'b1011011000011111111: color_data = Z;
		19'b1011011000100000000: color_data = Z;
		19'b1011011000100000001: color_data = Z;
		19'b1011011000100000010: color_data = Z;
		19'b1011011000100000011: color_data = Z;
		19'b1011011000100000100: color_data = Z;
		19'b1011011000100000101: color_data = Z;
		19'b1011011000100000110: color_data = Z;
		19'b1011011000100000111: color_data = Z;
		19'b1011011000100001000: color_data = Z;
		19'b1011011000100001001: color_data = Z;
		19'b1011011000100001010: color_data = Z;
		19'b1011011000100001011: color_data = Z;
		19'b1011011000100001100: color_data = Z;
		19'b1011011000100001101: color_data = Z;
		19'b1011011000100001110: color_data = Z;
		19'b1011011000100001111: color_data = Z;
		19'b1011011000100010000: color_data = Z;
		19'b1011011000100010001: color_data = Z;
		19'b1011011000100010010: color_data = Z;
		19'b1011011000100010011: color_data = Z;
		19'b1011011000100010100: color_data = Z;
		19'b1011011000100010101: color_data = Z;
		19'b1011011000100010110: color_data = Z;
		19'b1011011000100010111: color_data = Z;
		19'b1011011000100011000: color_data = Z;
		19'b1011011000100011001: color_data = Z;
		19'b1011011000100011010: color_data = Z;
		19'b1011011000100011011: color_data = Z;
		19'b1011011000100011100: color_data = Z;
		19'b1011011000100011101: color_data = Z;
		19'b1011011000100011110: color_data = Z;
		19'b1011011000100011111: color_data = Z;
		19'b1011011000100100000: color_data = Z;
		19'b1011011000100100001: color_data = Z;
		19'b1011011000100100010: color_data = Z;
		19'b1011011000100100011: color_data = Z;
		19'b1011011000100100100: color_data = Z;
		19'b1011011000100100101: color_data = Z;
		19'b1011011000100100110: color_data = Z;
		19'b1011011000100100111: color_data = Z;
		19'b1011011000100101000: color_data = Z;
		19'b1011011000100101001: color_data = Z;
		19'b1011011000101011010: color_data = Z;
		19'b1011011000101011011: color_data = Z;
		19'b1011011000101111010: color_data = Z;
		19'b1011011000101111011: color_data = Z;
		19'b1011011000101111100: color_data = Z;
		19'b1011011000101111101: color_data = Z;
		19'b1011011000101111110: color_data = Z;
		19'b1011011000101111111: color_data = Z;
		19'b1011011000110000000: color_data = Z;
		19'b1011011000110000001: color_data = Z;
		19'b1011011000110000010: color_data = Z;
		19'b1011011000110000011: color_data = Z;
		19'b1011011000110000100: color_data = Z;
		19'b1011011000110000101: color_data = Z;
		19'b1011011000110000110: color_data = Z;
		19'b1011011000110000111: color_data = Z;
		19'b1011011000110001000: color_data = Z;
		19'b1011011000110001001: color_data = Z;
		19'b1011011000110001010: color_data = Z;
		19'b1011011000110001011: color_data = Z;
		19'b1011011000110001100: color_data = Z;
		19'b1011011000110001101: color_data = Z;
		19'b1011011000110001110: color_data = Z;
		19'b1011011000110001111: color_data = Z;
		19'b1011011000110010000: color_data = Z;
		19'b1011011000110010001: color_data = Z;
		19'b1011011000110010010: color_data = Z;
		19'b1011011000110010011: color_data = Z;
		19'b1011011000110010100: color_data = Z;
		19'b1011011000110010101: color_data = Z;
		19'b1011011000110010110: color_data = Z;
		19'b1011011000110010111: color_data = Z;
		19'b1011011000110011000: color_data = Z;
		19'b1011011000110011001: color_data = Z;
		19'b1011011010011101111: color_data = Z;
		19'b1011011010011110000: color_data = Z;
		19'b1011011010011110001: color_data = Z;
		19'b1011011010011110010: color_data = Z;
		19'b1011011010011110011: color_data = Z;
		19'b1011011010011110100: color_data = Z;
		19'b1011011010011110101: color_data = Z;
		19'b1011011010011110110: color_data = Z;
		19'b1011011010011110111: color_data = Z;
		19'b1011011010011111000: color_data = Z;
		19'b1011011010011111001: color_data = Z;
		19'b1011011010011111010: color_data = Z;
		19'b1011011010011111011: color_data = Z;
		19'b1011011010011111100: color_data = Z;
		19'b1011011010011111101: color_data = Z;
		19'b1011011010011111110: color_data = Z;
		19'b1011011010011111111: color_data = Z;
		19'b1011011010100000000: color_data = Z;
		19'b1011011010100000001: color_data = Z;
		19'b1011011010100000010: color_data = Z;
		19'b1011011010100000011: color_data = Z;
		19'b1011011010100000100: color_data = Z;
		19'b1011011010100000101: color_data = Z;
		19'b1011011010100000110: color_data = Z;
		19'b1011011010100000111: color_data = Z;
		19'b1011011010100001000: color_data = Z;
		19'b1011011010100001001: color_data = Z;
		19'b1011011010100001010: color_data = Z;
		19'b1011011010100001011: color_data = Z;
		19'b1011011010100001100: color_data = Z;
		19'b1011011010100001101: color_data = Z;
		19'b1011011010100001110: color_data = Z;
		19'b1011011010100001111: color_data = Z;
		19'b1011011010100010000: color_data = Z;
		19'b1011011010100010001: color_data = Z;
		19'b1011011010100010010: color_data = Z;
		19'b1011011010100010011: color_data = Z;
		19'b1011011010100010100: color_data = Z;
		19'b1011011010100010101: color_data = Z;
		19'b1011011010100010110: color_data = Z;
		19'b1011011010100010111: color_data = Z;
		19'b1011011010100011000: color_data = Z;
		19'b1011011010100011001: color_data = Z;
		19'b1011011010100011010: color_data = Z;
		19'b1011011010100011011: color_data = Z;
		19'b1011011010100011100: color_data = Z;
		19'b1011011010100011101: color_data = Z;
		19'b1011011010100011110: color_data = Z;
		19'b1011011010100011111: color_data = Z;
		19'b1011011010100100000: color_data = Z;
		19'b1011011010100100001: color_data = Z;
		19'b1011011010100100010: color_data = Z;
		19'b1011011010100100011: color_data = Z;
		19'b1011011010100100100: color_data = Z;
		19'b1011011010100100101: color_data = Z;
		19'b1011011010100100110: color_data = Z;
		19'b1011011010100100111: color_data = Z;
		19'b1011011010100101000: color_data = Z;
		19'b1011011010100101001: color_data = Z;
		19'b1011011010100101010: color_data = Z;
		19'b1011011010101111000: color_data = Z;
		19'b1011011010101111001: color_data = Z;
		19'b1011011010101111010: color_data = Z;
		19'b1011011010101111011: color_data = Z;
		19'b1011011010101111100: color_data = Z;
		19'b1011011010101111101: color_data = Z;
		19'b1011011010101111110: color_data = Z;
		19'b1011011010101111111: color_data = Z;
		19'b1011011010110000000: color_data = Z;
		19'b1011011010110000001: color_data = Z;
		19'b1011011010110000010: color_data = Z;
		19'b1011011010110000011: color_data = Z;
		19'b1011011010110000100: color_data = Z;
		19'b1011011010110000101: color_data = Z;
		19'b1011011010110000110: color_data = Z;
		19'b1011011010110000111: color_data = Z;
		19'b1011011010110001000: color_data = Z;
		19'b1011011010110001001: color_data = Z;
		19'b1011011010110001010: color_data = Z;
		19'b1011011010110001011: color_data = Z;
		19'b1011011010110001100: color_data = Z;
		19'b1011011010110001101: color_data = Z;
		19'b1011011010110001110: color_data = Z;
		19'b1011011010110001111: color_data = Z;
		19'b1011011010110010000: color_data = Z;
		19'b1011011010110010001: color_data = Z;
		19'b1011011010110010010: color_data = Z;
		19'b1011011010110010011: color_data = Z;
		19'b1011011010110010100: color_data = Z;
		19'b1011011010110010101: color_data = Z;
		19'b1011011010110010110: color_data = Z;
		19'b1011011010110010111: color_data = Z;
		19'b1011011010110011000: color_data = Z;
		19'b1011011100011110000: color_data = Z;
		19'b1011011100011110001: color_data = Z;
		19'b1011011100011110010: color_data = Z;
		19'b1011011100011110011: color_data = Z;
		19'b1011011100011110100: color_data = Z;
		19'b1011011100011110101: color_data = Z;
		19'b1011011100011110110: color_data = Z;
		19'b1011011100011110111: color_data = Z;
		19'b1011011100011111000: color_data = Z;
		19'b1011011100011111001: color_data = Z;
		19'b1011011100011111010: color_data = Z;
		19'b1011011100011111011: color_data = Z;
		19'b1011011100011111100: color_data = Z;
		19'b1011011100011111101: color_data = Z;
		19'b1011011100011111110: color_data = Z;
		19'b1011011100011111111: color_data = Z;
		19'b1011011100100000000: color_data = Z;
		19'b1011011100100000001: color_data = Z;
		19'b1011011100100000010: color_data = Z;
		19'b1011011100100000011: color_data = Z;
		19'b1011011100100000100: color_data = Z;
		19'b1011011100100000101: color_data = Z;
		19'b1011011100100000110: color_data = Z;
		19'b1011011100100000111: color_data = Z;
		19'b1011011100100001000: color_data = Z;
		19'b1011011100100001001: color_data = Z;
		19'b1011011100100001010: color_data = Z;
		19'b1011011100100001011: color_data = Z;
		19'b1011011100100001100: color_data = Z;
		19'b1011011100100001101: color_data = Z;
		19'b1011011100100001110: color_data = Z;
		19'b1011011100100001111: color_data = Z;
		19'b1011011100100010000: color_data = Z;
		19'b1011011100100010001: color_data = Z;
		19'b1011011100100010010: color_data = Z;
		19'b1011011100100010011: color_data = Z;
		19'b1011011100100010100: color_data = Z;
		19'b1011011100100010101: color_data = Z;
		19'b1011011100100010110: color_data = Z;
		19'b1011011100100010111: color_data = Z;
		19'b1011011100100011000: color_data = Z;
		19'b1011011100100011001: color_data = Z;
		19'b1011011100100011010: color_data = Z;
		19'b1011011100100011011: color_data = Z;
		19'b1011011100100011100: color_data = Z;
		19'b1011011100100011101: color_data = Z;
		19'b1011011100100011110: color_data = Z;
		19'b1011011100100011111: color_data = Z;
		19'b1011011100100100000: color_data = Z;
		19'b1011011100100100001: color_data = Z;
		19'b1011011100100100010: color_data = Z;
		19'b1011011100100100011: color_data = Z;
		19'b1011011100100100100: color_data = Z;
		19'b1011011100100100101: color_data = Z;
		19'b1011011100100100110: color_data = Z;
		19'b1011011100100100111: color_data = Z;
		19'b1011011100100101000: color_data = Z;
		19'b1011011100100101001: color_data = Z;
		19'b1011011100100101010: color_data = Z;
		19'b1011011100100101011: color_data = Z;
		19'b1011011100100101100: color_data = Z;
		19'b1011011100100101101: color_data = Z;
		19'b1011011100101110110: color_data = Z;
		19'b1011011100101110111: color_data = Z;
		19'b1011011100101111000: color_data = Z;
		19'b1011011100101111001: color_data = Z;
		19'b1011011100101111010: color_data = Z;
		19'b1011011100101111011: color_data = Z;
		19'b1011011100101111100: color_data = Z;
		19'b1011011100101111101: color_data = Z;
		19'b1011011100101111110: color_data = Z;
		19'b1011011100101111111: color_data = Z;
		19'b1011011100110000000: color_data = Z;
		19'b1011011100110000001: color_data = Z;
		19'b1011011100110000010: color_data = Z;
		19'b1011011100110000011: color_data = Z;
		19'b1011011100110000100: color_data = Z;
		19'b1011011100110000101: color_data = Z;
		19'b1011011100110000110: color_data = Z;
		19'b1011011100110000111: color_data = Z;
		19'b1011011100110001000: color_data = Z;
		19'b1011011100110001001: color_data = Z;
		19'b1011011100110001010: color_data = Z;
		19'b1011011100110001011: color_data = Z;
		19'b1011011100110001100: color_data = Z;
		19'b1011011100110001101: color_data = Z;
		19'b1011011100110001110: color_data = Z;
		19'b1011011100110001111: color_data = Z;
		19'b1011011100110010000: color_data = Z;
		19'b1011011100110010001: color_data = Z;
		19'b1011011100110010010: color_data = Z;
		19'b1011011100110010011: color_data = Z;
		19'b1011011100110010100: color_data = Z;
		19'b1011011100110010101: color_data = Z;
		19'b1011011100110010110: color_data = Z;
		19'b1011011100110010111: color_data = Z;
		19'b1011011110011110010: color_data = Z;
		19'b1011011110011110011: color_data = Z;
		19'b1011011110011110100: color_data = Z;
		19'b1011011110011110101: color_data = Z;
		19'b1011011110011110110: color_data = Z;
		19'b1011011110011110111: color_data = Z;
		19'b1011011110011111000: color_data = Z;
		19'b1011011110011111001: color_data = Z;
		19'b1011011110011111010: color_data = Z;
		19'b1011011110011111011: color_data = Z;
		19'b1011011110011111100: color_data = Z;
		19'b1011011110011111101: color_data = Z;
		19'b1011011110011111110: color_data = Z;
		19'b1011011110011111111: color_data = Z;
		19'b1011011110100000000: color_data = Z;
		19'b1011011110100000001: color_data = Z;
		19'b1011011110100000010: color_data = Z;
		19'b1011011110100000011: color_data = Z;
		19'b1011011110100000100: color_data = Z;
		19'b1011011110100000101: color_data = Z;
		19'b1011011110100000110: color_data = Z;
		19'b1011011110100000111: color_data = Z;
		19'b1011011110100001000: color_data = Z;
		19'b1011011110100001001: color_data = Z;
		19'b1011011110100001010: color_data = Z;
		19'b1011011110100001011: color_data = Z;
		19'b1011011110100001100: color_data = Z;
		19'b1011011110100001101: color_data = Z;
		19'b1011011110100001110: color_data = Z;
		19'b1011011110100001111: color_data = Z;
		19'b1011011110100010000: color_data = Z;
		19'b1011011110100010001: color_data = Z;
		19'b1011011110100010010: color_data = Z;
		19'b1011011110100010011: color_data = Z;
		19'b1011011110100010100: color_data = Z;
		19'b1011011110100010101: color_data = Z;
		19'b1011011110100010110: color_data = Z;
		19'b1011011110100010111: color_data = Z;
		19'b1011011110100011000: color_data = Z;
		19'b1011011110100011001: color_data = Z;
		19'b1011011110100011010: color_data = Z;
		19'b1011011110100011011: color_data = Z;
		19'b1011011110100011100: color_data = Z;
		19'b1011011110100011101: color_data = Z;
		19'b1011011110100011110: color_data = Z;
		19'b1011011110100011111: color_data = Z;
		19'b1011011110100100000: color_data = Z;
		19'b1011011110100100001: color_data = Z;
		19'b1011011110100100010: color_data = Z;
		19'b1011011110100100011: color_data = Z;
		19'b1011011110100100100: color_data = Z;
		19'b1011011110100100101: color_data = Z;
		19'b1011011110100100110: color_data = Z;
		19'b1011011110100100111: color_data = Z;
		19'b1011011110100101000: color_data = Z;
		19'b1011011110100101001: color_data = Z;
		19'b1011011110100101010: color_data = Z;
		19'b1011011110100101011: color_data = Z;
		19'b1011011110100101100: color_data = Z;
		19'b1011011110100101101: color_data = Z;
		19'b1011011110100101110: color_data = Z;
		19'b1011011110100101111: color_data = Z;
		19'b1011011110100110000: color_data = Z;
		19'b1011011110100110011: color_data = Z;
		19'b1011011110101110100: color_data = Z;
		19'b1011011110101110101: color_data = Z;
		19'b1011011110101110110: color_data = Z;
		19'b1011011110101110111: color_data = Z;
		19'b1011011110101111000: color_data = Z;
		19'b1011011110101111001: color_data = Z;
		19'b1011011110101111010: color_data = Z;
		19'b1011011110101111011: color_data = Z;
		19'b1011011110101111100: color_data = Z;
		19'b1011011110101111101: color_data = Z;
		19'b1011011110101111110: color_data = Z;
		19'b1011011110101111111: color_data = Z;
		19'b1011011110110000000: color_data = Z;
		19'b1011011110110000001: color_data = Z;
		19'b1011011110110000010: color_data = Z;
		19'b1011011110110000011: color_data = Z;
		19'b1011011110110000100: color_data = Z;
		19'b1011011110110000101: color_data = Z;
		19'b1011011110110000110: color_data = Z;
		19'b1011011110110000111: color_data = Z;
		19'b1011011110110001000: color_data = Z;
		19'b1011011110110001001: color_data = Z;
		19'b1011011110110001010: color_data = Z;
		19'b1011011110110001011: color_data = Z;
		19'b1011011110110001100: color_data = Z;
		19'b1011011110110001101: color_data = Z;
		19'b1011011110110001110: color_data = Z;
		19'b1011011110110001111: color_data = Z;
		19'b1011011110110010000: color_data = Z;
		19'b1011011110110010001: color_data = Z;
		19'b1011011110110010010: color_data = Z;
		19'b1011011110110010011: color_data = Z;
		19'b1011011110110010100: color_data = Z;
		19'b1011011110110010101: color_data = Z;
		19'b1011011110110010110: color_data = Z;
		19'b1011100000011110011: color_data = Z;
		19'b1011100000011110100: color_data = Z;
		19'b1011100000011110101: color_data = Z;
		19'b1011100000011110110: color_data = Z;
		19'b1011100000011110111: color_data = Z;
		19'b1011100000011111000: color_data = Z;
		19'b1011100000011111001: color_data = Z;
		19'b1011100000011111010: color_data = Z;
		19'b1011100000011111011: color_data = Z;
		19'b1011100000011111100: color_data = Z;
		19'b1011100000011111101: color_data = Z;
		19'b1011100000011111110: color_data = Z;
		19'b1011100000011111111: color_data = Z;
		19'b1011100000100000000: color_data = Z;
		19'b1011100000100000001: color_data = Z;
		19'b1011100000100000010: color_data = Z;
		19'b1011100000100000011: color_data = Z;
		19'b1011100000100000100: color_data = Z;
		19'b1011100000100000101: color_data = Z;
		19'b1011100000100000110: color_data = Z;
		19'b1011100000100000111: color_data = Z;
		19'b1011100000100001000: color_data = Z;
		19'b1011100000100001001: color_data = Z;
		19'b1011100000100001010: color_data = Z;
		19'b1011100000100001011: color_data = Z;
		19'b1011100000100001100: color_data = Z;
		19'b1011100000100001101: color_data = Z;
		19'b1011100000100001110: color_data = Z;
		19'b1011100000100001111: color_data = Z;
		19'b1011100000100010000: color_data = Z;
		19'b1011100000100010001: color_data = Z;
		19'b1011100000100010010: color_data = Z;
		19'b1011100000100010011: color_data = Z;
		19'b1011100000100010100: color_data = Z;
		19'b1011100000100010101: color_data = Z;
		19'b1011100000100010110: color_data = Z;
		19'b1011100000100010111: color_data = Z;
		19'b1011100000100011000: color_data = Z;
		19'b1011100000100011001: color_data = Z;
		19'b1011100000100011010: color_data = Z;
		19'b1011100000100011011: color_data = Z;
		19'b1011100000100011100: color_data = Z;
		19'b1011100000100011101: color_data = Z;
		19'b1011100000100011110: color_data = Z;
		19'b1011100000100011111: color_data = Z;
		19'b1011100000100100000: color_data = Z;
		19'b1011100000100100001: color_data = Z;
		19'b1011100000100100010: color_data = Z;
		19'b1011100000100100011: color_data = Z;
		19'b1011100000100100100: color_data = Z;
		19'b1011100000100100101: color_data = Z;
		19'b1011100000100100110: color_data = Z;
		19'b1011100000100100111: color_data = Z;
		19'b1011100000100101000: color_data = Z;
		19'b1011100000100101001: color_data = Z;
		19'b1011100000100101010: color_data = Z;
		19'b1011100000100101011: color_data = Z;
		19'b1011100000100101100: color_data = Z;
		19'b1011100000100101101: color_data = Z;
		19'b1011100000100101110: color_data = Z;
		19'b1011100000100101111: color_data = Z;
		19'b1011100000100110000: color_data = Z;
		19'b1011100000100110001: color_data = Z;
		19'b1011100000100110010: color_data = Z;
		19'b1011100000100110011: color_data = Z;
		19'b1011100000100110100: color_data = Z;
		19'b1011100000100110101: color_data = Z;
		19'b1011100000101110001: color_data = Z;
		19'b1011100000101110010: color_data = Z;
		19'b1011100000101110011: color_data = Z;
		19'b1011100000101110100: color_data = Z;
		19'b1011100000101110101: color_data = Z;
		19'b1011100000101110110: color_data = Z;
		19'b1011100000101110111: color_data = Z;
		19'b1011100000101111000: color_data = Z;
		19'b1011100000101111001: color_data = Z;
		19'b1011100000101111010: color_data = Z;
		19'b1011100000101111011: color_data = Z;
		19'b1011100000101111100: color_data = Z;
		19'b1011100000101111101: color_data = Z;
		19'b1011100000101111110: color_data = Z;
		19'b1011100000101111111: color_data = Z;
		19'b1011100000110000000: color_data = Z;
		19'b1011100000110000001: color_data = Z;
		19'b1011100000110000010: color_data = Z;
		19'b1011100000110000011: color_data = Z;
		19'b1011100000110000100: color_data = Z;
		19'b1011100000110000101: color_data = Z;
		19'b1011100000110000110: color_data = Z;
		19'b1011100000110000111: color_data = Z;
		19'b1011100000110001000: color_data = Z;
		19'b1011100000110001001: color_data = Z;
		19'b1011100000110001010: color_data = Z;
		19'b1011100000110001011: color_data = Z;
		19'b1011100000110001100: color_data = Z;
		19'b1011100000110001101: color_data = Z;
		19'b1011100000110001110: color_data = Z;
		19'b1011100000110001111: color_data = Z;
		19'b1011100000110010000: color_data = Z;
		19'b1011100000110010001: color_data = Z;
		19'b1011100000110010010: color_data = Z;
		19'b1011100000110010011: color_data = Z;
		19'b1011100000110010100: color_data = Z;
		19'b1011100000110010101: color_data = Z;
		19'b1011100010011110100: color_data = Z;
		19'b1011100010011110101: color_data = Z;
		19'b1011100010011110110: color_data = Z;
		19'b1011100010011110111: color_data = Z;
		19'b1011100010011111000: color_data = Z;
		19'b1011100010011111001: color_data = Z;
		19'b1011100010011111010: color_data = Z;
		19'b1011100010011111011: color_data = Z;
		19'b1011100010011111100: color_data = Z;
		19'b1011100010011111101: color_data = Z;
		19'b1011100010011111110: color_data = Z;
		19'b1011100010011111111: color_data = Z;
		19'b1011100010100000000: color_data = Z;
		19'b1011100010100000001: color_data = Z;
		19'b1011100010100000010: color_data = Z;
		19'b1011100010100000011: color_data = Z;
		19'b1011100010100000100: color_data = Z;
		19'b1011100010100000101: color_data = Z;
		19'b1011100010100000110: color_data = Z;
		19'b1011100010100000111: color_data = Z;
		19'b1011100010100001000: color_data = Z;
		19'b1011100010100001001: color_data = Z;
		19'b1011100010100001010: color_data = Z;
		19'b1011100010100001011: color_data = Z;
		19'b1011100010100001100: color_data = Z;
		19'b1011100010100001101: color_data = Z;
		19'b1011100010100001110: color_data = Z;
		19'b1011100010100001111: color_data = Z;
		19'b1011100010100010000: color_data = Z;
		19'b1011100010100010001: color_data = Z;
		19'b1011100010100010010: color_data = Z;
		19'b1011100010100010011: color_data = Z;
		19'b1011100010100010100: color_data = Z;
		19'b1011100010100010101: color_data = Z;
		19'b1011100010100010110: color_data = Z;
		19'b1011100010100010111: color_data = Z;
		19'b1011100010100011000: color_data = Z;
		19'b1011100010100011001: color_data = Z;
		19'b1011100010100011010: color_data = Z;
		19'b1011100010100011011: color_data = Z;
		19'b1011100010100011100: color_data = Z;
		19'b1011100010100011101: color_data = Z;
		19'b1011100010100011110: color_data = Z;
		19'b1011100010100011111: color_data = Z;
		19'b1011100010100100000: color_data = Z;
		19'b1011100010100100001: color_data = Z;
		19'b1011100010100100010: color_data = Z;
		19'b1011100010100100011: color_data = Z;
		19'b1011100010100100100: color_data = Z;
		19'b1011100010100100101: color_data = Z;
		19'b1011100010100100110: color_data = Z;
		19'b1011100010100100111: color_data = Z;
		19'b1011100010100101000: color_data = Z;
		19'b1011100010100101001: color_data = Z;
		19'b1011100010100101010: color_data = Z;
		19'b1011100010100101011: color_data = Z;
		19'b1011100010100101100: color_data = Z;
		19'b1011100010100101101: color_data = Z;
		19'b1011100010100101110: color_data = Z;
		19'b1011100010100101111: color_data = Z;
		19'b1011100010100110000: color_data = Z;
		19'b1011100010100110001: color_data = Z;
		19'b1011100010100110010: color_data = Z;
		19'b1011100010100110011: color_data = Z;
		19'b1011100010100110100: color_data = Z;
		19'b1011100010100110101: color_data = Z;
		19'b1011100010100110110: color_data = Z;
		19'b1011100010100110111: color_data = Z;
		19'b1011100010101101010: color_data = Z;
		19'b1011100010101101011: color_data = Z;
		19'b1011100010101101100: color_data = Z;
		19'b1011100010101101101: color_data = Z;
		19'b1011100010101101110: color_data = Z;
		19'b1011100010101101111: color_data = Z;
		19'b1011100010101110000: color_data = Z;
		19'b1011100010101110001: color_data = Z;
		19'b1011100010101110010: color_data = Z;
		19'b1011100010101110011: color_data = Z;
		19'b1011100010101110100: color_data = Z;
		19'b1011100010101110101: color_data = Z;
		19'b1011100010101110110: color_data = Z;
		19'b1011100010101110111: color_data = Z;
		19'b1011100010101111000: color_data = Z;
		19'b1011100010101111001: color_data = Z;
		19'b1011100010101111010: color_data = Z;
		19'b1011100010101111011: color_data = Z;
		19'b1011100010101111100: color_data = Z;
		19'b1011100010101111101: color_data = Z;
		19'b1011100010101111110: color_data = Z;
		19'b1011100010101111111: color_data = Z;
		19'b1011100010110000000: color_data = Z;
		19'b1011100010110000001: color_data = Z;
		19'b1011100010110000010: color_data = Z;
		19'b1011100010110000011: color_data = Z;
		19'b1011100010110000100: color_data = Z;
		19'b1011100010110000101: color_data = Z;
		19'b1011100010110000110: color_data = Z;
		19'b1011100010110000111: color_data = Z;
		19'b1011100010110001000: color_data = Z;
		19'b1011100010110001001: color_data = Z;
		19'b1011100010110001010: color_data = Z;
		19'b1011100010110001011: color_data = Z;
		19'b1011100010110001100: color_data = Z;
		19'b1011100010110001101: color_data = Z;
		19'b1011100010110001110: color_data = Z;
		19'b1011100010110001111: color_data = Z;
		19'b1011100010110010000: color_data = Z;
		19'b1011100010110010001: color_data = Z;
		19'b1011100010110010010: color_data = Z;
		19'b1011100010110010011: color_data = Z;
		19'b1011100010110010100: color_data = Z;
		19'b1011100100011110110: color_data = Z;
		19'b1011100100011110111: color_data = Z;
		19'b1011100100011111000: color_data = Z;
		19'b1011100100011111001: color_data = Z;
		19'b1011100100011111010: color_data = Z;
		19'b1011100100011111011: color_data = Z;
		19'b1011100100011111100: color_data = Z;
		19'b1011100100011111101: color_data = Z;
		19'b1011100100011111110: color_data = Z;
		19'b1011100100011111111: color_data = Z;
		19'b1011100100100000000: color_data = Z;
		19'b1011100100100000001: color_data = Z;
		19'b1011100100100000010: color_data = Z;
		19'b1011100100100000011: color_data = Z;
		19'b1011100100100000100: color_data = Z;
		19'b1011100100100000101: color_data = Z;
		19'b1011100100100000110: color_data = Z;
		19'b1011100100100000111: color_data = Z;
		19'b1011100100100001000: color_data = Z;
		19'b1011100100100001001: color_data = Z;
		19'b1011100100100001010: color_data = Z;
		19'b1011100100100001011: color_data = Z;
		19'b1011100100100001100: color_data = Z;
		19'b1011100100100001101: color_data = Z;
		19'b1011100100100001110: color_data = Z;
		19'b1011100100100001111: color_data = Z;
		19'b1011100100100010000: color_data = Z;
		19'b1011100100100010001: color_data = Z;
		19'b1011100100100010010: color_data = Z;
		19'b1011100100100010011: color_data = Z;
		19'b1011100100100010100: color_data = Z;
		19'b1011100100100010101: color_data = Z;
		19'b1011100100100010110: color_data = Z;
		19'b1011100100100010111: color_data = Z;
		19'b1011100100100011000: color_data = Z;
		19'b1011100100100011001: color_data = Z;
		19'b1011100100100011010: color_data = Z;
		19'b1011100100100011011: color_data = Z;
		19'b1011100100100011100: color_data = Z;
		19'b1011100100100011101: color_data = Z;
		19'b1011100100100011110: color_data = Z;
		19'b1011100100100011111: color_data = Z;
		19'b1011100100100100000: color_data = Z;
		19'b1011100100100100001: color_data = Z;
		19'b1011100100100100010: color_data = Z;
		19'b1011100100100100011: color_data = Z;
		19'b1011100100100100100: color_data = Z;
		19'b1011100100100100101: color_data = Z;
		19'b1011100100100100110: color_data = Z;
		19'b1011100100100100111: color_data = Z;
		19'b1011100100100101000: color_data = Z;
		19'b1011100100100101001: color_data = Z;
		19'b1011100100100101010: color_data = Z;
		19'b1011100100100101011: color_data = Z;
		19'b1011100100100101100: color_data = Z;
		19'b1011100100100101101: color_data = Z;
		19'b1011100100100101110: color_data = Z;
		19'b1011100100100101111: color_data = Z;
		19'b1011100100100110000: color_data = Z;
		19'b1011100100100110001: color_data = Z;
		19'b1011100100100110010: color_data = Z;
		19'b1011100100100110011: color_data = Z;
		19'b1011100100100110100: color_data = Z;
		19'b1011100100100110101: color_data = Z;
		19'b1011100100100110110: color_data = Z;
		19'b1011100100100110111: color_data = Z;
		19'b1011100100100111000: color_data = Z;
		19'b1011100100101100001: color_data = Z;
		19'b1011100100101100010: color_data = Z;
		19'b1011100100101100011: color_data = Z;
		19'b1011100100101100100: color_data = Z;
		19'b1011100100101100101: color_data = Z;
		19'b1011100100101100110: color_data = Z;
		19'b1011100100101100111: color_data = Z;
		19'b1011100100101101000: color_data = Z;
		19'b1011100100101101001: color_data = Z;
		19'b1011100100101101010: color_data = Z;
		19'b1011100100101101011: color_data = Z;
		19'b1011100100101101100: color_data = Z;
		19'b1011100100101101101: color_data = Z;
		19'b1011100100101101110: color_data = Z;
		19'b1011100100101101111: color_data = Z;
		19'b1011100100101110000: color_data = Z;
		19'b1011100100101110001: color_data = Z;
		19'b1011100100101110010: color_data = Z;
		19'b1011100100101110011: color_data = Z;
		19'b1011100100101110100: color_data = Z;
		19'b1011100100101110101: color_data = Z;
		19'b1011100100101110110: color_data = Z;
		19'b1011100100101110111: color_data = Z;
		19'b1011100100101111000: color_data = Z;
		19'b1011100100101111001: color_data = Z;
		19'b1011100100101111010: color_data = Z;
		19'b1011100100101111011: color_data = Z;
		19'b1011100100101111100: color_data = Z;
		19'b1011100100101111101: color_data = Z;
		19'b1011100100101111110: color_data = Z;
		19'b1011100100101111111: color_data = Z;
		19'b1011100100110000000: color_data = Z;
		19'b1011100100110000001: color_data = Z;
		19'b1011100100110000010: color_data = Z;
		19'b1011100100110000011: color_data = Z;
		19'b1011100100110000100: color_data = Z;
		19'b1011100100110000101: color_data = Z;
		19'b1011100100110000110: color_data = Z;
		19'b1011100100110000111: color_data = Z;
		19'b1011100100110001000: color_data = Z;
		19'b1011100100110001001: color_data = Z;
		19'b1011100100110001010: color_data = Z;
		19'b1011100100110001011: color_data = Z;
		19'b1011100100110001100: color_data = Z;
		19'b1011100100110001101: color_data = Z;
		19'b1011100100110001110: color_data = Z;
		19'b1011100100110001111: color_data = Z;
		19'b1011100100110010000: color_data = Z;
		19'b1011100100110010001: color_data = Z;
		19'b1011100100110010010: color_data = Z;
		19'b1011100100110010011: color_data = Z;
		19'b1011100110011111000: color_data = Z;
		19'b1011100110011111001: color_data = Z;
		19'b1011100110011111010: color_data = Z;
		19'b1011100110011111011: color_data = Z;
		19'b1011100110011111100: color_data = Z;
		19'b1011100110011111101: color_data = Z;
		19'b1011100110011111110: color_data = Z;
		19'b1011100110011111111: color_data = Z;
		19'b1011100110100000000: color_data = Z;
		19'b1011100110100000001: color_data = Z;
		19'b1011100110100000010: color_data = Z;
		19'b1011100110100000011: color_data = Z;
		19'b1011100110100000100: color_data = Z;
		19'b1011100110100000101: color_data = Z;
		19'b1011100110100000110: color_data = Z;
		19'b1011100110100000111: color_data = Z;
		19'b1011100110100001000: color_data = Z;
		19'b1011100110100001001: color_data = Z;
		19'b1011100110100001010: color_data = Z;
		19'b1011100110100001011: color_data = Z;
		19'b1011100110100001100: color_data = Z;
		19'b1011100110100001101: color_data = Z;
		19'b1011100110100001110: color_data = Z;
		19'b1011100110100001111: color_data = Z;
		19'b1011100110100010000: color_data = Z;
		19'b1011100110100010001: color_data = Z;
		19'b1011100110100010010: color_data = Z;
		19'b1011100110100010011: color_data = Z;
		19'b1011100110100010100: color_data = Z;
		19'b1011100110100010101: color_data = Z;
		19'b1011100110100010110: color_data = Z;
		19'b1011100110100010111: color_data = Z;
		19'b1011100110100011000: color_data = Z;
		19'b1011100110100011001: color_data = Z;
		19'b1011100110100011010: color_data = Z;
		19'b1011100110100011011: color_data = Z;
		19'b1011100110100011100: color_data = Z;
		19'b1011100110100011101: color_data = Z;
		19'b1011100110100011110: color_data = Z;
		19'b1011100110100011111: color_data = Z;
		19'b1011100110100100000: color_data = Z;
		19'b1011100110100100001: color_data = Z;
		19'b1011100110100100010: color_data = Z;
		19'b1011100110100100011: color_data = Z;
		19'b1011100110100100100: color_data = Z;
		19'b1011100110100100101: color_data = Z;
		19'b1011100110100100110: color_data = Z;
		19'b1011100110100100111: color_data = Z;
		19'b1011100110100101000: color_data = Z;
		19'b1011100110100101001: color_data = Z;
		19'b1011100110100101010: color_data = Z;
		19'b1011100110100101011: color_data = Z;
		19'b1011100110100101100: color_data = Z;
		19'b1011100110100101101: color_data = Z;
		19'b1011100110100101110: color_data = Z;
		19'b1011100110100101111: color_data = Z;
		19'b1011100110100110000: color_data = Z;
		19'b1011100110100110001: color_data = Z;
		19'b1011100110100110010: color_data = Z;
		19'b1011100110100110011: color_data = Z;
		19'b1011100110100110100: color_data = Z;
		19'b1011100110100110101: color_data = Z;
		19'b1011100110100110110: color_data = Z;
		19'b1011100110100110111: color_data = Z;
		19'b1011100110100111000: color_data = Z;
		19'b1011100110100111001: color_data = Z;
		19'b1011100110100111010: color_data = Z;
		19'b1011100110101011101: color_data = Z;
		19'b1011100110101011110: color_data = Z;
		19'b1011100110101011111: color_data = Z;
		19'b1011100110101100000: color_data = Z;
		19'b1011100110101100001: color_data = Z;
		19'b1011100110101100010: color_data = Z;
		19'b1011100110101100011: color_data = Z;
		19'b1011100110101100100: color_data = Z;
		19'b1011100110101100101: color_data = Z;
		19'b1011100110101100110: color_data = Z;
		19'b1011100110101100111: color_data = Z;
		19'b1011100110101101000: color_data = Z;
		19'b1011100110101101001: color_data = Z;
		19'b1011100110101101010: color_data = Z;
		19'b1011100110101101011: color_data = Z;
		19'b1011100110101101100: color_data = Z;
		19'b1011100110101101101: color_data = Z;
		19'b1011100110101101110: color_data = Z;
		19'b1011100110101101111: color_data = Z;
		19'b1011100110101110000: color_data = Z;
		19'b1011100110101110001: color_data = Z;
		19'b1011100110101110010: color_data = Z;
		19'b1011100110101110011: color_data = Z;
		19'b1011100110101110100: color_data = Z;
		19'b1011100110101110101: color_data = Z;
		19'b1011100110101110110: color_data = Z;
		19'b1011100110101110111: color_data = Z;
		19'b1011100110101111000: color_data = Z;
		19'b1011100110101111001: color_data = Z;
		19'b1011100110101111010: color_data = Z;
		19'b1011100110101111011: color_data = Z;
		19'b1011100110101111100: color_data = Z;
		19'b1011100110101111101: color_data = Z;
		19'b1011100110101111110: color_data = Z;
		19'b1011100110101111111: color_data = Z;
		19'b1011100110110000000: color_data = Z;
		19'b1011100110110000001: color_data = Z;
		19'b1011100110110000010: color_data = Z;
		19'b1011100110110000011: color_data = Z;
		19'b1011100110110000100: color_data = Z;
		19'b1011100110110000101: color_data = Z;
		19'b1011100110110000110: color_data = Z;
		19'b1011100110110000111: color_data = Z;
		19'b1011100110110001000: color_data = Z;
		19'b1011100110110001001: color_data = Z;
		19'b1011100110110001010: color_data = Z;
		19'b1011100110110001011: color_data = Z;
		19'b1011100110110001100: color_data = Z;
		19'b1011100110110001101: color_data = Z;
		19'b1011100110110001110: color_data = Z;
		19'b1011100110110001111: color_data = Z;
		19'b1011100110110010000: color_data = Z;
		19'b1011100110110010001: color_data = Z;
		19'b1011100110110010010: color_data = Z;
		19'b1011101000011111001: color_data = Z;
		19'b1011101000011111010: color_data = Z;
		19'b1011101000011111011: color_data = Z;
		19'b1011101000011111100: color_data = Z;
		19'b1011101000011111101: color_data = Z;
		19'b1011101000011111110: color_data = Z;
		19'b1011101000011111111: color_data = Z;
		19'b1011101000100000000: color_data = Z;
		19'b1011101000100000001: color_data = Z;
		19'b1011101000100000010: color_data = Z;
		19'b1011101000100000011: color_data = Z;
		19'b1011101000100000100: color_data = Z;
		19'b1011101000100000101: color_data = Z;
		19'b1011101000100000110: color_data = Z;
		19'b1011101000100000111: color_data = Z;
		19'b1011101000100001000: color_data = Z;
		19'b1011101000100001001: color_data = Z;
		19'b1011101000100001010: color_data = Z;
		19'b1011101000100001011: color_data = Z;
		19'b1011101000100001100: color_data = Z;
		19'b1011101000100001101: color_data = Z;
		19'b1011101000100001110: color_data = Z;
		19'b1011101000100001111: color_data = Z;
		19'b1011101000100010000: color_data = Z;
		19'b1011101000100010001: color_data = Z;
		19'b1011101000100010010: color_data = Z;
		19'b1011101000100010011: color_data = Z;
		19'b1011101000100010100: color_data = Z;
		19'b1011101000100010101: color_data = Z;
		19'b1011101000100010110: color_data = Z;
		19'b1011101000100010111: color_data = Z;
		19'b1011101000100011000: color_data = Z;
		19'b1011101000100011001: color_data = Z;
		19'b1011101000100011010: color_data = Z;
		19'b1011101000100011011: color_data = Z;
		19'b1011101000100011100: color_data = Z;
		19'b1011101000100011101: color_data = Z;
		19'b1011101000100011110: color_data = Z;
		19'b1011101000100011111: color_data = Z;
		19'b1011101000100100000: color_data = Z;
		19'b1011101000100100001: color_data = Z;
		19'b1011101000100100010: color_data = Z;
		19'b1011101000100100011: color_data = Z;
		19'b1011101000100100100: color_data = Z;
		19'b1011101000100100101: color_data = Z;
		19'b1011101000100100110: color_data = Z;
		19'b1011101000100100111: color_data = Z;
		19'b1011101000100101000: color_data = Z;
		19'b1011101000100101001: color_data = Z;
		19'b1011101000100101010: color_data = Z;
		19'b1011101000100101011: color_data = Z;
		19'b1011101000100101100: color_data = Z;
		19'b1011101000100101101: color_data = Z;
		19'b1011101000100101110: color_data = Z;
		19'b1011101000100101111: color_data = Z;
		19'b1011101000100110000: color_data = Z;
		19'b1011101000100110001: color_data = Z;
		19'b1011101000100110010: color_data = Z;
		19'b1011101000100110011: color_data = Z;
		19'b1011101000100110100: color_data = Z;
		19'b1011101000100110101: color_data = Z;
		19'b1011101000100110110: color_data = Z;
		19'b1011101000100110111: color_data = Z;
		19'b1011101000100111000: color_data = Z;
		19'b1011101000100111001: color_data = Z;
		19'b1011101000100111010: color_data = Z;
		19'b1011101000100111011: color_data = Z;
		19'b1011101000100111100: color_data = Z;
		19'b1011101000101000000: color_data = Z;
		19'b1011101000101010010: color_data = Z;
		19'b1011101000101010011: color_data = Z;
		19'b1011101000101010100: color_data = Z;
		19'b1011101000101010101: color_data = Z;
		19'b1011101000101010110: color_data = Z;
		19'b1011101000101010111: color_data = Z;
		19'b1011101000101011000: color_data = Z;
		19'b1011101000101011001: color_data = Z;
		19'b1011101000101011010: color_data = Z;
		19'b1011101000101011011: color_data = Z;
		19'b1011101000101011100: color_data = Z;
		19'b1011101000101011101: color_data = Z;
		19'b1011101000101011110: color_data = Z;
		19'b1011101000101011111: color_data = Z;
		19'b1011101000101100000: color_data = Z;
		19'b1011101000101100001: color_data = Z;
		19'b1011101000101100010: color_data = Z;
		19'b1011101000101100011: color_data = Z;
		19'b1011101000101100100: color_data = Z;
		19'b1011101000101100101: color_data = Z;
		19'b1011101000101100110: color_data = Z;
		19'b1011101000101100111: color_data = Z;
		19'b1011101000101101000: color_data = Z;
		19'b1011101000101101001: color_data = Z;
		19'b1011101000101101010: color_data = Z;
		19'b1011101000101101011: color_data = Z;
		19'b1011101000101101100: color_data = Z;
		19'b1011101000101101101: color_data = Z;
		19'b1011101000101101110: color_data = Z;
		19'b1011101000101101111: color_data = Z;
		19'b1011101000101110000: color_data = Z;
		19'b1011101000101110001: color_data = Z;
		19'b1011101000101110010: color_data = Z;
		19'b1011101000101110011: color_data = Z;
		19'b1011101000101110100: color_data = Z;
		19'b1011101000101110101: color_data = Z;
		19'b1011101000101110110: color_data = Z;
		19'b1011101000101110111: color_data = Z;
		19'b1011101000101111000: color_data = Z;
		19'b1011101000101111001: color_data = Z;
		19'b1011101000101111010: color_data = Z;
		19'b1011101000101111011: color_data = Z;
		19'b1011101000101111100: color_data = Z;
		19'b1011101000101111101: color_data = Z;
		19'b1011101000101111110: color_data = Z;
		19'b1011101000101111111: color_data = Z;
		19'b1011101000110000000: color_data = Z;
		19'b1011101000110000001: color_data = Z;
		19'b1011101000110000010: color_data = Z;
		19'b1011101000110000011: color_data = Z;
		19'b1011101000110000100: color_data = Z;
		19'b1011101000110000101: color_data = Z;
		19'b1011101000110000110: color_data = Z;
		19'b1011101000110000111: color_data = Z;
		19'b1011101000110001000: color_data = Z;
		19'b1011101000110001001: color_data = Z;
		19'b1011101000110001010: color_data = Z;
		19'b1011101000110001011: color_data = Z;
		19'b1011101000110001100: color_data = Z;
		19'b1011101000110001101: color_data = Z;
		19'b1011101000110001110: color_data = Z;
		19'b1011101000110001111: color_data = Z;
		19'b1011101000110010000: color_data = Z;
		19'b1011101000110010001: color_data = Z;
		19'b1011101010011111011: color_data = Z;
		19'b1011101010011111100: color_data = Z;
		19'b1011101010011111101: color_data = Z;
		19'b1011101010011111110: color_data = Z;
		19'b1011101010011111111: color_data = Z;
		19'b1011101010100000000: color_data = Z;
		19'b1011101010100000001: color_data = Z;
		19'b1011101010100000010: color_data = Z;
		19'b1011101010100000011: color_data = Z;
		19'b1011101010100000100: color_data = Z;
		19'b1011101010100000101: color_data = Z;
		19'b1011101010100000110: color_data = Z;
		19'b1011101010100000111: color_data = Z;
		19'b1011101010100001000: color_data = Z;
		19'b1011101010100001001: color_data = Z;
		19'b1011101010100001010: color_data = Z;
		19'b1011101010100001011: color_data = Z;
		19'b1011101010100001100: color_data = Z;
		19'b1011101010100001101: color_data = Z;
		19'b1011101010100001110: color_data = Z;
		19'b1011101010100001111: color_data = Z;
		19'b1011101010100010000: color_data = Z;
		19'b1011101010100010001: color_data = Z;
		19'b1011101010100010010: color_data = Z;
		19'b1011101010100010011: color_data = Z;
		19'b1011101010100010100: color_data = Z;
		19'b1011101010100010101: color_data = Z;
		19'b1011101010100010110: color_data = Z;
		19'b1011101010100010111: color_data = Z;
		19'b1011101010100011000: color_data = Z;
		19'b1011101010100011001: color_data = Z;
		19'b1011101010100011010: color_data = Z;
		19'b1011101010100011011: color_data = Z;
		19'b1011101010100011100: color_data = Z;
		19'b1011101010100011101: color_data = Z;
		19'b1011101010100011110: color_data = Z;
		19'b1011101010100011111: color_data = Z;
		19'b1011101010100100000: color_data = Z;
		19'b1011101010100100001: color_data = Z;
		19'b1011101010100100010: color_data = Z;
		19'b1011101010100100011: color_data = Z;
		19'b1011101010100100100: color_data = Z;
		19'b1011101010100100101: color_data = Z;
		19'b1011101010100100110: color_data = Z;
		19'b1011101010100100111: color_data = Z;
		19'b1011101010100101000: color_data = Z;
		19'b1011101010100101001: color_data = Z;
		19'b1011101010100101010: color_data = Z;
		19'b1011101010100101011: color_data = Z;
		19'b1011101010100101100: color_data = Z;
		19'b1011101010100101101: color_data = Z;
		19'b1011101010100101110: color_data = Z;
		19'b1011101010100101111: color_data = Z;
		19'b1011101010100110000: color_data = Z;
		19'b1011101010100110001: color_data = Z;
		19'b1011101010100110010: color_data = Z;
		19'b1011101010100110011: color_data = Z;
		19'b1011101010100110100: color_data = Z;
		19'b1011101010100110101: color_data = Z;
		19'b1011101010100110110: color_data = Z;
		19'b1011101010100110111: color_data = Z;
		19'b1011101010100111000: color_data = Z;
		19'b1011101010100111001: color_data = Z;
		19'b1011101010100111010: color_data = Z;
		19'b1011101010100111011: color_data = Z;
		19'b1011101010100111100: color_data = Z;
		19'b1011101010100111101: color_data = Z;
		19'b1011101010100111110: color_data = Z;
		19'b1011101010100111111: color_data = Z;
		19'b1011101010101000000: color_data = Z;
		19'b1011101010101000001: color_data = Z;
		19'b1011101010101000010: color_data = Z;
		19'b1011101010101000011: color_data = Z;
		19'b1011101010101000100: color_data = Z;
		19'b1011101010101000101: color_data = Z;
		19'b1011101010101000110: color_data = Z;
		19'b1011101010101000111: color_data = Z;
		19'b1011101010101001000: color_data = Z;
		19'b1011101010101001001: color_data = Z;
		19'b1011101010101001010: color_data = Z;
		19'b1011101010101001011: color_data = Z;
		19'b1011101010101001100: color_data = Z;
		19'b1011101010101001101: color_data = Z;
		19'b1011101010101001110: color_data = Z;
		19'b1011101010101001111: color_data = Z;
		19'b1011101010101010000: color_data = Z;
		19'b1011101010101010001: color_data = Z;
		19'b1011101010101010010: color_data = Z;
		19'b1011101010101010011: color_data = Z;
		19'b1011101010101010100: color_data = Z;
		19'b1011101010101010101: color_data = Z;
		19'b1011101010101010110: color_data = Z;
		19'b1011101010101010111: color_data = Z;
		19'b1011101010101011000: color_data = Z;
		19'b1011101010101011001: color_data = Z;
		19'b1011101010101011010: color_data = Z;
		19'b1011101010101011011: color_data = Z;
		19'b1011101010101011100: color_data = Z;
		19'b1011101010101011101: color_data = Z;
		19'b1011101010101011110: color_data = Z;
		19'b1011101010101011111: color_data = Z;
		19'b1011101010101100000: color_data = Z;
		19'b1011101010101100001: color_data = Z;
		19'b1011101010101100010: color_data = Z;
		19'b1011101010101100011: color_data = Z;
		19'b1011101010101100100: color_data = Z;
		19'b1011101010101100101: color_data = Z;
		19'b1011101010101100110: color_data = Z;
		19'b1011101010101100111: color_data = Z;
		19'b1011101010101101000: color_data = Z;
		19'b1011101010101101001: color_data = Z;
		19'b1011101010101101010: color_data = Z;
		19'b1011101010101101011: color_data = Z;
		19'b1011101010101101100: color_data = Z;
		19'b1011101010101101101: color_data = Z;
		19'b1011101010101101110: color_data = Z;
		19'b1011101010101101111: color_data = Z;
		19'b1011101010101110000: color_data = Z;
		19'b1011101010101110001: color_data = Z;
		19'b1011101010101110010: color_data = Z;
		19'b1011101010101110011: color_data = Z;
		19'b1011101010101110100: color_data = Z;
		19'b1011101010101110101: color_data = Z;
		19'b1011101010101110110: color_data = Z;
		19'b1011101010101110111: color_data = Z;
		19'b1011101010101111000: color_data = Z;
		19'b1011101010101111001: color_data = Z;
		19'b1011101010101111010: color_data = Z;
		19'b1011101010101111011: color_data = Z;
		19'b1011101010101111100: color_data = Z;
		19'b1011101010101111101: color_data = Z;
		19'b1011101010101111110: color_data = Z;
		19'b1011101010101111111: color_data = Z;
		19'b1011101010110000000: color_data = Z;
		19'b1011101010110000001: color_data = Z;
		19'b1011101010110000010: color_data = Z;
		19'b1011101010110000011: color_data = Z;
		19'b1011101010110000100: color_data = Z;
		19'b1011101010110000101: color_data = Z;
		19'b1011101010110000110: color_data = Z;
		19'b1011101010110000111: color_data = Z;
		19'b1011101010110001000: color_data = Z;
		19'b1011101010110001001: color_data = Z;
		19'b1011101010110001010: color_data = Z;
		19'b1011101010110001011: color_data = Z;
		19'b1011101010110001100: color_data = Z;
		19'b1011101010110001101: color_data = Z;
		19'b1011101010110001110: color_data = Z;
		19'b1011101010110001111: color_data = Z;
		19'b1011101010110010000: color_data = Z;
		19'b1011101100011111101: color_data = Z;
		19'b1011101100011111110: color_data = Z;
		19'b1011101100011111111: color_data = Z;
		19'b1011101100100000000: color_data = Z;
		19'b1011101100100000001: color_data = Z;
		19'b1011101100100000010: color_data = Z;
		19'b1011101100100000011: color_data = Z;
		19'b1011101100100000100: color_data = Z;
		19'b1011101100100000101: color_data = Z;
		19'b1011101100100000110: color_data = Z;
		19'b1011101100100000111: color_data = Z;
		19'b1011101100100001000: color_data = Z;
		19'b1011101100100001001: color_data = Z;
		19'b1011101100100001010: color_data = Z;
		19'b1011101100100001011: color_data = Z;
		19'b1011101100100001100: color_data = Z;
		19'b1011101100100001101: color_data = Z;
		19'b1011101100100001110: color_data = Z;
		19'b1011101100100001111: color_data = Z;
		19'b1011101100100010000: color_data = Z;
		19'b1011101100100010001: color_data = Z;
		19'b1011101100100010010: color_data = Z;
		19'b1011101100100010011: color_data = Z;
		19'b1011101100100010100: color_data = Z;
		19'b1011101100100010101: color_data = Z;
		19'b1011101100100010110: color_data = Z;
		19'b1011101100100010111: color_data = Z;
		19'b1011101100100011000: color_data = Z;
		19'b1011101100100011001: color_data = Z;
		19'b1011101100100011010: color_data = Z;
		19'b1011101100100011011: color_data = Z;
		19'b1011101100100011100: color_data = Z;
		19'b1011101100100011101: color_data = Z;
		19'b1011101100100011110: color_data = Z;
		19'b1011101100100011111: color_data = Z;
		19'b1011101100100100000: color_data = Z;
		19'b1011101100100100001: color_data = Z;
		19'b1011101100100100010: color_data = Z;
		19'b1011101100100100011: color_data = Z;
		19'b1011101100100100100: color_data = Z;
		19'b1011101100100100101: color_data = Z;
		19'b1011101100100100110: color_data = Z;
		19'b1011101100100100111: color_data = Z;
		19'b1011101100100101000: color_data = Z;
		19'b1011101100100101001: color_data = Z;
		19'b1011101100100101010: color_data = Z;
		19'b1011101100100101011: color_data = Z;
		19'b1011101100100101100: color_data = Z;
		19'b1011101100100101101: color_data = Z;
		19'b1011101100100101110: color_data = Z;
		19'b1011101100100101111: color_data = Z;
		19'b1011101100100110000: color_data = Z;
		19'b1011101100100110001: color_data = Z;
		19'b1011101100100110010: color_data = Z;
		19'b1011101100100110011: color_data = Z;
		19'b1011101100100110100: color_data = Z;
		19'b1011101100100110101: color_data = Z;
		19'b1011101100100110110: color_data = Z;
		19'b1011101100100110111: color_data = Z;
		19'b1011101100100111000: color_data = Z;
		19'b1011101100100111001: color_data = Z;
		19'b1011101100100111010: color_data = Z;
		19'b1011101100100111011: color_data = Z;
		19'b1011101100100111100: color_data = Z;
		19'b1011101100100111101: color_data = Z;
		19'b1011101100100111110: color_data = Z;
		19'b1011101100100111111: color_data = Z;
		19'b1011101100101000000: color_data = Z;
		19'b1011101100101000001: color_data = Z;
		19'b1011101100101000010: color_data = Z;
		19'b1011101100101000011: color_data = Z;
		19'b1011101100101000100: color_data = Z;
		19'b1011101100101000101: color_data = Z;
		19'b1011101100101000110: color_data = Z;
		19'b1011101100101000111: color_data = Z;
		19'b1011101100101001000: color_data = Z;
		19'b1011101100101001001: color_data = Z;
		19'b1011101100101001010: color_data = Z;
		19'b1011101100101001011: color_data = Z;
		19'b1011101100101001100: color_data = Z;
		19'b1011101100101001101: color_data = Z;
		19'b1011101100101001110: color_data = Z;
		19'b1011101100101001111: color_data = Z;
		19'b1011101100101010000: color_data = Z;
		19'b1011101100101010001: color_data = Z;
		19'b1011101100101010010: color_data = Z;
		19'b1011101100101010011: color_data = Z;
		19'b1011101100101010100: color_data = Z;
		19'b1011101100101010101: color_data = Z;
		19'b1011101100101010110: color_data = Z;
		19'b1011101100101010111: color_data = Z;
		19'b1011101100101011000: color_data = Z;
		19'b1011101100101011001: color_data = Z;
		19'b1011101100101011010: color_data = Z;
		19'b1011101100101011011: color_data = Z;
		19'b1011101100101011100: color_data = Z;
		19'b1011101100101011101: color_data = Z;
		19'b1011101100101011110: color_data = Z;
		19'b1011101100101011111: color_data = Z;
		19'b1011101100101100000: color_data = Z;
		19'b1011101100101100001: color_data = Z;
		19'b1011101100101100010: color_data = Z;
		19'b1011101100101100011: color_data = Z;
		19'b1011101100101100100: color_data = Z;
		19'b1011101100101100101: color_data = Z;
		19'b1011101100101100110: color_data = Z;
		19'b1011101100101100111: color_data = Z;
		19'b1011101100101101000: color_data = Z;
		19'b1011101100101101001: color_data = Z;
		19'b1011101100101101010: color_data = Z;
		19'b1011101100101101011: color_data = Z;
		19'b1011101100101101100: color_data = Z;
		19'b1011101100101101101: color_data = Z;
		19'b1011101100101101110: color_data = Z;
		19'b1011101100101101111: color_data = Z;
		19'b1011101100101110000: color_data = Z;
		19'b1011101100101110001: color_data = Z;
		19'b1011101100101110010: color_data = Z;
		19'b1011101100101110011: color_data = Z;
		19'b1011101100101110100: color_data = Z;
		19'b1011101100101110101: color_data = Z;
		19'b1011101100101110110: color_data = Z;
		19'b1011101100101110111: color_data = Z;
		19'b1011101100101111000: color_data = Z;
		19'b1011101100101111001: color_data = Z;
		19'b1011101100101111010: color_data = Z;
		19'b1011101100101111011: color_data = Z;
		19'b1011101100101111100: color_data = Z;
		19'b1011101100101111101: color_data = Z;
		19'b1011101100101111110: color_data = Z;
		19'b1011101100101111111: color_data = Z;
		19'b1011101100110000000: color_data = Z;
		19'b1011101100110000001: color_data = Z;
		19'b1011101100110000010: color_data = Z;
		19'b1011101100110000011: color_data = Z;
		19'b1011101100110000100: color_data = Z;
		19'b1011101100110000101: color_data = Z;
		19'b1011101100110000110: color_data = Z;
		19'b1011101100110000111: color_data = Z;
		19'b1011101100110001000: color_data = Z;
		19'b1011101100110001001: color_data = Z;
		19'b1011101100110001010: color_data = Z;
		19'b1011101100110001011: color_data = Z;
		19'b1011101100110001100: color_data = Z;
		19'b1011101100110001101: color_data = Z;
		19'b1011101110100000000: color_data = Z;
		19'b1011101110100000001: color_data = Z;
		19'b1011101110100000010: color_data = Z;
		19'b1011101110100000011: color_data = Z;
		19'b1011101110100000100: color_data = Z;
		19'b1011101110100000101: color_data = Z;
		19'b1011101110100000110: color_data = Z;
		19'b1011101110100000111: color_data = Z;
		19'b1011101110100001000: color_data = Z;
		19'b1011101110100001001: color_data = Z;
		19'b1011101110100001010: color_data = Z;
		19'b1011101110100001011: color_data = Z;
		19'b1011101110100001100: color_data = Z;
		19'b1011101110100001101: color_data = Z;
		19'b1011101110100001110: color_data = Z;
		19'b1011101110100001111: color_data = Z;
		19'b1011101110100010000: color_data = Z;
		19'b1011101110100010001: color_data = Z;
		19'b1011101110100010010: color_data = Z;
		19'b1011101110100010011: color_data = Z;
		19'b1011101110100010100: color_data = Z;
		19'b1011101110100010101: color_data = Z;
		19'b1011101110100010110: color_data = Z;
		19'b1011101110100010111: color_data = Z;
		19'b1011101110100011000: color_data = Z;
		19'b1011101110100011001: color_data = Z;
		19'b1011101110100011010: color_data = Z;
		19'b1011101110100011011: color_data = Z;
		19'b1011101110100011100: color_data = Z;
		19'b1011101110100011101: color_data = Z;
		19'b1011101110100011110: color_data = Z;
		19'b1011101110100011111: color_data = Z;
		19'b1011101110100100000: color_data = Z;
		19'b1011101110100100001: color_data = Z;
		19'b1011101110100100010: color_data = Z;
		19'b1011101110100100011: color_data = Z;
		19'b1011101110100100100: color_data = Z;
		19'b1011101110100100101: color_data = Z;
		19'b1011101110100100110: color_data = Z;
		19'b1011101110100100111: color_data = Z;
		19'b1011101110100101000: color_data = Z;
		19'b1011101110100101001: color_data = Z;
		19'b1011101110100101010: color_data = Z;
		19'b1011101110100101011: color_data = Z;
		19'b1011101110100101100: color_data = Z;
		19'b1011101110100101101: color_data = Z;
		19'b1011101110100101110: color_data = Z;
		19'b1011101110100101111: color_data = Z;
		19'b1011101110100110000: color_data = Z;
		19'b1011101110100110001: color_data = Z;
		19'b1011101110100110010: color_data = Z;
		19'b1011101110100110011: color_data = Z;
		19'b1011101110100110100: color_data = Z;
		19'b1011101110100110101: color_data = Z;
		19'b1011101110100110110: color_data = Z;
		19'b1011101110100110111: color_data = Z;
		19'b1011101110100111000: color_data = Z;
		19'b1011101110100111001: color_data = Z;
		19'b1011101110100111010: color_data = Z;
		19'b1011101110100111011: color_data = Z;
		19'b1011101110100111100: color_data = Z;
		19'b1011101110100111101: color_data = Z;
		19'b1011101110100111110: color_data = Z;
		19'b1011101110100111111: color_data = Z;
		19'b1011101110101000000: color_data = Z;
		19'b1011101110101000001: color_data = Z;
		19'b1011101110101000010: color_data = Z;
		19'b1011101110101000011: color_data = Z;
		19'b1011101110101000100: color_data = Z;
		19'b1011101110101000101: color_data = Z;
		19'b1011101110101000110: color_data = Z;
		19'b1011101110101000111: color_data = Z;
		19'b1011101110101001000: color_data = Z;
		19'b1011101110101001001: color_data = Z;
		19'b1011101110101001010: color_data = Z;
		19'b1011101110101001011: color_data = Z;
		19'b1011101110101001100: color_data = Z;
		19'b1011101110101001101: color_data = Z;
		19'b1011101110101001110: color_data = Z;
		19'b1011101110101001111: color_data = Z;
		19'b1011101110101010000: color_data = Z;
		19'b1011101110101010001: color_data = Z;
		19'b1011101110101010010: color_data = Z;
		19'b1011101110101010011: color_data = Z;
		19'b1011101110101010100: color_data = Z;
		19'b1011101110101010101: color_data = Z;
		19'b1011101110101010110: color_data = Z;
		19'b1011101110101010111: color_data = Z;
		19'b1011101110101011000: color_data = Z;
		19'b1011101110101011001: color_data = Z;
		19'b1011101110101011010: color_data = Z;
		19'b1011101110101011011: color_data = Z;
		19'b1011101110101011100: color_data = Z;
		19'b1011101110101011101: color_data = Z;
		19'b1011101110101011110: color_data = Z;
		19'b1011101110101011111: color_data = Z;
		19'b1011101110101100000: color_data = Z;
		19'b1011101110101100001: color_data = Z;
		19'b1011101110101100010: color_data = Z;
		19'b1011101110101100011: color_data = Z;
		19'b1011101110101100100: color_data = Z;
		19'b1011101110101100101: color_data = Z;
		19'b1011101110101100110: color_data = Z;
		19'b1011101110101100111: color_data = Z;
		19'b1011101110101101000: color_data = Z;
		19'b1011101110101101001: color_data = Z;
		19'b1011101110101101010: color_data = Z;
		19'b1011101110101101011: color_data = Z;
		19'b1011101110101101100: color_data = Z;
		19'b1011101110101101101: color_data = Z;
		19'b1011101110101101110: color_data = Z;
		19'b1011101110101101111: color_data = Z;
		19'b1011101110101110000: color_data = Z;
		19'b1011101110101110001: color_data = Z;
		19'b1011101110101110010: color_data = Z;
		19'b1011101110101110011: color_data = Z;
		19'b1011101110101110100: color_data = Z;
		19'b1011101110101110101: color_data = Z;
		19'b1011101110101110110: color_data = Z;
		19'b1011101110101110111: color_data = Z;
		19'b1011101110101111000: color_data = Z;
		19'b1011101110101111001: color_data = Z;
		19'b1011101110101111010: color_data = Z;
		19'b1011101110101111011: color_data = Z;
		19'b1011101110101111100: color_data = Z;
		19'b1011101110101111101: color_data = Z;
		19'b1011101110101111110: color_data = Z;
		19'b1011101110101111111: color_data = Z;
		19'b1011101110110000000: color_data = Z;
		19'b1011101110110000001: color_data = Z;
		19'b1011101110110000010: color_data = Z;
		19'b1011101110110000011: color_data = Z;
		19'b1011101110110000100: color_data = Z;
		19'b1011101110110000101: color_data = Z;
		19'b1011101110110000110: color_data = Z;
		19'b1011101110110000111: color_data = Z;
		19'b1011101110110001000: color_data = Z;
		19'b1011101110110001001: color_data = Z;
		19'b1011101110110001010: color_data = Z;
		19'b1011101110110001011: color_data = Z;
		19'b1011110000100000011: color_data = Z;
		19'b1011110000100000100: color_data = Z;
		19'b1011110000100000101: color_data = Z;
		19'b1011110000100000110: color_data = Z;
		19'b1011110000100000111: color_data = Z;
		19'b1011110000100001000: color_data = Z;
		19'b1011110000100001001: color_data = Z;
		19'b1011110000100001010: color_data = Z;
		19'b1011110000100001011: color_data = Z;
		19'b1011110000100001100: color_data = Z;
		19'b1011110000100001101: color_data = Z;
		19'b1011110000100001110: color_data = Z;
		19'b1011110000100001111: color_data = Z;
		19'b1011110000100010000: color_data = Z;
		19'b1011110000100010001: color_data = Z;
		19'b1011110000100010010: color_data = Z;
		19'b1011110000100010011: color_data = Z;
		19'b1011110000100010100: color_data = Z;
		19'b1011110000100010101: color_data = Z;
		19'b1011110000100010110: color_data = Z;
		19'b1011110000100010111: color_data = Z;
		19'b1011110000100011000: color_data = Z;
		19'b1011110000100011001: color_data = Z;
		19'b1011110000100011010: color_data = Z;
		19'b1011110000100011011: color_data = Z;
		19'b1011110000100011100: color_data = Z;
		19'b1011110000100011101: color_data = Z;
		19'b1011110000100011110: color_data = Z;
		19'b1011110000100011111: color_data = Z;
		19'b1011110000100100000: color_data = Z;
		19'b1011110000100100001: color_data = Z;
		19'b1011110000100100010: color_data = Z;
		19'b1011110000100100011: color_data = Z;
		19'b1011110000100100100: color_data = Z;
		19'b1011110000100100101: color_data = Z;
		19'b1011110000100100110: color_data = Z;
		19'b1011110000100100111: color_data = Z;
		19'b1011110000100101000: color_data = Z;
		19'b1011110000100101001: color_data = Z;
		19'b1011110000100101010: color_data = Z;
		19'b1011110000100101011: color_data = Z;
		19'b1011110000100101100: color_data = Z;
		19'b1011110000100101101: color_data = Z;
		19'b1011110000100101110: color_data = Z;
		19'b1011110000100101111: color_data = Z;
		19'b1011110000100110000: color_data = Z;
		19'b1011110000100110001: color_data = Z;
		19'b1011110000100110010: color_data = Z;
		19'b1011110000100110011: color_data = Z;
		19'b1011110000100110100: color_data = Z;
		19'b1011110000100110101: color_data = Z;
		19'b1011110000100110110: color_data = Z;
		19'b1011110000100110111: color_data = Z;
		19'b1011110000100111000: color_data = Z;
		19'b1011110000100111001: color_data = Z;
		19'b1011110000100111010: color_data = Z;
		19'b1011110000100111011: color_data = Z;
		19'b1011110000100111100: color_data = Z;
		19'b1011110000100111101: color_data = Z;
		19'b1011110000100111110: color_data = Z;
		19'b1011110000100111111: color_data = Z;
		19'b1011110000101000000: color_data = Z;
		19'b1011110000101000001: color_data = Z;
		19'b1011110000101000010: color_data = Z;
		19'b1011110000101000011: color_data = Z;
		19'b1011110000101000100: color_data = Z;
		19'b1011110000101000101: color_data = Z;
		19'b1011110000101000110: color_data = Z;
		19'b1011110000101000111: color_data = Z;
		19'b1011110000101001000: color_data = Z;
		19'b1011110000101001001: color_data = Z;
		19'b1011110000101001010: color_data = Z;
		19'b1011110000101001011: color_data = Z;
		19'b1011110000101001100: color_data = Z;
		19'b1011110000101001101: color_data = Z;
		19'b1011110000101001110: color_data = Z;
		19'b1011110000101001111: color_data = Z;
		19'b1011110000101010000: color_data = Z;
		19'b1011110000101010001: color_data = Z;
		19'b1011110000101010010: color_data = Z;
		19'b1011110000101010011: color_data = Z;
		19'b1011110000101010100: color_data = Z;
		19'b1011110000101010101: color_data = Z;
		19'b1011110000101010110: color_data = Z;
		19'b1011110000101010111: color_data = Z;
		19'b1011110000101011000: color_data = Z;
		19'b1011110000101011001: color_data = Z;
		19'b1011110000101011010: color_data = Z;
		19'b1011110000101011011: color_data = Z;
		19'b1011110000101011100: color_data = Z;
		19'b1011110000101011101: color_data = Z;
		19'b1011110000101011110: color_data = Z;
		19'b1011110000101011111: color_data = Z;
		19'b1011110000101100000: color_data = Z;
		19'b1011110000101100001: color_data = Z;
		19'b1011110000101100010: color_data = Z;
		19'b1011110000101100011: color_data = Z;
		19'b1011110000101100100: color_data = Z;
		19'b1011110000101100101: color_data = Z;
		19'b1011110000101100110: color_data = Z;
		19'b1011110000101100111: color_data = Z;
		19'b1011110000101101000: color_data = Z;
		19'b1011110000101101001: color_data = Z;
		19'b1011110000101101010: color_data = Z;
		19'b1011110000101101011: color_data = Z;
		19'b1011110000101101100: color_data = Z;
		19'b1011110000101101101: color_data = Z;
		19'b1011110000101101110: color_data = Z;
		19'b1011110000101101111: color_data = Z;
		19'b1011110000101110000: color_data = Z;
		19'b1011110000101110001: color_data = Z;
		19'b1011110000101110010: color_data = Z;
		19'b1011110000101110011: color_data = Z;
		19'b1011110000101110100: color_data = Z;
		19'b1011110000101110101: color_data = Z;
		19'b1011110000101110110: color_data = Z;
		19'b1011110000101110111: color_data = Z;
		19'b1011110000101111000: color_data = Z;
		19'b1011110000101111001: color_data = Z;
		19'b1011110000101111010: color_data = Z;
		19'b1011110000101111011: color_data = Z;
		19'b1011110000101111100: color_data = Z;
		19'b1011110000101111101: color_data = Z;
		19'b1011110000101111110: color_data = Z;
		19'b1011110000101111111: color_data = Z;
		19'b1011110000110000000: color_data = Z;
		19'b1011110000110000001: color_data = Z;
		19'b1011110000110000010: color_data = Z;
		19'b1011110000110000011: color_data = Z;
		19'b1011110000110000100: color_data = Z;
		19'b1011110000110000101: color_data = Z;
		19'b1011110000110000110: color_data = Z;
		19'b1011110000110000111: color_data = Z;
		19'b1011110000110001000: color_data = Z;
		19'b1011110000110001001: color_data = Z;
		19'b1011110010100000101: color_data = Z;
		19'b1011110010100000110: color_data = Z;
		19'b1011110010100000111: color_data = Z;
		19'b1011110010100001000: color_data = Z;
		19'b1011110010100001001: color_data = Z;
		19'b1011110010100001010: color_data = Z;
		19'b1011110010100001011: color_data = Z;
		19'b1011110010100001100: color_data = Z;
		19'b1011110010100001101: color_data = Z;
		19'b1011110010100001110: color_data = Z;
		19'b1011110010100001111: color_data = Z;
		19'b1011110010100010000: color_data = Z;
		19'b1011110010100010001: color_data = Z;
		19'b1011110010100010010: color_data = Z;
		19'b1011110010100010011: color_data = Z;
		19'b1011110010100010100: color_data = Z;
		19'b1011110010100010101: color_data = Z;
		19'b1011110010100010110: color_data = Z;
		19'b1011110010100010111: color_data = Z;
		19'b1011110010100011000: color_data = Z;
		19'b1011110010100011001: color_data = Z;
		19'b1011110010100011010: color_data = Z;
		19'b1011110010100011011: color_data = Z;
		19'b1011110010100011100: color_data = Z;
		19'b1011110010100011101: color_data = Z;
		19'b1011110010100011110: color_data = Z;
		19'b1011110010100011111: color_data = Z;
		19'b1011110010100100000: color_data = Z;
		19'b1011110010100100001: color_data = Z;
		19'b1011110010100100010: color_data = Z;
		19'b1011110010100100011: color_data = Z;
		19'b1011110010100100100: color_data = Z;
		19'b1011110010100100101: color_data = Z;
		19'b1011110010100100110: color_data = Z;
		19'b1011110010100100111: color_data = Z;
		19'b1011110010100101000: color_data = Z;
		19'b1011110010100101001: color_data = Z;
		19'b1011110010100101010: color_data = Z;
		19'b1011110010100101011: color_data = Z;
		19'b1011110010100101100: color_data = Z;
		19'b1011110010100101101: color_data = Z;
		19'b1011110010100101110: color_data = Z;
		19'b1011110010100101111: color_data = Z;
		19'b1011110010100110000: color_data = Z;
		19'b1011110010100110001: color_data = Z;
		19'b1011110010100110010: color_data = Z;
		19'b1011110010100110011: color_data = Z;
		19'b1011110010100110100: color_data = Z;
		19'b1011110010100110101: color_data = Z;
		19'b1011110010100110110: color_data = Z;
		19'b1011110010100110111: color_data = Z;
		19'b1011110010100111000: color_data = Z;
		19'b1011110010100111001: color_data = Z;
		19'b1011110010100111010: color_data = Z;
		19'b1011110010100111011: color_data = Z;
		19'b1011110010100111100: color_data = Z;
		19'b1011110010100111101: color_data = Z;
		19'b1011110010100111110: color_data = Z;
		19'b1011110010100111111: color_data = Z;
		19'b1011110010101000000: color_data = Z;
		19'b1011110010101000001: color_data = Z;
		19'b1011110010101000010: color_data = Z;
		19'b1011110010101000011: color_data = Z;
		19'b1011110010101000100: color_data = Z;
		19'b1011110010101000101: color_data = Z;
		19'b1011110010101000110: color_data = Z;
		19'b1011110010101000111: color_data = Z;
		19'b1011110010101001000: color_data = Z;
		19'b1011110010101001001: color_data = Z;
		19'b1011110010101001010: color_data = Z;
		19'b1011110010101001011: color_data = Z;
		19'b1011110010101001100: color_data = Z;
		19'b1011110010101001101: color_data = Z;
		19'b1011110010101001110: color_data = Z;
		19'b1011110010101001111: color_data = Z;
		19'b1011110010101010000: color_data = Z;
		19'b1011110010101010001: color_data = Z;
		19'b1011110010101010010: color_data = Z;
		19'b1011110010101010011: color_data = Z;
		19'b1011110010101010100: color_data = Z;
		19'b1011110010101010101: color_data = Z;
		19'b1011110010101010110: color_data = Z;
		19'b1011110010101010111: color_data = Z;
		19'b1011110010101011000: color_data = Z;
		19'b1011110010101011001: color_data = Z;
		19'b1011110010101011010: color_data = Z;
		19'b1011110010101011011: color_data = Z;
		19'b1011110010101011100: color_data = Z;
		19'b1011110010101011101: color_data = Z;
		19'b1011110010101011110: color_data = Z;
		19'b1011110010101011111: color_data = Z;
		19'b1011110010101100000: color_data = Z;
		19'b1011110010101100001: color_data = Z;
		19'b1011110010101100010: color_data = Z;
		19'b1011110010101100011: color_data = Z;
		19'b1011110010101100100: color_data = Z;
		19'b1011110010101100101: color_data = Z;
		19'b1011110010101100110: color_data = Z;
		19'b1011110010101100111: color_data = Z;
		19'b1011110010101101000: color_data = Z;
		19'b1011110010101101001: color_data = Z;
		19'b1011110010101101010: color_data = Z;
		19'b1011110010101101011: color_data = Z;
		19'b1011110010101101100: color_data = Z;
		19'b1011110010101101101: color_data = Z;
		19'b1011110010101101110: color_data = Z;
		19'b1011110010101101111: color_data = Z;
		19'b1011110010101110000: color_data = Z;
		19'b1011110010101110001: color_data = Z;
		19'b1011110010101110010: color_data = Z;
		19'b1011110010101110011: color_data = Z;
		19'b1011110010101110100: color_data = Z;
		19'b1011110010101110101: color_data = Z;
		19'b1011110010101110110: color_data = Z;
		19'b1011110010101110111: color_data = Z;
		19'b1011110010101111000: color_data = Z;
		19'b1011110010101111001: color_data = Z;
		19'b1011110010101111010: color_data = Z;
		19'b1011110010101111011: color_data = Z;
		19'b1011110010101111100: color_data = Z;
		19'b1011110010101111101: color_data = Z;
		19'b1011110010101111110: color_data = Z;
		19'b1011110010101111111: color_data = Z;
		19'b1011110010110000000: color_data = Z;
		19'b1011110010110000001: color_data = Z;
		19'b1011110010110000010: color_data = Z;
		19'b1011110010110000011: color_data = Z;
		19'b1011110010110000100: color_data = Z;
		19'b1011110010110000101: color_data = Z;
		19'b1011110010110000110: color_data = Z;
		19'b1011110010110000111: color_data = Z;
		19'b1011110100100001000: color_data = Z;
		19'b1011110100100001001: color_data = Z;
		19'b1011110100100001010: color_data = Z;
		19'b1011110100100001011: color_data = Z;
		19'b1011110100100001100: color_data = Z;
		19'b1011110100100001101: color_data = Z;
		19'b1011110100100001110: color_data = Z;
		19'b1011110100100001111: color_data = Z;
		19'b1011110100100010000: color_data = Z;
		19'b1011110100100010001: color_data = Z;
		19'b1011110100100010010: color_data = Z;
		19'b1011110100100010011: color_data = Z;
		19'b1011110100100010100: color_data = Z;
		19'b1011110100100010101: color_data = Z;
		19'b1011110100100010110: color_data = Z;
		19'b1011110100100010111: color_data = Z;
		19'b1011110100100011000: color_data = Z;
		19'b1011110100100011001: color_data = Z;
		19'b1011110100100011010: color_data = Z;
		19'b1011110100100011011: color_data = Z;
		19'b1011110100100011100: color_data = Z;
		19'b1011110100100011101: color_data = Z;
		19'b1011110100100011110: color_data = Z;
		19'b1011110100100011111: color_data = Z;
		19'b1011110100100100000: color_data = Z;
		19'b1011110100100100001: color_data = Z;
		19'b1011110100100100010: color_data = Z;
		19'b1011110100100100011: color_data = Z;
		19'b1011110100100100100: color_data = Z;
		19'b1011110100100100101: color_data = Z;
		19'b1011110100100100110: color_data = Z;
		19'b1011110100100100111: color_data = Z;
		19'b1011110100100101000: color_data = Z;
		19'b1011110100100101001: color_data = Z;
		19'b1011110100100101010: color_data = Z;
		19'b1011110100100101011: color_data = Z;
		19'b1011110100100101100: color_data = Z;
		19'b1011110100100101101: color_data = Z;
		19'b1011110100100101110: color_data = Z;
		19'b1011110100100101111: color_data = Z;
		19'b1011110100100110000: color_data = Z;
		19'b1011110100100110001: color_data = Z;
		19'b1011110100100110010: color_data = Z;
		19'b1011110100100110011: color_data = Z;
		19'b1011110100100110100: color_data = Z;
		19'b1011110100100110101: color_data = Z;
		19'b1011110100100110110: color_data = Z;
		19'b1011110100100110111: color_data = Z;
		19'b1011110100100111000: color_data = Z;
		19'b1011110100100111001: color_data = Z;
		19'b1011110100100111010: color_data = Z;
		19'b1011110100100111011: color_data = Z;
		19'b1011110100100111100: color_data = Z;
		19'b1011110100100111101: color_data = Z;
		19'b1011110100100111110: color_data = Z;
		19'b1011110100100111111: color_data = Z;
		19'b1011110100101000000: color_data = Z;
		19'b1011110100101000001: color_data = Z;
		19'b1011110100101000010: color_data = Z;
		19'b1011110100101000011: color_data = Z;
		19'b1011110100101000100: color_data = Z;
		19'b1011110100101000101: color_data = Z;
		19'b1011110100101000110: color_data = Z;
		19'b1011110100101000111: color_data = Z;
		19'b1011110100101001000: color_data = Z;
		19'b1011110100101001001: color_data = Z;
		19'b1011110100101001010: color_data = Z;
		19'b1011110100101001011: color_data = Z;
		19'b1011110100101001100: color_data = Z;
		19'b1011110100101001101: color_data = Z;
		19'b1011110100101001110: color_data = Z;
		19'b1011110100101001111: color_data = Z;
		19'b1011110100101010000: color_data = Z;
		19'b1011110100101010001: color_data = Z;
		19'b1011110100101010010: color_data = Z;
		19'b1011110100101010011: color_data = Z;
		19'b1011110100101010100: color_data = Z;
		19'b1011110100101010101: color_data = Z;
		19'b1011110100101010110: color_data = Z;
		19'b1011110100101010111: color_data = Z;
		19'b1011110100101011000: color_data = Z;
		19'b1011110100101011001: color_data = Z;
		19'b1011110100101011010: color_data = Z;
		19'b1011110100101011011: color_data = Z;
		19'b1011110100101011100: color_data = Z;
		19'b1011110100101011101: color_data = Z;
		19'b1011110100101011110: color_data = Z;
		19'b1011110100101011111: color_data = Z;
		19'b1011110100101100000: color_data = Z;
		19'b1011110100101100001: color_data = Z;
		19'b1011110100101100010: color_data = Z;
		19'b1011110100101100011: color_data = Z;
		19'b1011110100101100100: color_data = Z;
		19'b1011110100101100101: color_data = Z;
		19'b1011110100101100110: color_data = Z;
		19'b1011110100101100111: color_data = Z;
		19'b1011110100101101000: color_data = Z;
		19'b1011110100101101001: color_data = Z;
		19'b1011110100101101010: color_data = Z;
		19'b1011110100101101011: color_data = Z;
		19'b1011110100101101100: color_data = Z;
		19'b1011110100101101101: color_data = Z;
		19'b1011110100101101110: color_data = Z;
		19'b1011110100101101111: color_data = Z;
		19'b1011110100101110000: color_data = Z;
		19'b1011110100101110001: color_data = Z;
		19'b1011110100101110010: color_data = Z;
		19'b1011110100101110011: color_data = Z;
		19'b1011110100101110100: color_data = Z;
		19'b1011110100101110101: color_data = Z;
		19'b1011110100101110110: color_data = Z;
		19'b1011110100101110111: color_data = Z;
		19'b1011110100101111000: color_data = Z;
		19'b1011110100101111001: color_data = Z;
		19'b1011110100101111010: color_data = Z;
		19'b1011110100101111011: color_data = Z;
		19'b1011110100101111100: color_data = Z;
		19'b1011110100101111101: color_data = Z;
		19'b1011110100101111110: color_data = Z;
		19'b1011110100101111111: color_data = Z;
		19'b1011110100110000000: color_data = Z;
		19'b1011110100110000001: color_data = Z;
		19'b1011110100110000010: color_data = Z;
		19'b1011110100110000011: color_data = Z;
		19'b1011110100110000100: color_data = Z;
		19'b1011110100110000101: color_data = Z;
		19'b1011110100110000110: color_data = Z;
		19'b1011110110100001011: color_data = Z;
		19'b1011110110100001100: color_data = Z;
		19'b1011110110100001101: color_data = Z;
		19'b1011110110100001110: color_data = Z;
		19'b1011110110100001111: color_data = Z;
		19'b1011110110100010000: color_data = Z;
		19'b1011110110100010001: color_data = Z;
		19'b1011110110100010010: color_data = Z;
		19'b1011110110100010011: color_data = Z;
		19'b1011110110100010100: color_data = Z;
		19'b1011110110100010101: color_data = Z;
		19'b1011110110100010110: color_data = Z;
		19'b1011110110100010111: color_data = Z;
		19'b1011110110100011000: color_data = Z;
		19'b1011110110100011001: color_data = Z;
		19'b1011110110100011010: color_data = Z;
		19'b1011110110100011011: color_data = Z;
		19'b1011110110100011100: color_data = Z;
		19'b1011110110100011101: color_data = Z;
		19'b1011110110100011110: color_data = Z;
		19'b1011110110100011111: color_data = Z;
		19'b1011110110100100000: color_data = Z;
		19'b1011110110100100001: color_data = Z;
		19'b1011110110100100010: color_data = Z;
		19'b1011110110100100011: color_data = Z;
		19'b1011110110100100100: color_data = Z;
		19'b1011110110100100101: color_data = Z;
		19'b1011110110100100110: color_data = Z;
		19'b1011110110100100111: color_data = Z;
		19'b1011110110100101000: color_data = Z;
		19'b1011110110100101001: color_data = Z;
		19'b1011110110100101010: color_data = Z;
		19'b1011110110100101011: color_data = Z;
		19'b1011110110100101100: color_data = Z;
		19'b1011110110100101101: color_data = Z;
		19'b1011110110100101110: color_data = Z;
		19'b1011110110100101111: color_data = Z;
		19'b1011110110100110000: color_data = Z;
		19'b1011110110100110001: color_data = Z;
		19'b1011110110100110010: color_data = Z;
		19'b1011110110100110011: color_data = Z;
		19'b1011110110100110100: color_data = Z;
		19'b1011110110100110101: color_data = Z;
		19'b1011110110100110110: color_data = Z;
		19'b1011110110100110111: color_data = Z;
		19'b1011110110100111000: color_data = Z;
		19'b1011110110100111001: color_data = Z;
		19'b1011110110100111010: color_data = Z;
		19'b1011110110100111011: color_data = Z;
		19'b1011110110100111100: color_data = Z;
		19'b1011110110100111101: color_data = Z;
		19'b1011110110100111110: color_data = Z;
		19'b1011110110100111111: color_data = Z;
		19'b1011110110101000000: color_data = Z;
		19'b1011110110101000001: color_data = Z;
		19'b1011110110101000010: color_data = Z;
		19'b1011110110101000011: color_data = Z;
		19'b1011110110101000100: color_data = Z;
		19'b1011110110101000101: color_data = Z;
		19'b1011110110101000110: color_data = Z;
		19'b1011110110101000111: color_data = Z;
		19'b1011110110101001000: color_data = Z;
		19'b1011110110101001001: color_data = Z;
		19'b1011110110101001010: color_data = Z;
		19'b1011110110101001011: color_data = Z;
		19'b1011110110101001100: color_data = Z;
		19'b1011110110101001101: color_data = Z;
		19'b1011110110101001110: color_data = Z;
		19'b1011110110101001111: color_data = Z;
		19'b1011110110101010000: color_data = Z;
		19'b1011110110101010001: color_data = Z;
		19'b1011110110101010010: color_data = Z;
		19'b1011110110101010011: color_data = Z;
		19'b1011110110101010100: color_data = Z;
		19'b1011110110101010101: color_data = Z;
		19'b1011110110101010110: color_data = Z;
		19'b1011110110101010111: color_data = Z;
		19'b1011110110101011000: color_data = Z;
		19'b1011110110101011001: color_data = Z;
		19'b1011110110101011010: color_data = Z;
		19'b1011110110101011011: color_data = Z;
		19'b1011110110101011100: color_data = Z;
		19'b1011110110101011101: color_data = Z;
		19'b1011110110101011110: color_data = Z;
		19'b1011110110101011111: color_data = Z;
		19'b1011110110101100000: color_data = Z;
		19'b1011110110101100001: color_data = Z;
		19'b1011110110101100010: color_data = Z;
		19'b1011110110101100011: color_data = Z;
		19'b1011110110101100100: color_data = Z;
		19'b1011110110101100101: color_data = Z;
		19'b1011110110101100110: color_data = Z;
		19'b1011110110101100111: color_data = Z;
		19'b1011110110101101000: color_data = Z;
		19'b1011110110101101001: color_data = Z;
		19'b1011110110101101010: color_data = Z;
		19'b1011110110101101011: color_data = Z;
		19'b1011110110101101100: color_data = Z;
		19'b1011110110101101101: color_data = Z;
		19'b1011110110101101110: color_data = Z;
		19'b1011110110101101111: color_data = Z;
		19'b1011110110101110000: color_data = Z;
		19'b1011110110101110001: color_data = Z;
		19'b1011110110101110010: color_data = Z;
		19'b1011110110101110011: color_data = Z;
		19'b1011110110101110100: color_data = Z;
		19'b1011110110101110101: color_data = Z;
		19'b1011110110101110110: color_data = Z;
		19'b1011110110101110111: color_data = Z;
		19'b1011110110101111000: color_data = Z;
		19'b1011110110101111001: color_data = Z;
		19'b1011110110101111010: color_data = Z;
		19'b1011110110101111011: color_data = Z;
		19'b1011110110101111100: color_data = Z;
		19'b1011110110101111101: color_data = Z;
		19'b1011110110101111110: color_data = Z;
		19'b1011110110101111111: color_data = Z;
		19'b1011110110110000000: color_data = Z;
		19'b1011110110110000001: color_data = Z;
		19'b1011110110110000010: color_data = Z;
		19'b1011110110110000011: color_data = Z;
		19'b1011110110110000100: color_data = Z;
		19'b1011111000100001110: color_data = Z;
		19'b1011111000100001111: color_data = Z;
		19'b1011111000100010000: color_data = Z;
		19'b1011111000100010001: color_data = Z;
		19'b1011111000100010010: color_data = Z;
		19'b1011111000100010011: color_data = Z;
		19'b1011111000100010100: color_data = Z;
		19'b1011111000100010101: color_data = Z;
		19'b1011111000100010110: color_data = Z;
		19'b1011111000100010111: color_data = Z;
		19'b1011111000100011000: color_data = Z;
		19'b1011111000100011001: color_data = Z;
		19'b1011111000100011010: color_data = Z;
		19'b1011111000100011011: color_data = Z;
		19'b1011111000100011100: color_data = Z;
		19'b1011111000100011101: color_data = Z;
		19'b1011111000100011110: color_data = Z;
		19'b1011111000100011111: color_data = Z;
		19'b1011111000100100000: color_data = Z;
		19'b1011111000100100001: color_data = Z;
		19'b1011111000100100010: color_data = Z;
		19'b1011111000100100011: color_data = Z;
		19'b1011111000100100100: color_data = Z;
		19'b1011111000100100101: color_data = Z;
		19'b1011111000100100110: color_data = Z;
		19'b1011111000100100111: color_data = Z;
		19'b1011111000100101000: color_data = Z;
		19'b1011111000100101001: color_data = Z;
		19'b1011111000100101010: color_data = Z;
		19'b1011111000100101011: color_data = Z;
		19'b1011111000100101100: color_data = Z;
		19'b1011111000100101101: color_data = Z;
		19'b1011111000100101110: color_data = Z;
		19'b1011111000100101111: color_data = Z;
		19'b1011111000100110000: color_data = Z;
		19'b1011111000100110001: color_data = Z;
		19'b1011111000100110010: color_data = Z;
		19'b1011111000100110011: color_data = Z;
		19'b1011111000100110100: color_data = Z;
		19'b1011111000100110101: color_data = Z;
		19'b1011111000100110110: color_data = Z;
		19'b1011111000100110111: color_data = Z;
		19'b1011111000100111000: color_data = Z;
		19'b1011111000100111001: color_data = Z;
		19'b1011111000100111010: color_data = Z;
		19'b1011111000100111011: color_data = Z;
		19'b1011111000100111100: color_data = Z;
		19'b1011111000100111101: color_data = Z;
		19'b1011111000100111110: color_data = Z;
		19'b1011111000100111111: color_data = Z;
		19'b1011111000101000000: color_data = Z;
		19'b1011111000101000001: color_data = Z;
		19'b1011111000101000010: color_data = Z;
		19'b1011111000101000011: color_data = Z;
		19'b1011111000101000100: color_data = Z;
		19'b1011111000101000101: color_data = Z;
		19'b1011111000101000110: color_data = Z;
		19'b1011111000101000111: color_data = Z;
		19'b1011111000101001000: color_data = Z;
		19'b1011111000101001001: color_data = Z;
		19'b1011111000101001010: color_data = Z;
		19'b1011111000101001011: color_data = Z;
		19'b1011111000101001100: color_data = Z;
		19'b1011111000101001101: color_data = Z;
		19'b1011111000101001110: color_data = Z;
		19'b1011111000101001111: color_data = Z;
		19'b1011111000101010000: color_data = Z;
		19'b1011111000101010001: color_data = Z;
		19'b1011111000101010010: color_data = Z;
		19'b1011111000101010011: color_data = Z;
		19'b1011111000101010100: color_data = Z;
		19'b1011111000101010101: color_data = Z;
		19'b1011111000101010110: color_data = Z;
		19'b1011111000101010111: color_data = Z;
		19'b1011111000101011000: color_data = Z;
		19'b1011111000101011001: color_data = Z;
		19'b1011111000101011010: color_data = Z;
		19'b1011111000101011011: color_data = Z;
		19'b1011111000101011100: color_data = Z;
		19'b1011111000101011101: color_data = Z;
		19'b1011111000101011110: color_data = Z;
		19'b1011111000101011111: color_data = Z;
		19'b1011111000101100000: color_data = Z;
		19'b1011111000101100001: color_data = Z;
		19'b1011111000101100010: color_data = Z;
		19'b1011111000101100011: color_data = Z;
		19'b1011111000101100100: color_data = Z;
		19'b1011111000101100101: color_data = Z;
		19'b1011111000101100110: color_data = Z;
		19'b1011111000101100111: color_data = Z;
		19'b1011111000101101000: color_data = Z;
		19'b1011111000101101001: color_data = Z;
		19'b1011111000101101010: color_data = Z;
		19'b1011111000101101011: color_data = Z;
		19'b1011111000101101100: color_data = Z;
		19'b1011111000101101101: color_data = Z;
		19'b1011111000101101110: color_data = Z;
		19'b1011111000101101111: color_data = Z;
		19'b1011111000101110000: color_data = Z;
		19'b1011111000101110001: color_data = Z;
		19'b1011111000101110010: color_data = Z;
		19'b1011111000101110011: color_data = Z;
		19'b1011111000101110100: color_data = Z;
		19'b1011111000101110101: color_data = Z;
		19'b1011111000101110110: color_data = Z;
		19'b1011111000101110111: color_data = Z;
		19'b1011111000101111000: color_data = Z;
		19'b1011111000101111001: color_data = Z;
		19'b1011111000101111010: color_data = Z;
		19'b1011111000101111011: color_data = Z;
		19'b1011111000101111100: color_data = Z;
		19'b1011111000101111101: color_data = Z;
		19'b1011111000101111110: color_data = Z;
		19'b1011111000101111111: color_data = Z;
		19'b1011111000110000000: color_data = Z;
		19'b1011111000110000001: color_data = Z;
		19'b1011111010100010001: color_data = Z;
		19'b1011111010100010010: color_data = Z;
		19'b1011111010100010011: color_data = Z;
		19'b1011111010100010100: color_data = Z;
		19'b1011111010100010101: color_data = Z;
		19'b1011111010100010110: color_data = Z;
		19'b1011111010100010111: color_data = Z;
		19'b1011111010100011000: color_data = Z;
		19'b1011111010100011001: color_data = Z;
		19'b1011111010100011010: color_data = Z;
		19'b1011111010100011011: color_data = Z;
		19'b1011111010100011100: color_data = Z;
		19'b1011111010100011101: color_data = Z;
		19'b1011111010100011110: color_data = Z;
		19'b1011111010100011111: color_data = Z;
		19'b1011111010100100000: color_data = Z;
		19'b1011111010100100001: color_data = Z;
		19'b1011111010100100010: color_data = Z;
		19'b1011111010100100011: color_data = Z;
		19'b1011111010100100100: color_data = Z;
		19'b1011111010100100101: color_data = Z;
		19'b1011111010100100110: color_data = Z;
		19'b1011111010100100111: color_data = Z;
		19'b1011111010100101000: color_data = Z;
		19'b1011111010100101001: color_data = Z;
		19'b1011111010100101010: color_data = Z;
		19'b1011111010100101011: color_data = Z;
		19'b1011111010100101100: color_data = Z;
		19'b1011111010100101101: color_data = Z;
		19'b1011111010100101110: color_data = Z;
		19'b1011111010100101111: color_data = Z;
		19'b1011111010100110000: color_data = Z;
		19'b1011111010100110001: color_data = Z;
		19'b1011111010100110010: color_data = Z;
		19'b1011111010100110011: color_data = Z;
		19'b1011111010100110100: color_data = Z;
		19'b1011111010100110101: color_data = Z;
		19'b1011111010100110110: color_data = Z;
		19'b1011111010100110111: color_data = Z;
		19'b1011111010100111000: color_data = Z;
		19'b1011111010100111001: color_data = Z;
		19'b1011111010100111010: color_data = Z;
		19'b1011111010100111011: color_data = Z;
		19'b1011111010100111100: color_data = Z;
		19'b1011111010100111101: color_data = Z;
		19'b1011111010100111110: color_data = Z;
		19'b1011111010100111111: color_data = Z;
		19'b1011111010101000000: color_data = Z;
		19'b1011111010101000001: color_data = Z;
		19'b1011111010101000010: color_data = Z;
		19'b1011111010101000011: color_data = Z;
		19'b1011111010101000100: color_data = Z;
		19'b1011111010101000101: color_data = Z;
		19'b1011111010101000110: color_data = Z;
		19'b1011111010101000111: color_data = Z;
		19'b1011111010101001000: color_data = Z;
		19'b1011111010101001001: color_data = Z;
		19'b1011111010101001010: color_data = Z;
		19'b1011111010101001011: color_data = Z;
		19'b1011111010101001100: color_data = Z;
		19'b1011111010101001101: color_data = Z;
		19'b1011111010101001110: color_data = Z;
		19'b1011111010101001111: color_data = Z;
		19'b1011111010101010000: color_data = Z;
		19'b1011111010101010001: color_data = Z;
		19'b1011111010101010010: color_data = Z;
		19'b1011111010101010011: color_data = Z;
		19'b1011111010101010100: color_data = Z;
		19'b1011111010101010101: color_data = Z;
		19'b1011111010101010110: color_data = Z;
		19'b1011111010101010111: color_data = Z;
		19'b1011111010101011000: color_data = Z;
		19'b1011111010101011001: color_data = Z;
		19'b1011111010101011010: color_data = Z;
		19'b1011111010101011011: color_data = Z;
		19'b1011111010101011100: color_data = Z;
		19'b1011111010101011101: color_data = Z;
		19'b1011111010101011110: color_data = Z;
		19'b1011111010101011111: color_data = Z;
		19'b1011111010101100000: color_data = Z;
		19'b1011111010101100001: color_data = Z;
		19'b1011111010101100010: color_data = Z;
		19'b1011111010101100011: color_data = Z;
		19'b1011111010101100100: color_data = Z;
		19'b1011111010101100101: color_data = Z;
		19'b1011111010101100110: color_data = Z;
		19'b1011111010101100111: color_data = Z;
		19'b1011111010101101000: color_data = Z;
		19'b1011111010101101001: color_data = Z;
		19'b1011111010101101010: color_data = Z;
		19'b1011111010101101011: color_data = Z;
		19'b1011111010101101100: color_data = Z;
		19'b1011111010101101101: color_data = Z;
		19'b1011111010101101110: color_data = Z;
		19'b1011111010101101111: color_data = Z;
		19'b1011111010101110000: color_data = Z;
		19'b1011111010101110001: color_data = Z;
		19'b1011111010101110010: color_data = Z;
		19'b1011111010101110011: color_data = Z;
		19'b1011111010101110100: color_data = Z;
		19'b1011111010101110101: color_data = Z;
		19'b1011111010101110110: color_data = Z;
		19'b1011111010101110111: color_data = Z;
		19'b1011111010101111000: color_data = Z;
		19'b1011111010101111001: color_data = Z;
		19'b1011111010101111010: color_data = Z;
		19'b1011111010101111011: color_data = Z;
		19'b1011111010101111100: color_data = Z;
		19'b1011111010101111101: color_data = Z;
		19'b1011111010101111110: color_data = Z;
		19'b1011111010101111111: color_data = Z;
		19'b1011111010110000000: color_data = Z;
		19'b1011111100100010011: color_data = Z;
		19'b1011111100100010100: color_data = Z;
		19'b1011111100100010101: color_data = Z;
		19'b1011111100100010110: color_data = Z;
		19'b1011111100100010111: color_data = Z;
		19'b1011111100100011000: color_data = Z;
		19'b1011111100100011001: color_data = Z;
		19'b1011111100100011010: color_data = Z;
		19'b1011111100100011011: color_data = Z;
		19'b1011111100100011100: color_data = Z;
		19'b1011111100100011101: color_data = Z;
		19'b1011111100100011110: color_data = Z;
		19'b1011111100100011111: color_data = Z;
		19'b1011111100100100000: color_data = Z;
		19'b1011111100100100001: color_data = Z;
		19'b1011111100100100010: color_data = Z;
		19'b1011111100100100011: color_data = Z;
		19'b1011111100100100100: color_data = Z;
		19'b1011111100100100101: color_data = Z;
		19'b1011111100100100110: color_data = Z;
		19'b1011111100100100111: color_data = Z;
		19'b1011111100100101000: color_data = Z;
		19'b1011111100100101001: color_data = Z;
		19'b1011111100100101010: color_data = Z;
		19'b1011111100100101011: color_data = Z;
		19'b1011111100100101100: color_data = Z;
		19'b1011111100100101101: color_data = Z;
		19'b1011111100100101110: color_data = Z;
		19'b1011111100100101111: color_data = Z;
		19'b1011111100100110000: color_data = Z;
		19'b1011111100100110001: color_data = Z;
		19'b1011111100100110010: color_data = Z;
		19'b1011111100100110011: color_data = Z;
		19'b1011111100100110100: color_data = Z;
		19'b1011111100100110101: color_data = Z;
		19'b1011111100100110110: color_data = Z;
		19'b1011111100100110111: color_data = Z;
		19'b1011111100100111000: color_data = Z;
		19'b1011111100100111001: color_data = Z;
		19'b1011111100100111010: color_data = Z;
		19'b1011111100100111011: color_data = Z;
		19'b1011111100100111100: color_data = Z;
		19'b1011111100100111101: color_data = Z;
		19'b1011111100100111110: color_data = Z;
		19'b1011111100100111111: color_data = Z;
		19'b1011111100101000000: color_data = Z;
		19'b1011111100101000001: color_data = Z;
		19'b1011111100101000010: color_data = Z;
		19'b1011111100101000011: color_data = Z;
		19'b1011111100101000100: color_data = Z;
		19'b1011111100101000101: color_data = Z;
		19'b1011111100101000110: color_data = Z;
		19'b1011111100101000111: color_data = Z;
		19'b1011111100101001000: color_data = Z;
		19'b1011111100101001001: color_data = Z;
		19'b1011111100101001010: color_data = Z;
		19'b1011111100101001011: color_data = Z;
		19'b1011111100101001100: color_data = Z;
		19'b1011111100101001101: color_data = Z;
		19'b1011111100101001110: color_data = Z;
		19'b1011111100101001111: color_data = Z;
		19'b1011111100101010000: color_data = Z;
		19'b1011111100101010001: color_data = Z;
		19'b1011111100101010010: color_data = Z;
		19'b1011111100101010011: color_data = Z;
		19'b1011111100101010100: color_data = Z;
		19'b1011111100101010101: color_data = Z;
		19'b1011111100101010110: color_data = Z;
		19'b1011111100101010111: color_data = Z;
		19'b1011111100101011000: color_data = Z;
		19'b1011111100101011001: color_data = Z;
		19'b1011111100101011010: color_data = Z;
		19'b1011111100101011011: color_data = Z;
		19'b1011111100101011100: color_data = Z;
		19'b1011111100101011101: color_data = Z;
		19'b1011111100101011110: color_data = Z;
		19'b1011111100101011111: color_data = Z;
		19'b1011111100101100000: color_data = Z;
		19'b1011111100101100001: color_data = Z;
		19'b1011111100101100010: color_data = Z;
		19'b1011111100101100011: color_data = Z;
		19'b1011111100101100100: color_data = Z;
		19'b1011111100101100101: color_data = Z;
		19'b1011111100101100110: color_data = Z;
		19'b1011111100101100111: color_data = Z;
		19'b1011111100101101000: color_data = Z;
		19'b1011111100101101001: color_data = Z;
		19'b1011111100101101010: color_data = Z;
		19'b1011111100101101011: color_data = Z;
		19'b1011111100101101100: color_data = Z;
		19'b1011111100101101101: color_data = Z;
		19'b1011111100101101110: color_data = Z;
		19'b1011111100101101111: color_data = Z;
		19'b1011111100101110000: color_data = Z;
		19'b1011111100101110001: color_data = Z;
		19'b1011111100101110010: color_data = Z;
		19'b1011111100101110011: color_data = Z;
		19'b1011111100101110100: color_data = Z;
		19'b1011111100101110101: color_data = Z;
		19'b1011111100101110110: color_data = Z;
		19'b1011111100101110111: color_data = Z;
		19'b1011111100101111000: color_data = Z;
		19'b1011111100101111001: color_data = Z;
		19'b1011111100101111010: color_data = Z;
		19'b1011111100101111011: color_data = Z;
		19'b1011111100101111100: color_data = Z;
		19'b1011111100101111101: color_data = Z;
		19'b1011111100101111110: color_data = Z;
		19'b1011111100101111111: color_data = Z;
		19'b1011111110100010100: color_data = Z;
		19'b1011111110100010101: color_data = Z;
		19'b1011111110100010110: color_data = Z;
		19'b1011111110100010111: color_data = Z;
		19'b1011111110100011000: color_data = Z;
		19'b1011111110100011001: color_data = Z;
		19'b1011111110100011010: color_data = Z;
		19'b1011111110100011011: color_data = Z;
		19'b1011111110100011100: color_data = Z;
		19'b1011111110100011101: color_data = Z;
		19'b1011111110100011110: color_data = Z;
		19'b1011111110100011111: color_data = Z;
		19'b1011111110100100000: color_data = Z;
		19'b1011111110100100001: color_data = Z;
		19'b1011111110100100010: color_data = Z;
		19'b1011111110100100011: color_data = Z;
		19'b1011111110100100100: color_data = Z;
		19'b1011111110100100101: color_data = Z;
		19'b1011111110100100110: color_data = Z;
		19'b1011111110100100111: color_data = Z;
		19'b1011111110100101000: color_data = Z;
		19'b1011111110100101001: color_data = Z;
		19'b1011111110100101010: color_data = Z;
		19'b1011111110100101011: color_data = Z;
		19'b1011111110100101100: color_data = Z;
		19'b1011111110100101101: color_data = Z;
		19'b1011111110100101110: color_data = Z;
		19'b1011111110100101111: color_data = Z;
		19'b1011111110100110000: color_data = Z;
		19'b1011111110100110001: color_data = Z;
		19'b1011111110100110010: color_data = Z;
		19'b1011111110100110011: color_data = Z;
		19'b1011111110100110100: color_data = Z;
		19'b1011111110100110101: color_data = Z;
		19'b1011111110100110110: color_data = Z;
		19'b1011111110100110111: color_data = Z;
		19'b1011111110100111000: color_data = Z;
		19'b1011111110100111001: color_data = Z;
		19'b1011111110100111010: color_data = Z;
		19'b1011111110100111011: color_data = Z;
		19'b1011111110100111100: color_data = Z;
		19'b1011111110100111101: color_data = Z;
		19'b1011111110100111110: color_data = Z;
		19'b1011111110100111111: color_data = Z;
		19'b1011111110101000000: color_data = Z;
		19'b1011111110101000001: color_data = Z;
		19'b1011111110101000010: color_data = Z;
		19'b1011111110101000011: color_data = Z;
		19'b1011111110101000100: color_data = Z;
		19'b1011111110101000101: color_data = Z;
		19'b1011111110101000110: color_data = Z;
		19'b1011111110101000111: color_data = Z;
		19'b1011111110101001000: color_data = Z;
		19'b1011111110101001001: color_data = Z;
		19'b1011111110101001010: color_data = Z;
		19'b1011111110101001011: color_data = Z;
		19'b1011111110101001100: color_data = Z;
		19'b1011111110101001101: color_data = Z;
		19'b1011111110101001110: color_data = Z;
		19'b1011111110101001111: color_data = Z;
		19'b1011111110101010000: color_data = Z;
		19'b1011111110101010001: color_data = Z;
		19'b1011111110101010010: color_data = Z;
		19'b1011111110101010011: color_data = Z;
		19'b1011111110101010100: color_data = Z;
		19'b1011111110101010101: color_data = Z;
		19'b1011111110101010110: color_data = Z;
		19'b1011111110101010111: color_data = Z;
		19'b1011111110101011000: color_data = Z;
		19'b1011111110101011001: color_data = Z;
		19'b1011111110101011010: color_data = Z;
		19'b1011111110101011011: color_data = Z;
		19'b1011111110101011100: color_data = Z;
		19'b1011111110101011101: color_data = Z;
		19'b1011111110101011110: color_data = Z;
		19'b1011111110101011111: color_data = Z;
		19'b1011111110101100000: color_data = Z;
		19'b1011111110101100001: color_data = Z;
		19'b1011111110101100010: color_data = Z;
		19'b1011111110101100011: color_data = Z;
		19'b1011111110101100100: color_data = Z;
		19'b1011111110101100101: color_data = Z;
		19'b1011111110101100110: color_data = Z;
		19'b1011111110101100111: color_data = Z;
		19'b1011111110101101000: color_data = Z;
		19'b1011111110101101001: color_data = Z;
		19'b1011111110101101010: color_data = Z;
		19'b1011111110101101011: color_data = Z;
		19'b1011111110101101100: color_data = Z;
		19'b1011111110101101101: color_data = Z;
		19'b1011111110101101110: color_data = Z;
		19'b1011111110101101111: color_data = Z;
		19'b1011111110101110000: color_data = Z;
		19'b1011111110101110001: color_data = Z;
		19'b1011111110101110010: color_data = Z;
		19'b1011111110101110011: color_data = Z;
		19'b1011111110101110100: color_data = Z;
		19'b1011111110101110101: color_data = Z;
		19'b1011111110101110110: color_data = Z;
		19'b1011111110101110111: color_data = Z;
		19'b1011111110101111000: color_data = Z;
		19'b1011111110101111001: color_data = Z;
		19'b1011111110101111010: color_data = Z;
		19'b1011111110101111011: color_data = Z;
		19'b1011111110101111100: color_data = Z;
		19'b1011111110101111101: color_data = Z;
		19'b1011111110101111110: color_data = Z;
		19'b1100000000100010110: color_data = Z;
		19'b1100000000100010111: color_data = Z;
		19'b1100000000100011000: color_data = Z;
		19'b1100000000100011001: color_data = Z;
		19'b1100000000100011010: color_data = Z;
		19'b1100000000100011011: color_data = Z;
		19'b1100000000100011100: color_data = Z;
		19'b1100000000100011101: color_data = Z;
		19'b1100000000100011110: color_data = Z;
		19'b1100000000100011111: color_data = Z;
		19'b1100000000100100000: color_data = Z;
		19'b1100000000100100001: color_data = Z;
		19'b1100000000100100010: color_data = Z;
		19'b1100000000100100011: color_data = Z;
		19'b1100000000100100100: color_data = Z;
		19'b1100000000100100101: color_data = Z;
		19'b1100000000100100110: color_data = Z;
		19'b1100000000100100111: color_data = Z;
		19'b1100000000100101000: color_data = Z;
		19'b1100000000100101001: color_data = Z;
		19'b1100000000100101010: color_data = Z;
		19'b1100000000100101011: color_data = Z;
		19'b1100000000100101100: color_data = Z;
		19'b1100000000100101101: color_data = Z;
		19'b1100000000100101110: color_data = Z;
		19'b1100000000100101111: color_data = Z;
		19'b1100000000100110000: color_data = Z;
		19'b1100000000100110001: color_data = Z;
		19'b1100000000100110010: color_data = Z;
		19'b1100000000100110011: color_data = Z;
		19'b1100000000100110100: color_data = Z;
		19'b1100000000100110101: color_data = Z;
		19'b1100000000100110110: color_data = Z;
		19'b1100000000100110111: color_data = Z;
		19'b1100000000100111000: color_data = Z;
		19'b1100000000100111001: color_data = Z;
		19'b1100000000100111010: color_data = Z;
		19'b1100000000100111011: color_data = Z;
		19'b1100000000100111100: color_data = Z;
		19'b1100000000100111101: color_data = Z;
		19'b1100000000100111110: color_data = Z;
		19'b1100000000100111111: color_data = Z;
		19'b1100000000101000000: color_data = Z;
		19'b1100000000101000001: color_data = Z;
		19'b1100000000101000010: color_data = Z;
		19'b1100000000101000011: color_data = Z;
		19'b1100000000101000100: color_data = Z;
		19'b1100000000101000101: color_data = Z;
		19'b1100000000101000110: color_data = Z;
		19'b1100000000101000111: color_data = Z;
		19'b1100000000101001000: color_data = Z;
		19'b1100000000101001001: color_data = Z;
		19'b1100000000101001010: color_data = Z;
		19'b1100000000101001011: color_data = Z;
		19'b1100000000101001100: color_data = Z;
		19'b1100000000101001101: color_data = Z;
		19'b1100000000101001110: color_data = Z;
		19'b1100000000101001111: color_data = Z;
		19'b1100000000101010000: color_data = Z;
		19'b1100000000101010001: color_data = Z;
		19'b1100000000101010010: color_data = Z;
		19'b1100000000101010011: color_data = Z;
		19'b1100000000101010100: color_data = Z;
		19'b1100000000101010101: color_data = Z;
		19'b1100000000101010110: color_data = Z;
		19'b1100000000101010111: color_data = Z;
		19'b1100000000101011111: color_data = Z;
		19'b1100000000101100001: color_data = Z;
		19'b1100000000101100010: color_data = Z;
		19'b1100000000101100011: color_data = Z;
		19'b1100000000101100100: color_data = Z;
		19'b1100000000101100101: color_data = Z;
		19'b1100000000101100110: color_data = Z;
		19'b1100000000101100111: color_data = Z;
		19'b1100000000101101000: color_data = Z;
		19'b1100000000101101001: color_data = Z;
		19'b1100000000101101010: color_data = Z;
		19'b1100000000101101011: color_data = Z;
		19'b1100000000101101100: color_data = Z;
		19'b1100000000101101101: color_data = Z;
		19'b1100000000101101110: color_data = Z;
		19'b1100000000101101111: color_data = Z;
		19'b1100000000101110000: color_data = Z;
		19'b1100000000101110001: color_data = Z;
		19'b1100000000101110010: color_data = Z;
		19'b1100000000101110011: color_data = Z;
		19'b1100000000101110100: color_data = Z;
		19'b1100000000101110101: color_data = Z;
		19'b1100000000101110110: color_data = Z;
		19'b1100000000101110111: color_data = Z;
		19'b1100000000101111000: color_data = Z;
		19'b1100000000101111001: color_data = Z;
		19'b1100000000101111010: color_data = Z;
		19'b1100000000101111011: color_data = Z;
		19'b1100000000101111100: color_data = Z;
		19'b1100000000101111101: color_data = Z;
		19'b1100000010100011001: color_data = Z;
		19'b1100000010100011010: color_data = Z;
		19'b1100000010100011011: color_data = Z;
		19'b1100000010100011100: color_data = Z;
		19'b1100000010100011101: color_data = Z;
		19'b1100000010100011110: color_data = Z;
		19'b1100000010100011111: color_data = Z;
		19'b1100000010100100000: color_data = Z;
		19'b1100000010100100001: color_data = Z;
		19'b1100000010100100010: color_data = Z;
		19'b1100000010100100011: color_data = Z;
		19'b1100000010100100100: color_data = Z;
		19'b1100000010100100101: color_data = Z;
		19'b1100000010100100110: color_data = Z;
		19'b1100000010100100111: color_data = Z;
		19'b1100000010100101000: color_data = Z;
		19'b1100000010100101001: color_data = Z;
		19'b1100000010100101010: color_data = Z;
		19'b1100000010100101011: color_data = Z;
		19'b1100000010100101100: color_data = Z;
		19'b1100000010100101101: color_data = Z;
		19'b1100000010100101110: color_data = Z;
		19'b1100000010100101111: color_data = Z;
		19'b1100000010100110000: color_data = Z;
		19'b1100000010100110001: color_data = Z;
		19'b1100000010100110010: color_data = Z;
		19'b1100000010100110011: color_data = Z;
		19'b1100000010100110100: color_data = Z;
		19'b1100000010100110101: color_data = Z;
		19'b1100000010100110110: color_data = Z;
		19'b1100000010100110111: color_data = Z;
		19'b1100000010100111000: color_data = Z;
		19'b1100000010100111001: color_data = Z;
		19'b1100000010100111010: color_data = Z;
		19'b1100000010100111011: color_data = Z;
		19'b1100000010100111100: color_data = Z;
		19'b1100000010100111101: color_data = Z;
		19'b1100000010100111110: color_data = Z;
		19'b1100000010100111111: color_data = Z;
		19'b1100000010101000000: color_data = Z;
		19'b1100000010101000001: color_data = Z;
		19'b1100000010101000010: color_data = Z;
		19'b1100000010101000011: color_data = Z;
		19'b1100000010101000100: color_data = Z;
		19'b1100000010101000101: color_data = Z;
		19'b1100000010101000110: color_data = Z;
		19'b1100000010101000111: color_data = Z;
		19'b1100000010101001000: color_data = Z;
		19'b1100000010101001001: color_data = Z;
		19'b1100000010101001010: color_data = Z;
		19'b1100000010101001011: color_data = Z;
		19'b1100000010101001100: color_data = Z;
		19'b1100000010101001101: color_data = Z;
		19'b1100000010101001110: color_data = Z;
		19'b1100000010101001111: color_data = Z;
		19'b1100000010101010000: color_data = Z;
		19'b1100000010101010001: color_data = Z;
		19'b1100000010101010010: color_data = Z;
		19'b1100000010101010011: color_data = Z;
		19'b1100000010101010100: color_data = Z;
		19'b1100000010101010101: color_data = Z;
		19'b1100000010101010110: color_data = Z;
		19'b1100000010101010111: color_data = Z;
		19'b1100000010101011100: color_data = Z;
		19'b1100000010101011101: color_data = Z;
		19'b1100000010101011110: color_data = Z;
		19'b1100000010101011111: color_data = Z;
		19'b1100000010101100000: color_data = Z;
		19'b1100000010101100001: color_data = Z;
		19'b1100000010101100010: color_data = Z;
		19'b1100000010101100011: color_data = Z;
		19'b1100000010101100100: color_data = Z;
		19'b1100000010101100101: color_data = Z;
		19'b1100000010101100110: color_data = Z;
		19'b1100000010101100111: color_data = Z;
		19'b1100000010101101000: color_data = Z;
		19'b1100000010101101001: color_data = Z;
		19'b1100000010101101010: color_data = Z;
		19'b1100000010101101011: color_data = Z;
		19'b1100000010101101100: color_data = Z;
		19'b1100000010101101101: color_data = Z;
		19'b1100000010101101110: color_data = Z;
		19'b1100000010101101111: color_data = Z;
		19'b1100000010101110000: color_data = Z;
		19'b1100000010101110001: color_data = Z;
		19'b1100000010101110010: color_data = Z;
		19'b1100000010101110011: color_data = Z;
		19'b1100000010101110100: color_data = Z;
		19'b1100000010101110101: color_data = Z;
		19'b1100000010101110110: color_data = Z;
		19'b1100000010101110111: color_data = Z;
		19'b1100000010101111000: color_data = Z;
		19'b1100000010101111001: color_data = Z;
		19'b1100000010101111010: color_data = Z;
		19'b1100000010101111011: color_data = Z;
		19'b1100000010101111100: color_data = Z;
		19'b1100000010101111101: color_data = Z;
		19'b1100000100100011100: color_data = Z;
		19'b1100000100100011101: color_data = Z;
		19'b1100000100100011110: color_data = Z;
		19'b1100000100100011111: color_data = Z;
		19'b1100000100100100000: color_data = Z;
		19'b1100000100100100001: color_data = Z;
		19'b1100000100100100010: color_data = Z;
		19'b1100000100100100011: color_data = Z;
		19'b1100000100100100100: color_data = Z;
		19'b1100000100100100101: color_data = Z;
		19'b1100000100100100110: color_data = Z;
		19'b1100000100100100111: color_data = Z;
		19'b1100000100100101000: color_data = Z;
		19'b1100000100100101001: color_data = Z;
		19'b1100000100100101010: color_data = Z;
		19'b1100000100100101011: color_data = Z;
		19'b1100000100100101100: color_data = Z;
		19'b1100000100100101101: color_data = Z;
		19'b1100000100100101110: color_data = Z;
		19'b1100000100100101111: color_data = Z;
		19'b1100000100100110000: color_data = Z;
		19'b1100000100100110001: color_data = Z;
		19'b1100000100100110010: color_data = Z;
		19'b1100000100100110011: color_data = Z;
		19'b1100000100100110100: color_data = Z;
		19'b1100000100100110101: color_data = Z;
		19'b1100000100100110110: color_data = Z;
		19'b1100000100100110111: color_data = Z;
		19'b1100000100100111000: color_data = Z;
		19'b1100000100100111001: color_data = Z;
		19'b1100000100100111010: color_data = Z;
		19'b1100000100100111011: color_data = Z;
		19'b1100000100100111100: color_data = Z;
		19'b1100000100100111101: color_data = Z;
		19'b1100000100100111110: color_data = Z;
		19'b1100000100100111111: color_data = Z;
		19'b1100000100101000000: color_data = Z;
		19'b1100000100101000001: color_data = Z;
		19'b1100000100101000010: color_data = Z;
		19'b1100000100101000011: color_data = Z;
		19'b1100000100101000100: color_data = Z;
		19'b1100000100101000101: color_data = Z;
		19'b1100000100101000110: color_data = Z;
		19'b1100000100101000111: color_data = Z;
		19'b1100000100101001000: color_data = Z;
		19'b1100000100101001001: color_data = Z;
		19'b1100000100101001010: color_data = Z;
		19'b1100000100101001011: color_data = Z;
		19'b1100000100101001100: color_data = Z;
		19'b1100000100101001101: color_data = Z;
		19'b1100000100101001110: color_data = Z;
		19'b1100000100101001111: color_data = Z;
		19'b1100000100101010000: color_data = Z;
		19'b1100000100101010001: color_data = Z;
		19'b1100000100101010010: color_data = Z;
		19'b1100000100101010011: color_data = Z;
		19'b1100000100101010100: color_data = Z;
		19'b1100000100101010101: color_data = Z;
		19'b1100000100101010110: color_data = Z;
		19'b1100000100101010111: color_data = Z;
		19'b1100000100101011000: color_data = Z;
		19'b1100000100101011001: color_data = Z;
		19'b1100000100101011010: color_data = Z;
		19'b1100000100101011011: color_data = Z;
		19'b1100000100101011100: color_data = Z;
		19'b1100000100101011101: color_data = Z;
		19'b1100000100101011110: color_data = Z;
		19'b1100000100101011111: color_data = Z;
		19'b1100000100101100000: color_data = Z;
		19'b1100000100101100001: color_data = Z;
		19'b1100000100101100010: color_data = Z;
		19'b1100000100101100011: color_data = Z;
		19'b1100000100101100100: color_data = Z;
		19'b1100000100101100101: color_data = Z;
		19'b1100000100101100110: color_data = Z;
		19'b1100000100101100111: color_data = Z;
		19'b1100000100101101000: color_data = Z;
		19'b1100000100101101001: color_data = Z;
		19'b1100000100101101010: color_data = Z;
		19'b1100000100101101011: color_data = Z;
		19'b1100000100101101100: color_data = Z;
		19'b1100000100101101101: color_data = Z;
		19'b1100000100101101110: color_data = Z;
		19'b1100000100101101111: color_data = Z;
		19'b1100000100101110000: color_data = Z;
		19'b1100000100101110001: color_data = Z;
		19'b1100000100101110010: color_data = Z;
		19'b1100000100101110011: color_data = Z;
		19'b1100000100101110100: color_data = Z;
		19'b1100000100101110101: color_data = Z;
		19'b1100000100101110110: color_data = Z;
		19'b1100000100101110111: color_data = Z;
		19'b1100000100101111000: color_data = Z;
		19'b1100000100101111001: color_data = Z;
		19'b1100000100101111010: color_data = Z;
		19'b1100000100101111011: color_data = Z;
		19'b1100000110100100000: color_data = Z;
		19'b1100000110100100001: color_data = Z;
		19'b1100000110100100010: color_data = Z;
		19'b1100000110100100011: color_data = Z;
		19'b1100000110100100100: color_data = Z;
		19'b1100000110100100101: color_data = Z;
		19'b1100000110100100110: color_data = Z;
		19'b1100000110100100111: color_data = Z;
		19'b1100000110100101000: color_data = Z;
		19'b1100000110100101001: color_data = Z;
		19'b1100000110100101010: color_data = Z;
		19'b1100000110100101011: color_data = Z;
		19'b1100000110100101100: color_data = Z;
		19'b1100000110100101101: color_data = Z;
		19'b1100000110100101110: color_data = Z;
		19'b1100000110100101111: color_data = Z;
		19'b1100000110100110000: color_data = Z;
		19'b1100000110100110001: color_data = Z;
		19'b1100000110100110010: color_data = Z;
		19'b1100000110100110011: color_data = Z;
		19'b1100000110100110100: color_data = Z;
		19'b1100000110100110101: color_data = Z;
		19'b1100000110100110110: color_data = Z;
		19'b1100000110100110111: color_data = Z;
		19'b1100000110100111000: color_data = Z;
		19'b1100000110100111001: color_data = Z;
		19'b1100000110100111010: color_data = Z;
		19'b1100000110100111011: color_data = Z;
		19'b1100000110100111100: color_data = Z;
		19'b1100000110100111101: color_data = Z;
		19'b1100000110100111110: color_data = Z;
		19'b1100000110100111111: color_data = Z;
		19'b1100000110101000000: color_data = Z;
		19'b1100000110101000001: color_data = Z;
		19'b1100000110101000010: color_data = Z;
		19'b1100000110101000011: color_data = Z;
		19'b1100000110101000100: color_data = Z;
		19'b1100000110101000101: color_data = Z;
		19'b1100000110101000110: color_data = Z;
		19'b1100000110101000111: color_data = Z;
		19'b1100000110101001000: color_data = Z;
		19'b1100000110101001001: color_data = Z;
		19'b1100000110101001010: color_data = Z;
		19'b1100000110101001011: color_data = Z;
		19'b1100000110101001100: color_data = Z;
		19'b1100000110101001101: color_data = Z;
		19'b1100000110101001110: color_data = Z;
		19'b1100000110101001111: color_data = Z;
		19'b1100000110101010000: color_data = Z;
		19'b1100000110101010001: color_data = Z;
		19'b1100000110101010010: color_data = Z;
		19'b1100000110101010011: color_data = Z;
		19'b1100000110101010100: color_data = Z;
		19'b1100000110101010101: color_data = Z;
		19'b1100000110101010110: color_data = Z;
		19'b1100000110101010111: color_data = Z;
		19'b1100000110101011000: color_data = Z;
		19'b1100000110101011001: color_data = Z;
		19'b1100000110101011010: color_data = Z;
		19'b1100000110101011011: color_data = Z;
		19'b1100000110101011100: color_data = Z;
		19'b1100000110101011101: color_data = Z;
		19'b1100000110101011110: color_data = Z;
		19'b1100000110101011111: color_data = Z;
		19'b1100000110101100000: color_data = Z;
		19'b1100000110101100001: color_data = Z;
		19'b1100000110101100010: color_data = Z;
		19'b1100000110101100011: color_data = Z;
		19'b1100000110101100100: color_data = Z;
		19'b1100000110101100101: color_data = Z;
		19'b1100000110101100110: color_data = Z;
		19'b1100000110101100111: color_data = Z;
		19'b1100000110101101000: color_data = Z;
		19'b1100000110101101001: color_data = Z;
		19'b1100000110101101010: color_data = Z;
		19'b1100000110101101011: color_data = Z;
		19'b1100000110101101100: color_data = Z;
		19'b1100000110101101101: color_data = Z;
		19'b1100000110101101110: color_data = Z;
		19'b1100000110101101111: color_data = Z;
		19'b1100000110101110000: color_data = Z;
		19'b1100000110101110001: color_data = Z;
		19'b1100000110101110010: color_data = Z;
		19'b1100000110101110011: color_data = Z;
		19'b1100000110101110100: color_data = Z;
		19'b1100000110101110101: color_data = Z;
		19'b1100000110101110110: color_data = Z;
		19'b1100000110101110111: color_data = Z;
		19'b1100000110101111000: color_data = Z;
		19'b1100000110101111001: color_data = Z;
		19'b1100000110101111010: color_data = Z;
		19'b1100001000100100010: color_data = Z;
		19'b1100001000100100011: color_data = Z;
		19'b1100001000100100100: color_data = Z;
		19'b1100001000100100101: color_data = Z;
		19'b1100001000100100110: color_data = Z;
		19'b1100001000100100111: color_data = Z;
		19'b1100001000100101000: color_data = Z;
		19'b1100001000100101001: color_data = Z;
		19'b1100001000100101010: color_data = Z;
		19'b1100001000100101011: color_data = Z;
		19'b1100001000100101100: color_data = Z;
		19'b1100001000100101101: color_data = Z;
		19'b1100001000100101110: color_data = Z;
		19'b1100001000100101111: color_data = Z;
		19'b1100001000100110000: color_data = Z;
		19'b1100001000100110001: color_data = Z;
		19'b1100001000100110010: color_data = Z;
		19'b1100001000100110011: color_data = Z;
		19'b1100001000100110100: color_data = Z;
		19'b1100001000100110101: color_data = Z;
		19'b1100001000100110110: color_data = Z;
		19'b1100001000100110111: color_data = Z;
		19'b1100001000100111000: color_data = Z;
		19'b1100001000100111001: color_data = Z;
		19'b1100001000100111010: color_data = Z;
		19'b1100001000100111011: color_data = Z;
		19'b1100001000100111100: color_data = Z;
		19'b1100001000100111101: color_data = Z;
		19'b1100001000100111110: color_data = Z;
		19'b1100001000100111111: color_data = Z;
		19'b1100001000101000000: color_data = Z;
		19'b1100001000101000001: color_data = Z;
		19'b1100001000101000010: color_data = Z;
		19'b1100001000101000011: color_data = Z;
		19'b1100001000101000100: color_data = Z;
		19'b1100001000101000101: color_data = Z;
		19'b1100001000101000110: color_data = Z;
		19'b1100001000101000111: color_data = Z;
		19'b1100001000101001000: color_data = Z;
		19'b1100001000101001001: color_data = Z;
		19'b1100001000101001010: color_data = Z;
		19'b1100001000101001011: color_data = Z;
		19'b1100001000101011111: color_data = Z;
		19'b1100001000101100000: color_data = Z;
		19'b1100001000101100001: color_data = Z;
		19'b1100001000101100010: color_data = Z;
		19'b1100001000101100011: color_data = Z;
		19'b1100001000101100100: color_data = Z;
		19'b1100001000101100101: color_data = Z;
		19'b1100001000101100110: color_data = Z;
		19'b1100001000101100111: color_data = Z;
		19'b1100001000101101000: color_data = Z;
		19'b1100001000101101001: color_data = Z;
		19'b1100001000101101010: color_data = Z;
		19'b1100001000101101011: color_data = Z;
		19'b1100001000101101100: color_data = Z;
		19'b1100001000101101101: color_data = Z;
		19'b1100001000101101110: color_data = Z;
		19'b1100001000101101111: color_data = Z;
		19'b1100001000101110000: color_data = Z;
		19'b1100001000101110001: color_data = Z;
		19'b1100001000101110010: color_data = Z;
		19'b1100001000101110011: color_data = Z;
		19'b1100001000101110100: color_data = Z;
		19'b1100001000101110101: color_data = Z;
		19'b1100001000101110110: color_data = Z;
		19'b1100001000101110111: color_data = Z;
		19'b1100001000101111000: color_data = Z;
		19'b1100001000101111001: color_data = Z;
		19'b1100001010100100100: color_data = Z;
		19'b1100001010100100101: color_data = Z;
		19'b1100001010100100110: color_data = Z;
		19'b1100001010100100111: color_data = Z;
		19'b1100001010100101000: color_data = Z;
		19'b1100001010100101001: color_data = Z;
		19'b1100001010100101010: color_data = Z;
		19'b1100001010100101011: color_data = Z;
		19'b1100001010100101100: color_data = Z;
		19'b1100001010100101101: color_data = Z;
		19'b1100001010100101110: color_data = Z;
		19'b1100001010100101111: color_data = Z;
		19'b1100001010100110000: color_data = Z;
		19'b1100001010100110001: color_data = Z;
		19'b1100001010100110010: color_data = Z;
		19'b1100001010100110011: color_data = Z;
		19'b1100001010100110100: color_data = Z;
		19'b1100001010100110101: color_data = Z;
		19'b1100001010100110110: color_data = Z;
		19'b1100001010100110111: color_data = Z;
		19'b1100001010100111000: color_data = Z;
		19'b1100001010100111001: color_data = Z;
		19'b1100001010100111010: color_data = Z;
		19'b1100001010100111011: color_data = Z;
		19'b1100001010100111100: color_data = Z;
		19'b1100001010100111101: color_data = Z;
		19'b1100001010100111110: color_data = Z;
		19'b1100001010100111111: color_data = Z;
		19'b1100001010101000000: color_data = Z;
		19'b1100001010101000001: color_data = Z;
		19'b1100001010101000010: color_data = Z;
		19'b1100001010101000011: color_data = Z;
		19'b1100001010101000100: color_data = Z;
		19'b1100001010101000101: color_data = Z;
		19'b1100001010101000110: color_data = Z;
		19'b1100001010101000111: color_data = Z;
		19'b1100001010101001000: color_data = Z;
		19'b1100001010101001001: color_data = Z;
		19'b1100001010101011111: color_data = Z;
		19'b1100001010101100010: color_data = Z;
		19'b1100001010101100011: color_data = Z;
		19'b1100001010101100100: color_data = Z;
		19'b1100001010101100101: color_data = Z;
		19'b1100001010101100110: color_data = Z;
		19'b1100001010101100111: color_data = Z;
		19'b1100001010101101000: color_data = Z;
		19'b1100001010101101001: color_data = Z;
		19'b1100001010101101010: color_data = Z;
		19'b1100001010101101011: color_data = Z;
		19'b1100001010101101100: color_data = Z;
		19'b1100001010101101101: color_data = Z;
		19'b1100001010101101110: color_data = Z;
		19'b1100001010101101111: color_data = Z;
		19'b1100001010101110000: color_data = Z;
		19'b1100001010101110001: color_data = Z;
		19'b1100001010101110010: color_data = Z;
		19'b1100001010101110011: color_data = Z;
		19'b1100001010101110100: color_data = Z;
		19'b1100001010101110101: color_data = Z;
		19'b1100001010101110110: color_data = Z;
		19'b1100001010101110111: color_data = Z;
		19'b1100001010101111000: color_data = Z;
		19'b1100001100100100101: color_data = Z;
		19'b1100001100100100110: color_data = Z;
		19'b1100001100100100111: color_data = Z;
		19'b1100001100100101000: color_data = Z;
		19'b1100001100100101001: color_data = Z;
		19'b1100001100100101010: color_data = Z;
		19'b1100001100100101011: color_data = Z;
		19'b1100001100100101100: color_data = Z;
		19'b1100001100100101101: color_data = Z;
		19'b1100001100100101110: color_data = Z;
		19'b1100001100100101111: color_data = Z;
		19'b1100001100100110000: color_data = Z;
		19'b1100001100100110001: color_data = Z;
		19'b1100001100100110010: color_data = Z;
		19'b1100001100100110011: color_data = Z;
		19'b1100001100100110100: color_data = Z;
		19'b1100001100100110101: color_data = Z;
		19'b1100001100100110110: color_data = Z;
		19'b1100001100100110111: color_data = Z;
		19'b1100001100100111000: color_data = Z;
		19'b1100001100100111001: color_data = Z;
		19'b1100001100100111010: color_data = Z;
		19'b1100001100100111011: color_data = Z;
		19'b1100001100100111100: color_data = Z;
		19'b1100001100100111101: color_data = Z;
		19'b1100001100100111110: color_data = Z;
		19'b1100001100100111111: color_data = Z;
		19'b1100001100101000000: color_data = Z;
		19'b1100001100101000001: color_data = Z;
		19'b1100001100101000010: color_data = Z;
		19'b1100001100101000011: color_data = Z;
		19'b1100001100101000100: color_data = Z;
		19'b1100001100101000101: color_data = Z;
		19'b1100001100101000110: color_data = Z;
		19'b1100001100101000111: color_data = Z;
		19'b1100001100101001000: color_data = Z;
		19'b1100001100101001001: color_data = Z;
		19'b1100001100101100000: color_data = Z;
		19'b1100001100101100001: color_data = Z;
		19'b1100001100101100010: color_data = Z;
		19'b1100001100101100011: color_data = Z;
		19'b1100001100101100100: color_data = Z;
		19'b1100001100101100101: color_data = Z;
		19'b1100001100101100110: color_data = Z;
		19'b1100001100101100111: color_data = Z;
		19'b1100001100101101000: color_data = Z;
		19'b1100001100101101001: color_data = Z;
		19'b1100001100101101010: color_data = Z;
		19'b1100001100101101011: color_data = Z;
		19'b1100001100101101100: color_data = Z;
		19'b1100001100101101101: color_data = Z;
		19'b1100001100101101110: color_data = Z;
		19'b1100001100101101111: color_data = Z;
		19'b1100001100101110000: color_data = Z;
		19'b1100001100101110001: color_data = Z;
		19'b1100001100101110010: color_data = Z;
		19'b1100001100101110011: color_data = Z;
		19'b1100001100101110100: color_data = Z;
		19'b1100001100101110101: color_data = Z;
		19'b1100001100101110110: color_data = Z;
		19'b1100001100101110111: color_data = Z;
		19'b1100001110100100110: color_data = Z;
		19'b1100001110100100111: color_data = Z;
		19'b1100001110100101000: color_data = Z;
		19'b1100001110100101001: color_data = Z;
		19'b1100001110100101010: color_data = Z;
		19'b1100001110100101011: color_data = Z;
		19'b1100001110100101100: color_data = Z;
		19'b1100001110100101101: color_data = Z;
		19'b1100001110100101110: color_data = Z;
		19'b1100001110100101111: color_data = Z;
		19'b1100001110100110000: color_data = Z;
		19'b1100001110100110001: color_data = Z;
		19'b1100001110100110010: color_data = Z;
		19'b1100001110100110011: color_data = Z;
		19'b1100001110100110100: color_data = Z;
		19'b1100001110100110101: color_data = Z;
		19'b1100001110100110110: color_data = Z;
		19'b1100001110100110111: color_data = Z;
		19'b1100001110100111000: color_data = Z;
		19'b1100001110100111001: color_data = Z;
		19'b1100001110100111010: color_data = Z;
		19'b1100001110100111011: color_data = Z;
		19'b1100001110100111100: color_data = Z;
		19'b1100001110100111101: color_data = Z;
		19'b1100001110100111110: color_data = Z;
		19'b1100001110100111111: color_data = Z;
		19'b1100001110101000000: color_data = Z;
		19'b1100001110101000001: color_data = Z;
		19'b1100001110101000010: color_data = Z;
		19'b1100001110101000011: color_data = Z;
		19'b1100001110101000100: color_data = Z;
		19'b1100001110101000101: color_data = Z;
		19'b1100001110101000110: color_data = Z;
		19'b1100001110101000111: color_data = Z;
		19'b1100001110101001000: color_data = Z;
		19'b1100001110101001001: color_data = Z;
		19'b1100001110101001010: color_data = Z;
		19'b1100001110101001011: color_data = Z;
		19'b1100001110101001100: color_data = Z;
		19'b1100001110101001101: color_data = Z;
		19'b1100001110101001110: color_data = Z;
		19'b1100001110101001111: color_data = Z;
		19'b1100001110101010000: color_data = Z;
		19'b1100001110101011101: color_data = Z;
		19'b1100001110101011110: color_data = Z;
		19'b1100001110101011111: color_data = Z;
		19'b1100001110101100000: color_data = Z;
		19'b1100001110101100001: color_data = Z;
		19'b1100001110101100010: color_data = Z;
		19'b1100001110101100011: color_data = Z;
		19'b1100001110101100100: color_data = Z;
		19'b1100001110101100101: color_data = Z;
		19'b1100001110101100110: color_data = Z;
		19'b1100001110101100111: color_data = Z;
		19'b1100001110101101000: color_data = Z;
		19'b1100001110101101001: color_data = Z;
		19'b1100001110101101010: color_data = Z;
		19'b1100001110101101011: color_data = Z;
		19'b1100001110101101100: color_data = Z;
		19'b1100001110101101101: color_data = Z;
		19'b1100001110101101110: color_data = Z;
		19'b1100001110101101111: color_data = Z;
		19'b1100001110101110000: color_data = Z;
		19'b1100001110101110001: color_data = Z;
		19'b1100001110101110010: color_data = Z;
		19'b1100001110101110011: color_data = Z;
		19'b1100001110101110100: color_data = Z;
		19'b1100001110101110101: color_data = Z;
		19'b1100001110101110110: color_data = Z;
		19'b1100010000100100111: color_data = Z;
		19'b1100010000100101000: color_data = Z;
		19'b1100010000100101001: color_data = Z;
		19'b1100010000100101010: color_data = Z;
		19'b1100010000100101011: color_data = Z;
		19'b1100010000100101100: color_data = Z;
		19'b1100010000100101101: color_data = Z;
		19'b1100010000100101110: color_data = Z;
		19'b1100010000100101111: color_data = Z;
		19'b1100010000100110000: color_data = Z;
		19'b1100010000100110001: color_data = Z;
		19'b1100010000100110010: color_data = Z;
		19'b1100010000100110011: color_data = Z;
		19'b1100010000100110100: color_data = Z;
		19'b1100010000100110101: color_data = Z;
		19'b1100010000100110110: color_data = Z;
		19'b1100010000100110111: color_data = Z;
		19'b1100010000100111000: color_data = Z;
		19'b1100010000100111001: color_data = Z;
		19'b1100010000100111010: color_data = Z;
		19'b1100010000100111011: color_data = Z;
		19'b1100010000100111100: color_data = Z;
		19'b1100010000100111101: color_data = Z;
		19'b1100010000100111110: color_data = Z;
		19'b1100010000100111111: color_data = Z;
		19'b1100010000101000000: color_data = Z;
		19'b1100010000101000001: color_data = Z;
		19'b1100010000101000010: color_data = Z;
		19'b1100010000101000011: color_data = Z;
		19'b1100010000101000100: color_data = Z;
		19'b1100010000101000101: color_data = Z;
		19'b1100010000101000110: color_data = Z;
		19'b1100010000101000111: color_data = Z;
		19'b1100010000101001000: color_data = Z;
		19'b1100010000101001001: color_data = Z;
		19'b1100010000101001010: color_data = Z;
		19'b1100010000101001011: color_data = Z;
		19'b1100010000101001100: color_data = Z;
		19'b1100010000101001101: color_data = Z;
		19'b1100010000101001110: color_data = Z;
		19'b1100010000101001111: color_data = Z;
		19'b1100010000101010000: color_data = Z;
		19'b1100010000101010001: color_data = Z;
		19'b1100010000101010010: color_data = Z;
		19'b1100010000101010011: color_data = Z;
		19'b1100010000101010111: color_data = Z;
		19'b1100010000101011000: color_data = Z;
		19'b1100010000101011001: color_data = Z;
		19'b1100010000101011010: color_data = Z;
		19'b1100010000101011011: color_data = Z;
		19'b1100010000101011100: color_data = Z;
		19'b1100010000101011101: color_data = Z;
		19'b1100010000101011110: color_data = Z;
		19'b1100010000101011111: color_data = Z;
		19'b1100010000101100000: color_data = Z;
		19'b1100010000101100001: color_data = Z;
		19'b1100010000101100010: color_data = Z;
		19'b1100010000101100011: color_data = Z;
		19'b1100010000101100100: color_data = Z;
		19'b1100010000101100101: color_data = Z;
		19'b1100010000101100110: color_data = Z;
		19'b1100010000101100111: color_data = Z;
		19'b1100010000101101000: color_data = Z;
		19'b1100010000101101001: color_data = Z;
		19'b1100010000101101010: color_data = Z;
		19'b1100010000101101011: color_data = Z;
		19'b1100010000101101100: color_data = Z;
		19'b1100010000101101101: color_data = Z;
		19'b1100010000101101110: color_data = Z;
		19'b1100010000101101111: color_data = Z;
		19'b1100010000101110000: color_data = Z;
		19'b1100010000101110001: color_data = Z;
		19'b1100010000101110010: color_data = Z;
		19'b1100010000101110011: color_data = Z;
		19'b1100010000101110100: color_data = Z;
		19'b1100010010100101001: color_data = Z;
		19'b1100010010100101010: color_data = Z;
		19'b1100010010100101011: color_data = Z;
		19'b1100010010100101100: color_data = Z;
		19'b1100010010100101101: color_data = Z;
		19'b1100010010100101110: color_data = Z;
		19'b1100010010100101111: color_data = Z;
		19'b1100010010100110000: color_data = Z;
		19'b1100010010100110001: color_data = Z;
		19'b1100010010100110010: color_data = Z;
		19'b1100010010100110011: color_data = Z;
		19'b1100010010100110100: color_data = Z;
		19'b1100010010100110101: color_data = Z;
		19'b1100010010100110110: color_data = Z;
		19'b1100010010100110111: color_data = Z;
		19'b1100010010100111000: color_data = Z;
		19'b1100010010100111001: color_data = Z;
		19'b1100010010100111010: color_data = Z;
		19'b1100010010100111011: color_data = Z;
		19'b1100010010100111100: color_data = Z;
		19'b1100010010100111101: color_data = Z;
		19'b1100010010100111110: color_data = Z;
		19'b1100010010100111111: color_data = Z;
		19'b1100010010101000000: color_data = Z;
		19'b1100010010101000001: color_data = Z;
		19'b1100010010101000010: color_data = Z;
		19'b1100010010101000011: color_data = Z;
		19'b1100010010101000100: color_data = Z;
		19'b1100010010101000101: color_data = Z;
		19'b1100010010101000110: color_data = Z;
		19'b1100010010101000111: color_data = Z;
		19'b1100010010101001000: color_data = Z;
		19'b1100010010101001001: color_data = Z;
		19'b1100010010101001010: color_data = Z;
		19'b1100010010101001011: color_data = Z;
		19'b1100010010101001100: color_data = Z;
		19'b1100010010101001101: color_data = Z;
		19'b1100010010101001110: color_data = Z;
		19'b1100010010101001111: color_data = Z;
		19'b1100010010101010000: color_data = Z;
		19'b1100010010101010001: color_data = Z;
		19'b1100010010101010010: color_data = Z;
		19'b1100010010101010011: color_data = Z;
		19'b1100010010101010100: color_data = Z;
		19'b1100010010101010101: color_data = Z;
		19'b1100010010101010110: color_data = Z;
		19'b1100010010101010111: color_data = Z;
		19'b1100010010101011000: color_data = Z;
		19'b1100010010101011001: color_data = Z;
		19'b1100010010101011010: color_data = Z;
		19'b1100010010101011011: color_data = Z;
		19'b1100010010101011100: color_data = Z;
		19'b1100010010101011101: color_data = Z;
		19'b1100010010101011110: color_data = Z;
		19'b1100010010101011111: color_data = Z;
		19'b1100010010101100000: color_data = Z;
		19'b1100010010101100001: color_data = Z;
		19'b1100010010101100010: color_data = Z;
		19'b1100010010101100011: color_data = Z;
		19'b1100010010101100100: color_data = Z;
		19'b1100010010101100101: color_data = Z;
		19'b1100010010101100110: color_data = Z;
		19'b1100010010101100111: color_data = Z;
		19'b1100010010101101000: color_data = Z;
		19'b1100010010101101001: color_data = Z;
		19'b1100010010101101010: color_data = Z;
		19'b1100010010101101011: color_data = Z;
		19'b1100010010101101100: color_data = Z;
		19'b1100010010101101101: color_data = Z;
		19'b1100010010101101110: color_data = Z;
		19'b1100010010101101111: color_data = Z;
		19'b1100010010101110000: color_data = Z;
		19'b1100010010101110001: color_data = Z;
		19'b1100010010101110010: color_data = Z;
		19'b1100010100100101011: color_data = Z;
		19'b1100010100100101100: color_data = Z;
		19'b1100010100100101101: color_data = Z;
		19'b1100010100100101110: color_data = Z;
		19'b1100010100100101111: color_data = Z;
		19'b1100010100100110000: color_data = Z;
		19'b1100010100100110001: color_data = Z;
		19'b1100010100100110010: color_data = Z;
		19'b1100010100100110011: color_data = Z;
		19'b1100010100100110100: color_data = Z;
		19'b1100010100100110101: color_data = Z;
		19'b1100010100100110110: color_data = Z;
		19'b1100010100100110111: color_data = Z;
		19'b1100010100100111000: color_data = Z;
		19'b1100010100100111001: color_data = Z;
		19'b1100010100100111010: color_data = Z;
		19'b1100010100100111011: color_data = Z;
		19'b1100010100100111100: color_data = Z;
		19'b1100010100100111101: color_data = Z;
		19'b1100010100100111110: color_data = Z;
		19'b1100010100100111111: color_data = Z;
		19'b1100010100101000000: color_data = Z;
		19'b1100010100101000001: color_data = Z;
		19'b1100010100101000010: color_data = Z;
		19'b1100010100101000011: color_data = Z;
		19'b1100010100101000100: color_data = Z;
		19'b1100010100101000101: color_data = Z;
		19'b1100010100101000110: color_data = Z;
		19'b1100010100101000111: color_data = Z;
		19'b1100010100101001000: color_data = Z;
		19'b1100010100101001001: color_data = Z;
		19'b1100010100101001010: color_data = Z;
		19'b1100010100101001011: color_data = Z;
		19'b1100010100101001100: color_data = Z;
		19'b1100010100101001101: color_data = Z;
		19'b1100010100101001110: color_data = Z;
		19'b1100010100101001111: color_data = Z;
		19'b1100010100101010000: color_data = Z;
		19'b1100010100101010001: color_data = Z;
		19'b1100010100101010010: color_data = Z;
		19'b1100010100101010011: color_data = Z;
		19'b1100010100101010100: color_data = Z;
		19'b1100010100101010101: color_data = Z;
		19'b1100010100101010110: color_data = Z;
		19'b1100010100101010111: color_data = Z;
		19'b1100010100101011000: color_data = Z;
		19'b1100010100101011001: color_data = Z;
		19'b1100010100101011010: color_data = Z;
		19'b1100010100101011011: color_data = Z;
		19'b1100010100101011100: color_data = Z;
		19'b1100010100101011101: color_data = Z;
		19'b1100010100101011110: color_data = Z;
		19'b1100010100101011111: color_data = Z;
		19'b1100010100101100000: color_data = Z;
		19'b1100010100101100001: color_data = Z;
		19'b1100010100101100010: color_data = Z;
		19'b1100010100101100011: color_data = Z;
		19'b1100010100101100100: color_data = Z;
		19'b1100010100101100101: color_data = Z;
		19'b1100010100101100110: color_data = Z;
		19'b1100010100101100111: color_data = Z;
		19'b1100010100101101000: color_data = Z;
		19'b1100010100101101001: color_data = Z;
		19'b1100010100101101010: color_data = Z;
		19'b1100010100101101011: color_data = Z;
		19'b1100010100101101100: color_data = Z;
		19'b1100010100101101101: color_data = Z;
		19'b1100010100101101110: color_data = Z;
		19'b1100010100101101111: color_data = Z;
		19'b1100010100101110000: color_data = Z;
		19'b1100010100101110001: color_data = Z;
		19'b1100010110100101100: color_data = Z;
		19'b1100010110100101101: color_data = Z;
		19'b1100010110100101110: color_data = Z;
		19'b1100010110100101111: color_data = Z;
		19'b1100010110100110000: color_data = Z;
		19'b1100010110100110001: color_data = Z;
		19'b1100010110100110010: color_data = Z;
		19'b1100010110100110011: color_data = Z;
		19'b1100010110100110100: color_data = Z;
		19'b1100010110100110101: color_data = Z;
		19'b1100010110100110110: color_data = Z;
		19'b1100010110100110111: color_data = Z;
		19'b1100010110100111000: color_data = Z;
		19'b1100010110100111001: color_data = Z;
		19'b1100010110100111010: color_data = Z;
		19'b1100010110100111011: color_data = Z;
		19'b1100010110100111100: color_data = Z;
		19'b1100010110100111101: color_data = Z;
		19'b1100010110100111110: color_data = Z;
		19'b1100010110100111111: color_data = Z;
		19'b1100010110101000000: color_data = Z;
		19'b1100010110101000001: color_data = Z;
		19'b1100010110101000010: color_data = Z;
		19'b1100010110101000011: color_data = Z;
		19'b1100010110101000100: color_data = Z;
		19'b1100010110101000101: color_data = Z;
		19'b1100010110101000110: color_data = Z;
		19'b1100010110101000111: color_data = Z;
		19'b1100010110101001000: color_data = Z;
		19'b1100010110101001001: color_data = Z;
		19'b1100010110101001010: color_data = Z;
		19'b1100010110101001011: color_data = Z;
		19'b1100010110101001100: color_data = Z;
		19'b1100010110101001101: color_data = Z;
		19'b1100010110101001110: color_data = Z;
		19'b1100010110101001111: color_data = Z;
		19'b1100010110101010000: color_data = Z;
		19'b1100010110101010001: color_data = Z;
		19'b1100010110101010010: color_data = Z;
		19'b1100010110101010011: color_data = Z;
		19'b1100010110101010100: color_data = Z;
		19'b1100010110101010101: color_data = Z;
		19'b1100010110101010110: color_data = Z;
		19'b1100010110101010111: color_data = Z;
		19'b1100010110101011000: color_data = Z;
		19'b1100010110101011001: color_data = Z;
		19'b1100010110101011010: color_data = Z;
		19'b1100010110101011011: color_data = Z;
		19'b1100010110101011100: color_data = Z;
		19'b1100010110101011101: color_data = Z;
		19'b1100010110101011110: color_data = Z;
		19'b1100010110101011111: color_data = Z;
		19'b1100010110101100000: color_data = Z;
		19'b1100010110101100001: color_data = Z;
		19'b1100010110101100010: color_data = Z;
		19'b1100010110101100011: color_data = Z;
		19'b1100010110101100100: color_data = Z;
		19'b1100010110101100101: color_data = Z;
		19'b1100010110101100110: color_data = Z;
		19'b1100010110101100111: color_data = Z;
		19'b1100010110101101000: color_data = Z;
		19'b1100010110101101001: color_data = Z;
		19'b1100010110101101010: color_data = Z;
		19'b1100010110101101011: color_data = Z;
		19'b1100010110101101100: color_data = Z;
		19'b1100010110101101101: color_data = Z;
		19'b1100010110101101110: color_data = Z;
		19'b1100010110101101111: color_data = Z;
		19'b1100010110101110000: color_data = Z;
		19'b1100010110101110001: color_data = Z;
		19'b1100011000100101110: color_data = Z;
		19'b1100011000100101111: color_data = Z;
		19'b1100011000100110000: color_data = Z;
		19'b1100011000100110001: color_data = Z;
		19'b1100011000100110010: color_data = Z;
		19'b1100011000100110011: color_data = Z;
		19'b1100011000100110100: color_data = Z;
		19'b1100011000100110101: color_data = Z;
		19'b1100011000100110110: color_data = Z;
		19'b1100011000100110111: color_data = Z;
		19'b1100011000100111000: color_data = Z;
		19'b1100011000100111001: color_data = Z;
		19'b1100011000100111010: color_data = Z;
		19'b1100011000100111011: color_data = Z;
		19'b1100011000100111100: color_data = Z;
		19'b1100011000100111101: color_data = Z;
		19'b1100011000100111110: color_data = Z;
		19'b1100011000100111111: color_data = Z;
		19'b1100011000101000000: color_data = Z;
		19'b1100011000101000001: color_data = Z;
		19'b1100011000101000010: color_data = Z;
		19'b1100011000101000011: color_data = Z;
		19'b1100011000101000100: color_data = Z;
		19'b1100011000101000101: color_data = Z;
		19'b1100011000101000110: color_data = Z;
		19'b1100011000101000111: color_data = Z;
		19'b1100011000101001000: color_data = Z;
		19'b1100011000101001001: color_data = Z;
		19'b1100011000101001010: color_data = Z;
		19'b1100011000101001011: color_data = Z;
		19'b1100011000101001100: color_data = Z;
		19'b1100011000101001101: color_data = Z;
		19'b1100011000101001110: color_data = Z;
		19'b1100011000101001111: color_data = Z;
		19'b1100011000101010000: color_data = Z;
		19'b1100011000101010001: color_data = Z;
		19'b1100011000101010010: color_data = Z;
		19'b1100011000101010011: color_data = Z;
		19'b1100011000101010100: color_data = Z;
		19'b1100011000101010101: color_data = Z;
		19'b1100011000101010110: color_data = Z;
		19'b1100011000101010111: color_data = Z;
		19'b1100011000101011000: color_data = Z;
		19'b1100011000101011001: color_data = Z;
		19'b1100011000101011010: color_data = Z;
		19'b1100011000101011011: color_data = Z;
		19'b1100011000101011100: color_data = Z;
		19'b1100011000101011101: color_data = Z;
		19'b1100011000101011110: color_data = Z;
		19'b1100011000101011111: color_data = Z;
		19'b1100011000101100000: color_data = Z;
		19'b1100011000101100001: color_data = Z;
		19'b1100011000101100010: color_data = Z;
		19'b1100011000101100011: color_data = Z;
		19'b1100011000101100100: color_data = Z;
		19'b1100011000101100101: color_data = Z;
		19'b1100011000101100110: color_data = Z;
		19'b1100011000101100111: color_data = Z;
		19'b1100011000101101000: color_data = Z;
		19'b1100011000101101001: color_data = Z;
		19'b1100011000101101010: color_data = Z;
		19'b1100011000101101011: color_data = Z;
		19'b1100011000101101100: color_data = Z;
		19'b1100011000101101101: color_data = Z;
		19'b1100011000101101110: color_data = Z;
		19'b1100011000101101111: color_data = Z;
		19'b1100011000101110000: color_data = Z;
		19'b1100011010100110000: color_data = Z;
		19'b1100011010100110001: color_data = Z;
		19'b1100011010100110010: color_data = Z;
		19'b1100011010100110011: color_data = Z;
		19'b1100011010100110100: color_data = Z;
		19'b1100011010100110101: color_data = Z;
		19'b1100011010100110110: color_data = Z;
		19'b1100011010100110111: color_data = Z;
		19'b1100011010100111000: color_data = Z;
		19'b1100011010100111001: color_data = Z;
		19'b1100011010100111010: color_data = Z;
		19'b1100011010100111011: color_data = Z;
		19'b1100011010100111100: color_data = Z;
		19'b1100011010100111101: color_data = Z;
		19'b1100011010100111110: color_data = Z;
		19'b1100011010100111111: color_data = Z;
		19'b1100011010101000000: color_data = Z;
		19'b1100011010101000001: color_data = Z;
		19'b1100011010101000010: color_data = Z;
		19'b1100011010101000011: color_data = Z;
		19'b1100011010101000100: color_data = Z;
		19'b1100011010101000101: color_data = Z;
		19'b1100011010101000110: color_data = Z;
		19'b1100011010101000111: color_data = Z;
		19'b1100011010101001000: color_data = Z;
		19'b1100011010101001001: color_data = Z;
		19'b1100011010101001010: color_data = Z;
		19'b1100011010101001011: color_data = Z;
		19'b1100011010101001100: color_data = Z;
		19'b1100011010101001101: color_data = Z;
		19'b1100011010101001110: color_data = Z;
		19'b1100011010101001111: color_data = Z;
		19'b1100011010101010000: color_data = Z;
		19'b1100011010101010001: color_data = Z;
		19'b1100011010101010010: color_data = Z;
		19'b1100011010101010011: color_data = Z;
		19'b1100011010101010100: color_data = Z;
		19'b1100011010101010101: color_data = Z;
		19'b1100011010101010110: color_data = Z;
		19'b1100011010101010111: color_data = Z;
		19'b1100011010101011000: color_data = Z;
		19'b1100011010101011001: color_data = Z;
		19'b1100011010101011010: color_data = Z;
		19'b1100011010101011011: color_data = Z;
		19'b1100011010101011100: color_data = Z;
		19'b1100011010101011101: color_data = Z;
		19'b1100011010101011110: color_data = Z;
		19'b1100011010101011111: color_data = Z;
		19'b1100011010101100000: color_data = Z;
		19'b1100011010101100001: color_data = Z;
		19'b1100011010101100010: color_data = Z;
		19'b1100011010101100011: color_data = Z;
		19'b1100011010101100100: color_data = Z;
		19'b1100011010101100101: color_data = Z;
		19'b1100011010101100110: color_data = Z;
		19'b1100011010101100111: color_data = Z;
		19'b1100011010101101000: color_data = Z;
		19'b1100011010101101001: color_data = Z;
		19'b1100011010101101010: color_data = Z;
		19'b1100011010101101011: color_data = Z;
		19'b1100011010101101100: color_data = Z;
		19'b1100011010101101101: color_data = Z;
		19'b1100011010101101110: color_data = Z;
		19'b1100011010101101111: color_data = Z;
		19'b1100011100100110010: color_data = Z;
		19'b1100011100100110011: color_data = Z;
		19'b1100011100100110100: color_data = Z;
		19'b1100011100100110101: color_data = Z;
		19'b1100011100100110110: color_data = Z;
		19'b1100011100100110111: color_data = Z;
		19'b1100011100100111000: color_data = Z;
		19'b1100011100100111001: color_data = Z;
		19'b1100011100100111010: color_data = Z;
		19'b1100011100100111011: color_data = Z;
		19'b1100011100100111100: color_data = Z;
		19'b1100011100100111101: color_data = Z;
		19'b1100011100100111110: color_data = Z;
		19'b1100011100100111111: color_data = Z;
		19'b1100011100101000000: color_data = Z;
		19'b1100011100101000001: color_data = Z;
		19'b1100011100101000010: color_data = Z;
		19'b1100011100101000011: color_data = Z;
		19'b1100011100101000100: color_data = Z;
		19'b1100011100101000101: color_data = Z;
		19'b1100011100101000110: color_data = Z;
		19'b1100011100101000111: color_data = Z;
		19'b1100011100101001000: color_data = Z;
		19'b1100011100101001001: color_data = Z;
		19'b1100011100101001010: color_data = Z;
		19'b1100011100101001011: color_data = Z;
		19'b1100011100101001100: color_data = Z;
		19'b1100011100101001101: color_data = Z;
		19'b1100011100101001110: color_data = Z;
		19'b1100011100101001111: color_data = Z;
		19'b1100011100101010000: color_data = Z;
		19'b1100011100101010001: color_data = Z;
		19'b1100011100101010010: color_data = Z;
		19'b1100011100101010011: color_data = Z;
		19'b1100011100101010100: color_data = Z;
		19'b1100011100101010101: color_data = Z;
		19'b1100011100101010110: color_data = Z;
		19'b1100011100101010111: color_data = Z;
		19'b1100011100101011000: color_data = Z;
		19'b1100011100101011001: color_data = Z;
		19'b1100011100101011010: color_data = Z;
		19'b1100011100101011011: color_data = Z;
		19'b1100011100101011100: color_data = Z;
		19'b1100011100101011101: color_data = Z;
		19'b1100011100101011110: color_data = Z;
		19'b1100011100101011111: color_data = Z;
		19'b1100011100101100000: color_data = Z;
		19'b1100011100101100001: color_data = Z;
		19'b1100011100101100010: color_data = Z;
		19'b1100011100101100011: color_data = Z;
		19'b1100011100101100100: color_data = Z;
		19'b1100011100101100101: color_data = Z;
		19'b1100011100101100110: color_data = Z;
		19'b1100011100101100111: color_data = Z;
		19'b1100011100101101000: color_data = Z;
		19'b1100011100101101001: color_data = Z;
		19'b1100011100101101010: color_data = Z;
		19'b1100011100101101011: color_data = Z;
		19'b1100011100101101100: color_data = Z;
		19'b1100011100101101101: color_data = Z;
		19'b1100011100101101110: color_data = Z;
		19'b1100011110100110100: color_data = Z;
		19'b1100011110100110101: color_data = Z;
		19'b1100011110100110110: color_data = Z;
		19'b1100011110100110111: color_data = Z;
		19'b1100011110100111000: color_data = Z;
		19'b1100011110100111001: color_data = Z;
		19'b1100011110100111010: color_data = Z;
		19'b1100011110100111011: color_data = Z;
		19'b1100011110100111100: color_data = Z;
		19'b1100011110100111101: color_data = Z;
		19'b1100011110100111110: color_data = Z;
		19'b1100011110100111111: color_data = Z;
		19'b1100011110101000000: color_data = Z;
		19'b1100011110101000001: color_data = Z;
		19'b1100011110101000010: color_data = Z;
		19'b1100011110101000011: color_data = Z;
		19'b1100011110101000100: color_data = Z;
		19'b1100011110101000101: color_data = Z;
		19'b1100011110101000110: color_data = Z;
		19'b1100011110101000111: color_data = Z;
		19'b1100011110101001000: color_data = Z;
		19'b1100011110101001001: color_data = Z;
		19'b1100011110101001010: color_data = Z;
		19'b1100011110101001011: color_data = Z;
		19'b1100011110101001100: color_data = Z;
		19'b1100011110101001101: color_data = Z;
		19'b1100011110101001110: color_data = Z;
		19'b1100011110101001111: color_data = Z;
		19'b1100011110101010000: color_data = Z;
		19'b1100011110101010001: color_data = Z;
		19'b1100011110101010010: color_data = Z;
		19'b1100011110101010011: color_data = Z;
		19'b1100011110101010100: color_data = Z;
		19'b1100011110101010101: color_data = Z;
		19'b1100011110101010110: color_data = Z;
		19'b1100011110101010111: color_data = Z;
		19'b1100011110101011000: color_data = Z;
		19'b1100011110101011001: color_data = Z;
		19'b1100011110101011010: color_data = Z;
		19'b1100011110101011011: color_data = Z;
		19'b1100011110101011100: color_data = Z;
		19'b1100011110101011101: color_data = Z;
		19'b1100011110101011110: color_data = Z;
		19'b1100011110101011111: color_data = Z;
		19'b1100011110101100000: color_data = Z;
		19'b1100011110101100001: color_data = Z;
		19'b1100011110101100010: color_data = Z;
		19'b1100011110101100011: color_data = Z;
		19'b1100011110101100100: color_data = Z;
		19'b1100011110101100101: color_data = Z;
		19'b1100011110101100110: color_data = Z;
		19'b1100011110101100111: color_data = Z;
		19'b1100011110101101000: color_data = Z;
		19'b1100011110101101001: color_data = Z;
		19'b1100011110101101010: color_data = Z;
		19'b1100011110101101011: color_data = Z;
		19'b1100011110101101100: color_data = Z;
		19'b1100011110101101101: color_data = Z;
		19'b1100100000100110110: color_data = Z;
		19'b1100100000100110111: color_data = Z;
		19'b1100100000100111000: color_data = Z;
		19'b1100100000100111001: color_data = Z;
		19'b1100100000100111010: color_data = Z;
		19'b1100100000100111011: color_data = Z;
		19'b1100100000100111100: color_data = Z;
		19'b1100100000100111101: color_data = Z;
		19'b1100100000100111110: color_data = Z;
		19'b1100100000100111111: color_data = Z;
		19'b1100100000101000000: color_data = Z;
		19'b1100100000101000001: color_data = Z;
		19'b1100100000101000010: color_data = Z;
		19'b1100100000101000011: color_data = Z;
		19'b1100100000101000100: color_data = Z;
		19'b1100100000101000101: color_data = Z;
		19'b1100100000101000110: color_data = Z;
		19'b1100100000101000111: color_data = Z;
		19'b1100100000101001000: color_data = Z;
		19'b1100100000101001001: color_data = Z;
		19'b1100100000101001010: color_data = Z;
		19'b1100100000101001011: color_data = Z;
		19'b1100100000101001100: color_data = Z;
		19'b1100100000101001101: color_data = Z;
		19'b1100100000101001110: color_data = Z;
		19'b1100100000101001111: color_data = Z;
		19'b1100100000101010000: color_data = Z;
		19'b1100100000101010001: color_data = Z;
		19'b1100100000101010010: color_data = Z;
		19'b1100100000101010011: color_data = Z;
		19'b1100100000101010100: color_data = Z;
		19'b1100100000101010101: color_data = Z;
		19'b1100100000101010110: color_data = Z;
		19'b1100100000101010111: color_data = Z;
		19'b1100100000101011000: color_data = Z;
		19'b1100100000101011001: color_data = Z;
		19'b1100100000101011010: color_data = Z;
		19'b1100100000101011011: color_data = Z;
		19'b1100100000101011100: color_data = Z;
		19'b1100100000101011101: color_data = Z;
		19'b1100100000101011110: color_data = Z;
		19'b1100100000101011111: color_data = Z;
		19'b1100100000101100000: color_data = Z;
		19'b1100100000101100001: color_data = Z;
		19'b1100100000101100010: color_data = Z;
		19'b1100100000101100011: color_data = Z;
		19'b1100100000101100100: color_data = Z;
		19'b1100100000101100101: color_data = Z;
		19'b1100100000101100110: color_data = Z;
		19'b1100100000101100111: color_data = Z;
		19'b1100100000101101000: color_data = Z;
		19'b1100100000101101001: color_data = Z;
		19'b1100100000101101010: color_data = Z;
		19'b1100100000101101011: color_data = Z;
		19'b1100100010100111000: color_data = Z;
		19'b1100100010100111001: color_data = Z;
		19'b1100100010100111010: color_data = Z;
		19'b1100100010100111011: color_data = Z;
		19'b1100100010100111100: color_data = Z;
		19'b1100100010100111101: color_data = Z;
		19'b1100100010100111110: color_data = Z;
		19'b1100100010100111111: color_data = Z;
		19'b1100100010101000000: color_data = Z;
		19'b1100100010101000001: color_data = Z;
		19'b1100100010101000010: color_data = Z;
		19'b1100100010101000011: color_data = Z;
		19'b1100100010101000100: color_data = Z;
		19'b1100100010101000101: color_data = Z;
		19'b1100100010101000110: color_data = Z;
		19'b1100100010101000111: color_data = Z;
		19'b1100100010101001000: color_data = Z;
		19'b1100100010101001001: color_data = Z;
		19'b1100100010101001010: color_data = Z;
		19'b1100100010101001011: color_data = Z;
		19'b1100100010101001100: color_data = Z;
		19'b1100100010101001101: color_data = Z;
		19'b1100100010101001110: color_data = Z;
		19'b1100100010101001111: color_data = Z;
		19'b1100100010101010000: color_data = Z;
		19'b1100100010101010001: color_data = Z;
		19'b1100100010101010010: color_data = Z;
		19'b1100100010101010011: color_data = Z;
		19'b1100100010101010100: color_data = Z;
		19'b1100100010101010101: color_data = Z;
		19'b1100100010101010110: color_data = Z;
		19'b1100100010101010111: color_data = Z;
		19'b1100100010101011000: color_data = Z;
		19'b1100100010101011001: color_data = Z;
		19'b1100100010101011010: color_data = Z;
		19'b1100100010101011011: color_data = Z;
		19'b1100100010101011100: color_data = Z;
		19'b1100100010101011101: color_data = Z;
		19'b1100100010101011110: color_data = Z;
		19'b1100100010101011111: color_data = Z;
		19'b1100100010101100000: color_data = Z;
		19'b1100100010101100001: color_data = Z;
		19'b1100100010101100010: color_data = Z;
		19'b1100100010101100011: color_data = Z;
		19'b1100100010101100100: color_data = Z;
		19'b1100100010101100101: color_data = Z;
		19'b1100100010101100110: color_data = Z;
		19'b1100100010101100111: color_data = Z;
		19'b1100100010101101000: color_data = Z;
		19'b1100100010101101001: color_data = Z;
		19'b1100100010101101010: color_data = Z;
		19'b1100100100100111011: color_data = Z;
		19'b1100100100100111100: color_data = Z;
		19'b1100100100100111101: color_data = Z;
		19'b1100100100100111110: color_data = Z;
		19'b1100100100100111111: color_data = Z;
		19'b1100100100101000000: color_data = Z;
		19'b1100100100101000001: color_data = Z;
		19'b1100100100101000010: color_data = Z;
		19'b1100100100101000011: color_data = Z;
		19'b1100100100101000100: color_data = Z;
		19'b1100100100101000101: color_data = Z;
		19'b1100100100101000110: color_data = Z;
		19'b1100100100101000111: color_data = Z;
		19'b1100100100101001000: color_data = Z;
		19'b1100100100101001001: color_data = Z;
		19'b1100100100101001010: color_data = Z;
		19'b1100100100101001011: color_data = Z;
		19'b1100100100101001100: color_data = Z;
		19'b1100100100101001101: color_data = Z;
		19'b1100100100101001110: color_data = Z;
		19'b1100100100101001111: color_data = Z;
		19'b1100100100101010000: color_data = Z;
		19'b1100100100101010001: color_data = Z;
		19'b1100100100101010010: color_data = Z;
		19'b1100100100101010011: color_data = Z;
		19'b1100100100101010100: color_data = Z;
		19'b1100100100101010101: color_data = Z;
		19'b1100100100101010110: color_data = Z;
		19'b1100100100101010111: color_data = Z;
		19'b1100100100101011000: color_data = Z;
		19'b1100100100101011001: color_data = Z;
		19'b1100100100101011010: color_data = Z;
		19'b1100100100101011011: color_data = Z;
		19'b1100100100101011100: color_data = Z;
		19'b1100100100101011101: color_data = Z;
		19'b1100100100101011110: color_data = Z;
		19'b1100100100101011111: color_data = Z;
		19'b1100100100101100000: color_data = Z;
		19'b1100100100101100001: color_data = Z;
		19'b1100100100101100010: color_data = Z;
		19'b1100100100101100011: color_data = Z;
		19'b1100100100101100100: color_data = Z;
		19'b1100100100101100101: color_data = Z;
		19'b1100100100101100110: color_data = Z;
		19'b1100100100101100111: color_data = Z;
		19'b1100100100101101000: color_data = Z;
		19'b1100100100101101001: color_data = Z;
		19'b1100100110100111101: color_data = Z;
		19'b1100100110100111110: color_data = Z;
		19'b1100100110100111111: color_data = Z;
		19'b1100100110101000000: color_data = Z;
		19'b1100100110101000001: color_data = Z;
		19'b1100100110101000010: color_data = Z;
		19'b1100100110101000011: color_data = Z;
		19'b1100100110101000100: color_data = Z;
		19'b1100100110101000101: color_data = Z;
		19'b1100100110101000110: color_data = Z;
		19'b1100100110101000111: color_data = Z;
		19'b1100100110101001000: color_data = Z;
		19'b1100100110101001001: color_data = Z;
		19'b1100100110101001010: color_data = Z;
		19'b1100100110101001011: color_data = Z;
		19'b1100100110101001100: color_data = Z;
		19'b1100100110101001101: color_data = Z;
		19'b1100100110101001110: color_data = Z;
		19'b1100100110101001111: color_data = Z;
		19'b1100100110101010000: color_data = Z;
		19'b1100100110101010001: color_data = Z;
		19'b1100100110101010010: color_data = Z;
		19'b1100100110101010011: color_data = Z;
		19'b1100100110101010100: color_data = Z;
		19'b1100100110101010101: color_data = Z;
		19'b1100100110101010110: color_data = Z;
		19'b1100100110101010111: color_data = Z;
		19'b1100100110101011000: color_data = Z;
		19'b1100100110101011001: color_data = Z;
		19'b1100100110101011010: color_data = Z;
		19'b1100100110101011011: color_data = Z;
		19'b1100100110101011100: color_data = Z;
		19'b1100100110101011101: color_data = Z;
		19'b1100100110101011110: color_data = Z;
		19'b1100100110101011111: color_data = Z;
		19'b1100100110101100000: color_data = Z;
		19'b1100100110101100001: color_data = Z;
		19'b1100100110101100010: color_data = Z;
		19'b1100100110101100011: color_data = Z;
		19'b1100100110101100100: color_data = Z;
		19'b1100100110101100101: color_data = Z;
		19'b1100100110101100110: color_data = Z;
		19'b1100100110101100111: color_data = Z;
		19'b1100100110101101000: color_data = Z;
		19'b1100101000100111111: color_data = Z;
		19'b1100101000101000000: color_data = Z;
		19'b1100101000101000001: color_data = Z;
		19'b1100101000101000010: color_data = Z;
		19'b1100101000101000011: color_data = Z;
		19'b1100101000101000100: color_data = Z;
		19'b1100101000101000101: color_data = Z;
		19'b1100101000101000110: color_data = Z;
		19'b1100101000101000111: color_data = Z;
		19'b1100101000101001000: color_data = Z;
		19'b1100101000101001001: color_data = Z;
		19'b1100101000101001010: color_data = Z;
		19'b1100101000101001011: color_data = Z;
		19'b1100101000101001100: color_data = Z;
		19'b1100101000101001101: color_data = Z;
		19'b1100101000101001110: color_data = Z;
		19'b1100101000101001111: color_data = Z;
		19'b1100101000101010000: color_data = Z;
		19'b1100101000101010001: color_data = Z;
		19'b1100101000101010010: color_data = Z;
		19'b1100101000101010011: color_data = Z;
		19'b1100101000101010100: color_data = Z;
		19'b1100101000101010101: color_data = Z;
		19'b1100101000101010110: color_data = Z;
		19'b1100101000101010111: color_data = Z;
		19'b1100101000101011000: color_data = Z;
		19'b1100101000101011001: color_data = Z;
		19'b1100101000101011010: color_data = Z;
		19'b1100101000101011011: color_data = Z;
		19'b1100101000101011100: color_data = Z;
		19'b1100101000101011101: color_data = Z;
		19'b1100101000101011110: color_data = Z;
		19'b1100101000101011111: color_data = Z;
		19'b1100101000101100000: color_data = Z;
		19'b1100101000101100001: color_data = Z;
		19'b1100101000101100010: color_data = Z;
		19'b1100101000101100011: color_data = Z;
		19'b1100101000101100100: color_data = Z;
		19'b1100101000101100101: color_data = Z;
		19'b1100101000101100110: color_data = Z;
		19'b1100101000101100111: color_data = Z;
		19'b1100101010101000001: color_data = Z;
		19'b1100101010101000010: color_data = Z;
		19'b1100101010101000011: color_data = Z;
		19'b1100101010101000100: color_data = Z;
		19'b1100101010101000101: color_data = Z;
		19'b1100101010101000110: color_data = Z;
		19'b1100101010101000111: color_data = Z;
		19'b1100101010101001000: color_data = Z;
		19'b1100101010101001001: color_data = Z;
		19'b1100101010101001010: color_data = Z;
		19'b1100101010101001011: color_data = Z;
		19'b1100101010101001100: color_data = Z;
		19'b1100101010101001101: color_data = Z;
		19'b1100101010101001110: color_data = Z;
		19'b1100101010101001111: color_data = Z;
		19'b1100101010101010000: color_data = Z;
		19'b1100101010101010001: color_data = Z;
		19'b1100101010101010010: color_data = Z;
		19'b1100101010101010011: color_data = Z;
		19'b1100101010101010100: color_data = Z;
		19'b1100101010101010101: color_data = Z;
		19'b1100101010101010110: color_data = Z;
		19'b1100101010101010111: color_data = Z;
		19'b1100101010101011000: color_data = Z;
		19'b1100101010101011001: color_data = Z;
		19'b1100101010101011010: color_data = Z;
		19'b1100101010101011011: color_data = Z;
		19'b1100101010101011100: color_data = Z;
		19'b1100101010101011101: color_data = Z;
		19'b1100101010101011110: color_data = Z;
		19'b1100101010101011111: color_data = Z;
		19'b1100101010101100000: color_data = Z;
		19'b1100101010101100001: color_data = Z;
		19'b1100101010101100010: color_data = Z;
		19'b1100101010101100011: color_data = Z;
		19'b1100101010101100100: color_data = Z;
		19'b1100101010101100101: color_data = Z;
		19'b1100101010101100110: color_data = Z;
		19'b1100101100101000010: color_data = Z;
		19'b1100101100101000011: color_data = Z;
		19'b1100101100101000100: color_data = Z;
		19'b1100101100101000101: color_data = Z;
		19'b1100101100101000110: color_data = Z;
		19'b1100101100101000111: color_data = Z;
		19'b1100101100101001000: color_data = Z;
		19'b1100101100101001001: color_data = Z;
		19'b1100101100101001010: color_data = Z;
		19'b1100101100101001011: color_data = Z;
		19'b1100101100101001100: color_data = Z;
		19'b1100101100101001101: color_data = Z;
		19'b1100101100101001110: color_data = Z;
		19'b1100101100101001111: color_data = Z;
		19'b1100101100101010000: color_data = Z;
		19'b1100101100101010001: color_data = Z;
		19'b1100101100101010010: color_data = Z;
		19'b1100101100101010011: color_data = Z;
		19'b1100101100101010100: color_data = Z;
		19'b1100101100101010101: color_data = Z;
		19'b1100101100101010110: color_data = Z;
		19'b1100101100101010111: color_data = Z;
		19'b1100101100101011000: color_data = Z;
		19'b1100101100101011001: color_data = Z;
		19'b1100101100101011010: color_data = Z;
		19'b1100101100101011011: color_data = Z;
		19'b1100101100101011100: color_data = Z;
		19'b1100101100101011101: color_data = Z;
		19'b1100101100101011110: color_data = Z;
		19'b1100101100101011111: color_data = Z;
		19'b1100101100101100000: color_data = Z;
		19'b1100101100101100001: color_data = Z;
		19'b1100101100101100010: color_data = Z;
		19'b1100101100101100011: color_data = Z;
		19'b1100101100101100100: color_data = Z;
		19'b1100101100101100101: color_data = Z;
		19'b1100101110101000100: color_data = Z;
		19'b1100101110101000101: color_data = Z;
		19'b1100101110101000110: color_data = Z;
		19'b1100101110101000111: color_data = Z;
		19'b1100101110101001000: color_data = Z;
		19'b1100101110101001001: color_data = Z;
		19'b1100101110101001010: color_data = Z;
		19'b1100101110101001011: color_data = Z;
		19'b1100101110101001100: color_data = Z;
		19'b1100101110101001101: color_data = Z;
		19'b1100101110101001110: color_data = Z;
		19'b1100101110101001111: color_data = Z;
		19'b1100101110101010000: color_data = Z;
		19'b1100101110101010001: color_data = Z;
		19'b1100101110101010010: color_data = Z;
		19'b1100101110101010011: color_data = Z;
		19'b1100101110101010100: color_data = Z;
		19'b1100101110101010101: color_data = Z;
		19'b1100101110101010110: color_data = Z;
		19'b1100101110101010111: color_data = Z;
		19'b1100101110101011000: color_data = Z;
		19'b1100101110101011001: color_data = Z;
		19'b1100101110101011010: color_data = Z;
		19'b1100101110101011011: color_data = Z;
		19'b1100101110101011100: color_data = Z;
		19'b1100101110101011101: color_data = Z;
		19'b1100101110101011110: color_data = Z;
		19'b1100101110101011111: color_data = Z;
		19'b1100101110101100000: color_data = Z;
		19'b1100101110101100001: color_data = Z;
		19'b1100101110101100010: color_data = Z;
		19'b1100101110101100011: color_data = Z;
		19'b1100110000101000110: color_data = Z;
		19'b1100110000101000111: color_data = Z;
		19'b1100110000101001000: color_data = Z;
		19'b1100110000101001001: color_data = Z;
		19'b1100110000101001010: color_data = Z;
		19'b1100110000101001011: color_data = Z;
		19'b1100110000101001100: color_data = Z;
		19'b1100110000101001101: color_data = Z;
		19'b1100110000101001110: color_data = Z;
		19'b1100110000101001111: color_data = Z;
		19'b1100110000101010000: color_data = Z;
		19'b1100110000101010001: color_data = Z;
		19'b1100110000101010010: color_data = Z;
		19'b1100110000101010011: color_data = Z;
		19'b1100110000101010100: color_data = Z;
		19'b1100110000101010101: color_data = Z;
		19'b1100110000101010110: color_data = Z;
		19'b1100110000101010111: color_data = Z;
		19'b1100110000101011000: color_data = Z;
		19'b1100110000101011001: color_data = Z;
		19'b1100110000101011010: color_data = Z;
		19'b1100110000101011011: color_data = Z;
		19'b1100110000101011100: color_data = Z;
		19'b1100110000101011101: color_data = Z;
		19'b1100110000101011110: color_data = Z;
		19'b1100110000101011111: color_data = Z;
		19'b1100110000101100000: color_data = Z;
		19'b1100110000101100001: color_data = Z;
		19'b1100110010101001001: color_data = Z;
		19'b1100110010101001010: color_data = Z;
		19'b1100110010101001011: color_data = Z;
		19'b1100110010101001100: color_data = Z;
		19'b1100110010101001101: color_data = Z;
		19'b1100110010101001110: color_data = Z;
		19'b1100110010101001111: color_data = Z;
		19'b1100110010101010000: color_data = Z;
		19'b1100110010101010001: color_data = Z;
		19'b1100110010101010010: color_data = Z;
		19'b1100110010101010011: color_data = Z;
		19'b1100110010101010100: color_data = Z;
		19'b1100110010101010101: color_data = Z;
		19'b1100110010101010110: color_data = Z;
		19'b1101001000100101000: color_data = Z;
		19'b1101001000100101001: color_data = Z;
		19'b1101001010100101000: color_data = Z;
		19'b1101001010100101001: color_data = Z;
		19'b1101001010100101010: color_data = Z;
		19'b1101001010100101011: color_data = Z;
		19'b1101001100100100111: color_data = Z;
		19'b1101001100100101000: color_data = Z;
		19'b1101001100100101001: color_data = Z;
		19'b1101001100100101010: color_data = Z;
		19'b1101001100100101011: color_data = Z;
		19'b1101001100100101100: color_data = Z;
		19'b1101001100100101101: color_data = Z;
		19'b1101001100100101110: color_data = Z;
		19'b1101001110100100111: color_data = Z;
		19'b1101001110100101000: color_data = Z;
		19'b1101001110100101001: color_data = Z;
		19'b1101001110100101010: color_data = Z;
		19'b1101001110100101011: color_data = Z;
		19'b1101001110100101100: color_data = Z;
		19'b1101001110100101101: color_data = Z;
		19'b1101001110100101110: color_data = Z;
		19'b1101001110100101111: color_data = Z;
		19'b1101001110100110000: color_data = Z;
		19'b1101010000100100111: color_data = Z;
		19'b1101010000100101000: color_data = Z;
		19'b1101010000100101001: color_data = Z;
		19'b1101010000100101010: color_data = Z;
		19'b1101010000100101011: color_data = Z;
		19'b1101010000100101100: color_data = Z;
		19'b1101010000100101101: color_data = Z;
		19'b1101010000100101110: color_data = Z;
		19'b1101010000100101111: color_data = Z;
		19'b1101010000100110000: color_data = Z;
		19'b1101010000100110001: color_data = Z;
		19'b1101010000100110010: color_data = Z;
		19'b1101010000101101001: color_data = Z;
		19'b1101010000101101010: color_data = Z;
		19'b1101010000101101011: color_data = Z;
		19'b1101010000101101100: color_data = Z;
		19'b1101010000101101101: color_data = Z;
		19'b1101010000101101110: color_data = Z;
		19'b1101010010100100111: color_data = Z;
		19'b1101010010100101000: color_data = Z;
		19'b1101010010100101001: color_data = Z;
		19'b1101010010100101010: color_data = Z;
		19'b1101010010100101011: color_data = Z;
		19'b1101010010100101100: color_data = Z;
		19'b1101010010100101101: color_data = Z;
		19'b1101010010100101110: color_data = Z;
		19'b1101010010100101111: color_data = Z;
		19'b1101010010100110000: color_data = Z;
		19'b1101010010100110001: color_data = Z;
		19'b1101010010100110010: color_data = Z;
		19'b1101010010100110011: color_data = Z;
		19'b1101010010100110100: color_data = Z;
		19'b1101010010100110101: color_data = Z;
		19'b1101010010101100110: color_data = Z;
		19'b1101010010101100111: color_data = Z;
		19'b1101010010101101000: color_data = Z;
		19'b1101010010101101001: color_data = Z;
		19'b1101010010101101010: color_data = Z;
		19'b1101010010101101011: color_data = Z;
		19'b1101010010101101100: color_data = Z;
		19'b1101010010101101101: color_data = Z;
		19'b1101010010101101110: color_data = Z;
		19'b1101010100100100111: color_data = Z;
		19'b1101010100100101000: color_data = Z;
		19'b1101010100100101001: color_data = Z;
		19'b1101010100100101010: color_data = Z;
		19'b1101010100100101011: color_data = Z;
		19'b1101010100100101100: color_data = Z;
		19'b1101010100100101101: color_data = Z;
		19'b1101010100100101110: color_data = Z;
		19'b1101010100100101111: color_data = Z;
		19'b1101010100100110000: color_data = Z;
		19'b1101010100100110001: color_data = Z;
		19'b1101010100100110010: color_data = Z;
		19'b1101010100100110011: color_data = Z;
		19'b1101010100100110100: color_data = Z;
		19'b1101010100100110101: color_data = Z;
		19'b1101010100100110110: color_data = Z;
		19'b1101010100100110111: color_data = Z;
		19'b1101010100101100011: color_data = Z;
		19'b1101010100101100100: color_data = Z;
		19'b1101010100101100101: color_data = Z;
		19'b1101010100101100110: color_data = Z;
		19'b1101010100101100111: color_data = Z;
		19'b1101010100101101000: color_data = Z;
		19'b1101010100101101001: color_data = Z;
		19'b1101010100101101010: color_data = Z;
		19'b1101010100101101011: color_data = Z;
		19'b1101010100101101100: color_data = Z;
		19'b1101010100101101101: color_data = Z;
		19'b1101010100101101110: color_data = Z;
		19'b1101010110100100111: color_data = Z;
		19'b1101010110100101000: color_data = Z;
		19'b1101010110100101001: color_data = Z;
		19'b1101010110100101010: color_data = Z;
		19'b1101010110100101011: color_data = Z;
		19'b1101010110100101100: color_data = Z;
		19'b1101010110100101101: color_data = Z;
		19'b1101010110100101110: color_data = Z;
		19'b1101010110100101111: color_data = Z;
		19'b1101010110100110000: color_data = Z;
		19'b1101010110100110001: color_data = Z;
		19'b1101010110100110010: color_data = Z;
		19'b1101010110100110011: color_data = Z;
		19'b1101010110100110100: color_data = Z;
		19'b1101010110100110101: color_data = Z;
		19'b1101010110100110110: color_data = Z;
		19'b1101010110100110111: color_data = Z;
		19'b1101010110101100001: color_data = Z;
		19'b1101010110101100010: color_data = Z;
		19'b1101010110101100011: color_data = Z;
		19'b1101010110101100100: color_data = Z;
		19'b1101010110101100101: color_data = Z;
		19'b1101010110101100110: color_data = Z;
		19'b1101010110101100111: color_data = Z;
		19'b1101010110101101000: color_data = Z;
		19'b1101010110101101001: color_data = Z;
		19'b1101010110101101010: color_data = Z;
		19'b1101010110101101011: color_data = Z;
		19'b1101010110101101100: color_data = Z;
		19'b1101010110101101101: color_data = Z;
		19'b1101010110101101110: color_data = Z;
		19'b1101011000100100111: color_data = Z;
		19'b1101011000100101000: color_data = Z;
		19'b1101011000100101001: color_data = Z;
		19'b1101011000100101010: color_data = Z;
		19'b1101011000100101011: color_data = Z;
		19'b1101011000100101100: color_data = Z;
		19'b1101011000100101101: color_data = Z;
		19'b1101011000100101110: color_data = Z;
		19'b1101011000100101111: color_data = Z;
		19'b1101011000100110000: color_data = Z;
		19'b1101011000100110001: color_data = Z;
		19'b1101011000100110010: color_data = Z;
		19'b1101011000100110011: color_data = Z;
		19'b1101011000100110100: color_data = Z;
		19'b1101011000100110101: color_data = Z;
		19'b1101011000100110110: color_data = Z;
		19'b1101011000100110111: color_data = Z;
		19'b1101011000100111000: color_data = Z;
		19'b1101011000100111001: color_data = Z;
		19'b1101011000101011101: color_data = Z;
		19'b1101011000101011110: color_data = Z;
		19'b1101011000101011111: color_data = Z;
		19'b1101011000101100000: color_data = Z;
		19'b1101011000101100001: color_data = Z;
		19'b1101011000101100010: color_data = Z;
		19'b1101011000101100011: color_data = Z;
		19'b1101011000101100100: color_data = Z;
		19'b1101011000101100101: color_data = Z;
		19'b1101011000101100110: color_data = Z;
		19'b1101011000101100111: color_data = Z;
		19'b1101011000101101000: color_data = Z;
		19'b1101011000101101001: color_data = Z;
		19'b1101011000101101010: color_data = Z;
		19'b1101011000101101011: color_data = Z;
		19'b1101011000101101100: color_data = Z;
		19'b1101011000101101101: color_data = Z;
		19'b1101011000101101110: color_data = Z;
		19'b1101011000101111001: color_data = Z;
		19'b1101011010100100111: color_data = Z;
		19'b1101011010100101000: color_data = Z;
		19'b1101011010100101001: color_data = Z;
		19'b1101011010100101010: color_data = Z;
		19'b1101011010100101011: color_data = Z;
		19'b1101011010100101100: color_data = Z;
		19'b1101011010100101101: color_data = Z;
		19'b1101011010100101110: color_data = Z;
		19'b1101011010100101111: color_data = Z;
		19'b1101011010100110000: color_data = Z;
		19'b1101011010100110001: color_data = Z;
		19'b1101011010100110010: color_data = Z;
		19'b1101011010100110011: color_data = Z;
		19'b1101011010100110100: color_data = Z;
		19'b1101011010100110101: color_data = Z;
		19'b1101011010100110110: color_data = Z;
		19'b1101011010100110111: color_data = Z;
		19'b1101011010100111000: color_data = Z;
		19'b1101011010100111001: color_data = Z;
		19'b1101011010100111010: color_data = Z;
		19'b1101011010101011001: color_data = Z;
		19'b1101011010101011010: color_data = Z;
		19'b1101011010101011011: color_data = Z;
		19'b1101011010101011100: color_data = Z;
		19'b1101011010101011101: color_data = Z;
		19'b1101011010101011110: color_data = Z;
		19'b1101011010101011111: color_data = Z;
		19'b1101011010101100000: color_data = Z;
		19'b1101011010101100001: color_data = Z;
		19'b1101011010101100010: color_data = Z;
		19'b1101011010101100011: color_data = Z;
		19'b1101011010101100100: color_data = Z;
		19'b1101011010101100101: color_data = Z;
		19'b1101011010101100110: color_data = Z;
		19'b1101011010101100111: color_data = Z;
		19'b1101011010101101000: color_data = Z;
		19'b1101011010101101001: color_data = Z;
		19'b1101011010101101010: color_data = Z;
		19'b1101011010101101011: color_data = Z;
		19'b1101011010101101100: color_data = Z;
		19'b1101011010101101101: color_data = Z;
		19'b1101011010101101110: color_data = Z;
		19'b1101011100100100111: color_data = Z;
		19'b1101011100100101000: color_data = Z;
		19'b1101011100100101001: color_data = Z;
		19'b1101011100100101010: color_data = Z;
		19'b1101011100100101011: color_data = Z;
		19'b1101011100100101100: color_data = Z;
		19'b1101011100100101101: color_data = Z;
		19'b1101011100100101110: color_data = Z;
		19'b1101011100100101111: color_data = Z;
		19'b1101011100100110000: color_data = Z;
		19'b1101011100100110001: color_data = Z;
		19'b1101011100100110010: color_data = Z;
		19'b1101011100100110011: color_data = Z;
		19'b1101011100100110100: color_data = Z;
		19'b1101011100100110101: color_data = Z;
		19'b1101011100100110110: color_data = Z;
		19'b1101011100100110111: color_data = Z;
		19'b1101011100100111000: color_data = Z;
		19'b1101011100100111001: color_data = Z;
		19'b1101011100100111010: color_data = Z;
		19'b1101011100100111011: color_data = Z;
		19'b1101011100101001011: color_data = Z;
		19'b1101011100101010110: color_data = Z;
		19'b1101011100101010111: color_data = Z;
		19'b1101011100101011000: color_data = Z;
		19'b1101011100101011001: color_data = Z;
		19'b1101011100101011010: color_data = Z;
		19'b1101011100101011011: color_data = Z;
		19'b1101011100101011100: color_data = Z;
		19'b1101011100101011101: color_data = Z;
		19'b1101011100101011110: color_data = Z;
		19'b1101011100101011111: color_data = Z;
		19'b1101011100101100000: color_data = Z;
		19'b1101011100101100001: color_data = Z;
		19'b1101011100101100010: color_data = Z;
		19'b1101011100101100011: color_data = Z;
		19'b1101011100101100100: color_data = Z;
		19'b1101011100101100101: color_data = Z;
		19'b1101011100101100110: color_data = Z;
		19'b1101011100101100111: color_data = Z;
		19'b1101011100101101000: color_data = Z;
		19'b1101011100101101001: color_data = Z;
		19'b1101011100101101010: color_data = Z;
		19'b1101011100101101011: color_data = Z;
		19'b1101011100101101100: color_data = Z;
		19'b1101011100101101101: color_data = Z;
		19'b1101011100101101110: color_data = Z;
		19'b1101011110100100110: color_data = Z;
		19'b1101011110100100111: color_data = Z;
		19'b1101011110100101000: color_data = Z;
		19'b1101011110100101001: color_data = Z;
		19'b1101011110100101010: color_data = Z;
		19'b1101011110100101011: color_data = Z;
		19'b1101011110100101100: color_data = Z;
		19'b1101011110100101101: color_data = Z;
		19'b1101011110100101110: color_data = Z;
		19'b1101011110100101111: color_data = Z;
		19'b1101011110100110000: color_data = Z;
		19'b1101011110100110001: color_data = Z;
		19'b1101011110100110010: color_data = Z;
		19'b1101011110100110011: color_data = Z;
		19'b1101011110100110100: color_data = Z;
		19'b1101011110100110101: color_data = Z;
		19'b1101011110100110110: color_data = Z;
		19'b1101011110100110111: color_data = Z;
		19'b1101011110100111000: color_data = Z;
		19'b1101011110100111001: color_data = Z;
		19'b1101011110100111010: color_data = Z;
		19'b1101011110100111011: color_data = Z;
		19'b1101011110101001001: color_data = Z;
		19'b1101011110101001010: color_data = Z;
		19'b1101011110101001011: color_data = Z;
		19'b1101011110101001100: color_data = Z;
		19'b1101011110101001101: color_data = Z;
		19'b1101011110101001110: color_data = Z;
		19'b1101011110101001111: color_data = Z;
		19'b1101011110101010000: color_data = Z;
		19'b1101011110101010001: color_data = Z;
		19'b1101011110101010010: color_data = Z;
		19'b1101011110101010011: color_data = Z;
		19'b1101011110101010100: color_data = Z;
		19'b1101011110101010101: color_data = Z;
		19'b1101011110101010110: color_data = Z;
		19'b1101011110101010111: color_data = Z;
		19'b1101011110101011000: color_data = Z;
		19'b1101011110101011001: color_data = Z;
		19'b1101011110101011010: color_data = Z;
		19'b1101011110101011011: color_data = Z;
		19'b1101011110101011100: color_data = Z;
		19'b1101011110101011101: color_data = Z;
		19'b1101011110101011110: color_data = Z;
		19'b1101011110101011111: color_data = Z;
		19'b1101011110101100000: color_data = Z;
		19'b1101011110101100001: color_data = Z;
		19'b1101011110101100010: color_data = Z;
		19'b1101011110101100011: color_data = Z;
		19'b1101011110101100100: color_data = Z;
		19'b1101011110101100101: color_data = Z;
		19'b1101011110101100110: color_data = Z;
		19'b1101011110101100111: color_data = Z;
		19'b1101011110101101000: color_data = Z;
		19'b1101011110101101001: color_data = Z;
		19'b1101011110101101010: color_data = Z;
		19'b1101011110101101011: color_data = Z;
		19'b1101011110101101100: color_data = Z;
		19'b1101011110101101101: color_data = Z;
		19'b1101011110101101110: color_data = Z;
		19'b1101100000100100110: color_data = Z;
		19'b1101100000100100111: color_data = Z;
		19'b1101100000100101000: color_data = Z;
		19'b1101100000100101001: color_data = Z;
		19'b1101100000100101010: color_data = Z;
		19'b1101100000100101011: color_data = Z;
		19'b1101100000100101100: color_data = Z;
		19'b1101100000100101101: color_data = Z;
		19'b1101100000100101110: color_data = Z;
		19'b1101100000100101111: color_data = Z;
		19'b1101100000100110000: color_data = Z;
		19'b1101100000100110001: color_data = Z;
		19'b1101100000100110010: color_data = Z;
		19'b1101100000100110011: color_data = Z;
		19'b1101100000100110100: color_data = Z;
		19'b1101100000100110101: color_data = Z;
		19'b1101100000100110110: color_data = Z;
		19'b1101100000100110111: color_data = Z;
		19'b1101100000100111000: color_data = Z;
		19'b1101100000100111001: color_data = Z;
		19'b1101100000100111010: color_data = Z;
		19'b1101100000100111011: color_data = Z;
		19'b1101100000100111100: color_data = Z;
		19'b1101100000100111101: color_data = Z;
		19'b1101100000100111110: color_data = Z;
		19'b1101100000100111111: color_data = Z;
		19'b1101100000101000000: color_data = Z;
		19'b1101100000101000001: color_data = Z;
		19'b1101100000101000011: color_data = Z;
		19'b1101100000101000100: color_data = Z;
		19'b1101100000101000101: color_data = Z;
		19'b1101100000101000110: color_data = Z;
		19'b1101100000101000111: color_data = Z;
		19'b1101100000101001000: color_data = Z;
		19'b1101100000101001001: color_data = Z;
		19'b1101100000101001010: color_data = Z;
		19'b1101100000101001011: color_data = Z;
		19'b1101100000101001100: color_data = Z;
		19'b1101100000101001101: color_data = Z;
		19'b1101100000101001110: color_data = Z;
		19'b1101100000101001111: color_data = Z;
		19'b1101100000101010000: color_data = Z;
		19'b1101100000101010001: color_data = Z;
		19'b1101100000101010010: color_data = Z;
		19'b1101100000101010011: color_data = Z;
		19'b1101100000101010100: color_data = Z;
		19'b1101100000101010101: color_data = Z;
		19'b1101100000101010110: color_data = Z;
		19'b1101100000101010111: color_data = Z;
		19'b1101100000101011000: color_data = Z;
		19'b1101100000101011001: color_data = Z;
		19'b1101100000101011010: color_data = Z;
		19'b1101100000101011011: color_data = Z;
		19'b1101100000101011100: color_data = Z;
		19'b1101100000101011101: color_data = Z;
		19'b1101100000101011110: color_data = Z;
		19'b1101100000101011111: color_data = Z;
		19'b1101100000101100000: color_data = Z;
		19'b1101100000101100001: color_data = Z;
		19'b1101100000101100010: color_data = Z;
		19'b1101100000101100011: color_data = Z;
		19'b1101100000101100100: color_data = Z;
		19'b1101100000101100101: color_data = Z;
		19'b1101100000101100110: color_data = Z;
		19'b1101100000101100111: color_data = Z;
		19'b1101100000101101000: color_data = Z;
		19'b1101100000101101001: color_data = Z;
		19'b1101100000101101010: color_data = Z;
		19'b1101100000101101011: color_data = Z;
		19'b1101100000101101100: color_data = Z;
		19'b1101100000101101101: color_data = Z;
		19'b1101100000101101110: color_data = Z;
		19'b1101100010100100110: color_data = Z;
		19'b1101100010100100111: color_data = Z;
		19'b1101100010100101000: color_data = Z;
		19'b1101100010100101001: color_data = Z;
		19'b1101100010100101010: color_data = Z;
		19'b1101100010100101011: color_data = Z;
		19'b1101100010100101100: color_data = Z;
		19'b1101100010100101101: color_data = Z;
		19'b1101100010100101110: color_data = Z;
		19'b1101100010100101111: color_data = Z;
		19'b1101100010100110000: color_data = Z;
		19'b1101100010100110001: color_data = Z;
		19'b1101100010100110010: color_data = Z;
		19'b1101100010100110011: color_data = Z;
		19'b1101100010100110100: color_data = Z;
		19'b1101100010100110101: color_data = Z;
		19'b1101100010100110110: color_data = Z;
		19'b1101100010100110111: color_data = Z;
		19'b1101100010100111000: color_data = Z;
		19'b1101100010100111001: color_data = Z;
		19'b1101100010100111010: color_data = Z;
		19'b1101100010100111011: color_data = Z;
		19'b1101100010100111100: color_data = Z;
		19'b1101100010100111101: color_data = Z;
		19'b1101100010100111110: color_data = Z;
		19'b1101100010100111111: color_data = Z;
		19'b1101100010101000000: color_data = Z;
		19'b1101100010101000001: color_data = Z;
		19'b1101100010101000010: color_data = Z;
		19'b1101100010101000011: color_data = Z;
		19'b1101100010101000100: color_data = Z;
		19'b1101100010101000101: color_data = Z;
		19'b1101100010101000110: color_data = Z;
		19'b1101100010101000111: color_data = Z;
		19'b1101100010101001000: color_data = Z;
		19'b1101100010101001001: color_data = Z;
		19'b1101100010101001010: color_data = Z;
		19'b1101100010101001011: color_data = Z;
		19'b1101100010101001100: color_data = Z;
		19'b1101100010101001101: color_data = Z;
		19'b1101100010101001110: color_data = Z;
		19'b1101100010101001111: color_data = Z;
		19'b1101100010101010000: color_data = Z;
		19'b1101100010101010001: color_data = Z;
		19'b1101100010101010010: color_data = Z;
		19'b1101100010101010011: color_data = Z;
		19'b1101100010101010100: color_data = Z;
		19'b1101100010101010101: color_data = Z;
		19'b1101100010101010110: color_data = Z;
		19'b1101100010101010111: color_data = Z;
		19'b1101100010101011000: color_data = Z;
		19'b1101100010101011001: color_data = Z;
		19'b1101100010101011010: color_data = Z;
		19'b1101100010101011011: color_data = Z;
		19'b1101100010101011100: color_data = Z;
		19'b1101100010101011101: color_data = Z;
		19'b1101100010101011110: color_data = Z;
		19'b1101100010101011111: color_data = Z;
		19'b1101100010101100000: color_data = Z;
		19'b1101100010101100001: color_data = Z;
		19'b1101100010101100010: color_data = Z;
		19'b1101100010101100011: color_data = Z;
		19'b1101100010101100100: color_data = Z;
		19'b1101100010101100101: color_data = Z;
		19'b1101100010101100110: color_data = Z;
		19'b1101100010101100111: color_data = Z;
		19'b1101100010101101000: color_data = Z;
		19'b1101100010101101001: color_data = Z;
		19'b1101100010101101010: color_data = Z;
		19'b1101100010101101011: color_data = Z;
		19'b1101100010101101100: color_data = Z;
		19'b1101100010101101101: color_data = Z;
		19'b1101100010101101110: color_data = Z;
		19'b1101100100100100110: color_data = Z;
		19'b1101100100100100111: color_data = Z;
		19'b1101100100100101000: color_data = Z;
		19'b1101100100100101001: color_data = Z;
		19'b1101100100100101010: color_data = Z;
		19'b1101100100100101011: color_data = Z;
		19'b1101100100100101100: color_data = Z;
		19'b1101100100100101101: color_data = Z;
		19'b1101100100100101110: color_data = Z;
		19'b1101100100100101111: color_data = Z;
		19'b1101100100100110000: color_data = Z;
		19'b1101100100100110001: color_data = Z;
		19'b1101100100100110010: color_data = Z;
		19'b1101100100100110011: color_data = Z;
		19'b1101100100100110100: color_data = Z;
		19'b1101100100100110101: color_data = Z;
		19'b1101100100100110110: color_data = Z;
		19'b1101100100100110111: color_data = Z;
		19'b1101100100100111000: color_data = Z;
		19'b1101100100100111001: color_data = Z;
		19'b1101100100100111010: color_data = Z;
		19'b1101100100100111011: color_data = Z;
		19'b1101100100100111100: color_data = Z;
		19'b1101100100100111101: color_data = Z;
		19'b1101100100100111110: color_data = Z;
		19'b1101100100100111111: color_data = Z;
		19'b1101100100101000000: color_data = Z;
		19'b1101100100101000001: color_data = Z;
		19'b1101100100101000010: color_data = Z;
		19'b1101100100101000011: color_data = Z;
		19'b1101100100101000100: color_data = Z;
		19'b1101100100101000101: color_data = Z;
		19'b1101100100101000110: color_data = Z;
		19'b1101100100101000111: color_data = Z;
		19'b1101100100101001000: color_data = Z;
		19'b1101100100101001001: color_data = Z;
		19'b1101100100101001010: color_data = Z;
		19'b1101100100101001011: color_data = Z;
		19'b1101100100101001100: color_data = Z;
		19'b1101100100101001101: color_data = Z;
		19'b1101100100101001110: color_data = Z;
		19'b1101100100101001111: color_data = Z;
		19'b1101100100101010000: color_data = Z;
		19'b1101100100101010001: color_data = Z;
		19'b1101100100101010010: color_data = Z;
		19'b1101100100101010011: color_data = Z;
		19'b1101100100101010100: color_data = Z;
		19'b1101100100101010101: color_data = Z;
		19'b1101100100101010110: color_data = Z;
		19'b1101100100101010111: color_data = Z;
		19'b1101100100101011000: color_data = Z;
		19'b1101100100101011001: color_data = Z;
		19'b1101100100101011010: color_data = Z;
		19'b1101100100101011011: color_data = Z;
		19'b1101100100101011100: color_data = Z;
		19'b1101100100101011101: color_data = Z;
		19'b1101100100101011110: color_data = Z;
		19'b1101100100101011111: color_data = Z;
		19'b1101100100101100000: color_data = Z;
		19'b1101100100101100001: color_data = Z;
		19'b1101100100101100010: color_data = Z;
		19'b1101100100101100011: color_data = Z;
		19'b1101100100101100100: color_data = Z;
		19'b1101100100101100101: color_data = Z;
		19'b1101100100101100110: color_data = Z;
		19'b1101100100101100111: color_data = Z;
		19'b1101100100101101000: color_data = Z;
		19'b1101100100101101001: color_data = Z;
		19'b1101100100101101010: color_data = Z;
		19'b1101100100101101011: color_data = Z;
		19'b1101100100101101100: color_data = Z;
		19'b1101100100101101101: color_data = Z;
		19'b1101100100101101110: color_data = Z;
		19'b1101100110100011010: color_data = Z;
		19'b1101100110100100110: color_data = Z;
		19'b1101100110100100111: color_data = Z;
		19'b1101100110100101000: color_data = Z;
		19'b1101100110100101001: color_data = Z;
		19'b1101100110100101010: color_data = Z;
		19'b1101100110100101011: color_data = Z;
		19'b1101100110100101100: color_data = Z;
		19'b1101100110100101101: color_data = Z;
		19'b1101100110100101110: color_data = Z;
		19'b1101100110100101111: color_data = Z;
		19'b1101100110100110000: color_data = Z;
		19'b1101100110100110001: color_data = Z;
		19'b1101100110100110010: color_data = Z;
		19'b1101100110100110011: color_data = Z;
		19'b1101100110100110100: color_data = Z;
		19'b1101100110100110101: color_data = Z;
		19'b1101100110100110110: color_data = Z;
		19'b1101100110100110111: color_data = Z;
		19'b1101100110100111000: color_data = Z;
		19'b1101100110100111001: color_data = Z;
		19'b1101100110100111010: color_data = Z;
		19'b1101100110100111011: color_data = Z;
		19'b1101100110100111100: color_data = Z;
		19'b1101100110100111101: color_data = Z;
		19'b1101100110100111110: color_data = Z;
		19'b1101100110100111111: color_data = Z;
		19'b1101100110101000000: color_data = Z;
		19'b1101100110101000001: color_data = Z;
		19'b1101100110101000010: color_data = Z;
		19'b1101100110101000011: color_data = Z;
		19'b1101100110101000100: color_data = Z;
		19'b1101100110101000101: color_data = Z;
		19'b1101100110101000110: color_data = Z;
		19'b1101100110101000111: color_data = Z;
		19'b1101100110101001000: color_data = Z;
		19'b1101100110101001001: color_data = Z;
		19'b1101100110101001010: color_data = Z;
		19'b1101100110101001011: color_data = Z;
		19'b1101100110101001100: color_data = Z;
		19'b1101100110101001101: color_data = Z;
		19'b1101100110101001110: color_data = Z;
		19'b1101100110101001111: color_data = Z;
		19'b1101100110101010000: color_data = Z;
		19'b1101100110101010001: color_data = Z;
		19'b1101100110101010010: color_data = Z;
		19'b1101100110101010011: color_data = Z;
		19'b1101100110101010100: color_data = Z;
		19'b1101100110101010101: color_data = Z;
		19'b1101100110101010110: color_data = Z;
		19'b1101100110101010111: color_data = Z;
		19'b1101100110101011000: color_data = Z;
		19'b1101100110101011001: color_data = Z;
		19'b1101100110101011010: color_data = Z;
		19'b1101100110101011011: color_data = Z;
		19'b1101100110101011100: color_data = Z;
		19'b1101100110101011101: color_data = Z;
		19'b1101100110101011110: color_data = Z;
		19'b1101100110101011111: color_data = Z;
		19'b1101100110101100000: color_data = Z;
		19'b1101100110101100001: color_data = Z;
		19'b1101100110101100010: color_data = Z;
		19'b1101100110101100011: color_data = Z;
		19'b1101100110101100100: color_data = Z;
		19'b1101100110101100101: color_data = Z;
		19'b1101100110101100110: color_data = Z;
		19'b1101100110101100111: color_data = Z;
		19'b1101100110101101000: color_data = Z;
		19'b1101100110101101001: color_data = Z;
		19'b1101100110101101010: color_data = Z;
		19'b1101100110101101011: color_data = Z;
		19'b1101100110101101100: color_data = Z;
		19'b1101100110101101101: color_data = Z;
		19'b1101101000100011010: color_data = Z;
		19'b1101101000100100101: color_data = Z;
		19'b1101101000100100110: color_data = Z;
		19'b1101101000100100111: color_data = Z;
		19'b1101101000100101000: color_data = Z;
		19'b1101101000100101001: color_data = Z;
		19'b1101101000100101010: color_data = Z;
		19'b1101101000100101011: color_data = Z;
		19'b1101101000100101100: color_data = Z;
		19'b1101101000100101101: color_data = Z;
		19'b1101101000100101110: color_data = Z;
		19'b1101101000100101111: color_data = Z;
		19'b1101101000100110000: color_data = Z;
		19'b1101101000100110001: color_data = Z;
		19'b1101101000100110010: color_data = Z;
		19'b1101101000100110011: color_data = Z;
		19'b1101101000100110100: color_data = Z;
		19'b1101101000100110101: color_data = Z;
		19'b1101101000100110110: color_data = Z;
		19'b1101101000100110111: color_data = Z;
		19'b1101101000100111000: color_data = Z;
		19'b1101101000100111001: color_data = Z;
		19'b1101101000100111010: color_data = Z;
		19'b1101101000100111011: color_data = Z;
		19'b1101101000100111100: color_data = Z;
		19'b1101101000100111101: color_data = Z;
		19'b1101101000100111110: color_data = Z;
		19'b1101101000100111111: color_data = Z;
		19'b1101101000101000000: color_data = Z;
		19'b1101101000101000001: color_data = Z;
		19'b1101101000101000010: color_data = Z;
		19'b1101101000101000011: color_data = Z;
		19'b1101101000101000100: color_data = Z;
		19'b1101101000101000101: color_data = Z;
		19'b1101101000101000110: color_data = Z;
		19'b1101101000101000111: color_data = Z;
		19'b1101101000101001000: color_data = Z;
		19'b1101101000101001001: color_data = Z;
		19'b1101101000101001010: color_data = Z;
		19'b1101101000101001011: color_data = Z;
		19'b1101101000101001100: color_data = Z;
		19'b1101101000101001101: color_data = Z;
		19'b1101101000101001110: color_data = Z;
		19'b1101101000101001111: color_data = Z;
		19'b1101101000101010000: color_data = Z;
		19'b1101101000101010001: color_data = Z;
		19'b1101101000101010010: color_data = Z;
		19'b1101101000101010011: color_data = Z;
		19'b1101101000101010100: color_data = Z;
		19'b1101101000101010101: color_data = Z;
		19'b1101101000101010110: color_data = Z;
		19'b1101101000101010111: color_data = Z;
		19'b1101101000101011000: color_data = Z;
		19'b1101101000101011001: color_data = Z;
		19'b1101101000101011010: color_data = Z;
		19'b1101101000101011011: color_data = Z;
		19'b1101101000101011100: color_data = Z;
		19'b1101101000101011101: color_data = Z;
		19'b1101101000101011110: color_data = Z;
		19'b1101101000101011111: color_data = Z;
		19'b1101101000101100000: color_data = Z;
		19'b1101101000101100001: color_data = Z;
		19'b1101101000101100010: color_data = Z;
		19'b1101101000101100011: color_data = Z;
		19'b1101101000101100100: color_data = Z;
		19'b1101101000101100101: color_data = Z;
		19'b1101101000101100110: color_data = Z;
		19'b1101101000101100111: color_data = Z;
		19'b1101101000101101000: color_data = Z;
		19'b1101101000101101001: color_data = Z;
		19'b1101101000101101010: color_data = Z;
		19'b1101101000101101011: color_data = Z;
		19'b1101101000101101100: color_data = Z;
		19'b1101101000101101101: color_data = Z;
		19'b1101101000101101110: color_data = Z;
		19'b1101101000101101111: color_data = Z;
		19'b1101101000101110000: color_data = Z;
		19'b1101101010100011011: color_data = Z;
		19'b1101101010100100101: color_data = Z;
		19'b1101101010100100110: color_data = Z;
		19'b1101101010100100111: color_data = Z;
		19'b1101101010100101000: color_data = Z;
		19'b1101101010100101001: color_data = Z;
		19'b1101101010100101010: color_data = Z;
		19'b1101101010100101011: color_data = Z;
		19'b1101101010100101100: color_data = Z;
		19'b1101101010100101101: color_data = Z;
		19'b1101101010100101110: color_data = Z;
		19'b1101101010100101111: color_data = Z;
		19'b1101101010100110000: color_data = Z;
		19'b1101101010100110001: color_data = Z;
		19'b1101101010100110010: color_data = Z;
		19'b1101101010100110011: color_data = Z;
		19'b1101101010100110100: color_data = Z;
		19'b1101101010100110101: color_data = Z;
		19'b1101101010100110110: color_data = Z;
		19'b1101101010100110111: color_data = Z;
		19'b1101101010100111000: color_data = Z;
		19'b1101101010100111001: color_data = Z;
		19'b1101101010100111010: color_data = Z;
		19'b1101101010100111011: color_data = Z;
		19'b1101101010100111100: color_data = Z;
		19'b1101101010100111101: color_data = Z;
		19'b1101101010100111110: color_data = Z;
		19'b1101101010100111111: color_data = Z;
		19'b1101101010101000000: color_data = Z;
		19'b1101101010101000001: color_data = Z;
		19'b1101101010101000010: color_data = Z;
		19'b1101101010101000011: color_data = Z;
		19'b1101101010101000100: color_data = Z;
		19'b1101101010101000101: color_data = Z;
		19'b1101101010101000110: color_data = Z;
		19'b1101101010101000111: color_data = Z;
		19'b1101101010101001000: color_data = Z;
		19'b1101101010101001001: color_data = Z;
		19'b1101101010101001010: color_data = Z;
		19'b1101101010101001011: color_data = Z;
		19'b1101101010101001100: color_data = Z;
		19'b1101101010101001101: color_data = Z;
		19'b1101101010101001110: color_data = Z;
		19'b1101101010101001111: color_data = Z;
		19'b1101101010101010000: color_data = Z;
		19'b1101101010101010001: color_data = Z;
		19'b1101101010101010010: color_data = Z;
		19'b1101101010101010011: color_data = Z;
		19'b1101101010101010100: color_data = Z;
		19'b1101101010101010101: color_data = Z;
		19'b1101101010101010110: color_data = Z;
		19'b1101101010101010111: color_data = Z;
		19'b1101101010101011000: color_data = Z;
		19'b1101101010101011001: color_data = Z;
		19'b1101101010101011010: color_data = Z;
		19'b1101101010101011011: color_data = Z;
		19'b1101101010101011100: color_data = Z;
		19'b1101101010101011101: color_data = Z;
		19'b1101101010101011110: color_data = Z;
		19'b1101101010101011111: color_data = Z;
		19'b1101101010101100000: color_data = Z;
		19'b1101101010101100001: color_data = Z;
		19'b1101101010101100010: color_data = Z;
		19'b1101101010101100011: color_data = Z;
		19'b1101101010101100100: color_data = Z;
		19'b1101101010101100101: color_data = Z;
		19'b1101101010101100110: color_data = Z;
		19'b1101101010101100111: color_data = Z;
		19'b1101101010101101000: color_data = Z;
		19'b1101101010101101001: color_data = Z;
		19'b1101101010101101010: color_data = Z;
		19'b1101101010101101011: color_data = Z;
		19'b1101101010101101100: color_data = Z;
		19'b1101101010101101101: color_data = Z;
		19'b1101101010101101110: color_data = Z;
		19'b1101101010101101111: color_data = Z;
		19'b1101101010101110000: color_data = Z;
		19'b1101101100100011011: color_data = Z;
		19'b1101101100100100101: color_data = Z;
		19'b1101101100100100110: color_data = Z;
		19'b1101101100100100111: color_data = Z;
		19'b1101101100100101000: color_data = Z;
		19'b1101101100100101001: color_data = Z;
		19'b1101101100100101010: color_data = Z;
		19'b1101101100100101011: color_data = Z;
		19'b1101101100100101100: color_data = Z;
		19'b1101101100100101101: color_data = Z;
		19'b1101101100100101110: color_data = Z;
		19'b1101101100100101111: color_data = Z;
		19'b1101101100100110000: color_data = Z;
		19'b1101101100100110001: color_data = Z;
		19'b1101101100100110010: color_data = Z;
		19'b1101101100100110011: color_data = Z;
		19'b1101101100100110100: color_data = Z;
		19'b1101101100100110101: color_data = Z;
		19'b1101101100100110110: color_data = Z;
		19'b1101101100100110111: color_data = Z;
		19'b1101101100100111000: color_data = Z;
		19'b1101101100100111001: color_data = Z;
		19'b1101101100100111010: color_data = Z;
		19'b1101101100100111011: color_data = Z;
		19'b1101101100100111100: color_data = Z;
		19'b1101101100100111101: color_data = Z;
		19'b1101101100100111110: color_data = Z;
		19'b1101101100100111111: color_data = Z;
		19'b1101101100101000000: color_data = Z;
		19'b1101101100101000001: color_data = Z;
		19'b1101101100101000010: color_data = Z;
		19'b1101101100101000011: color_data = Z;
		19'b1101101100101000100: color_data = Z;
		19'b1101101100101000101: color_data = Z;
		19'b1101101100101000110: color_data = Z;
		19'b1101101100101000111: color_data = Z;
		19'b1101101100101001000: color_data = Z;
		19'b1101101100101001001: color_data = Z;
		19'b1101101100101001010: color_data = Z;
		19'b1101101100101001011: color_data = Z;
		19'b1101101100101001100: color_data = Z;
		19'b1101101100101001101: color_data = Z;
		19'b1101101100101001110: color_data = Z;
		19'b1101101100101001111: color_data = Z;
		19'b1101101100101010000: color_data = Z;
		19'b1101101100101010001: color_data = Z;
		19'b1101101100101010010: color_data = Z;
		19'b1101101100101010011: color_data = Z;
		19'b1101101100101010100: color_data = Z;
		19'b1101101100101010101: color_data = Z;
		19'b1101101100101010110: color_data = Z;
		19'b1101101100101010111: color_data = Z;
		19'b1101101100101011000: color_data = Z;
		19'b1101101100101011001: color_data = Z;
		19'b1101101100101011010: color_data = Z;
		19'b1101101100101011011: color_data = Z;
		19'b1101101100101011100: color_data = Z;
		19'b1101101100101011101: color_data = Z;
		19'b1101101100101011110: color_data = Z;
		19'b1101101100101011111: color_data = Z;
		19'b1101101100101100000: color_data = Z;
		19'b1101101100101100001: color_data = Z;
		19'b1101101100101100010: color_data = Z;
		19'b1101101100101100011: color_data = Z;
		19'b1101101100101100100: color_data = Z;
		19'b1101101100101100101: color_data = Z;
		19'b1101101100101100110: color_data = Z;
		19'b1101101100101100111: color_data = Z;
		19'b1101101100101101000: color_data = Z;
		19'b1101101100101101001: color_data = Z;
		19'b1101101100101101010: color_data = Z;
		19'b1101101100101101011: color_data = Z;
		19'b1101101100101101100: color_data = Z;
		19'b1101101100101101101: color_data = Z;
		19'b1101101100101101110: color_data = Z;
		19'b1101101100101101111: color_data = Z;
		19'b1101101100101110000: color_data = Z;
		19'b1101101100101110001: color_data = Z;
		19'b1101101110100011011: color_data = Z;
		19'b1101101110100100101: color_data = Z;
		19'b1101101110100100110: color_data = Z;
		19'b1101101110100100111: color_data = Z;
		19'b1101101110100101000: color_data = Z;
		19'b1101101110100101001: color_data = Z;
		19'b1101101110100101010: color_data = Z;
		19'b1101101110100101011: color_data = Z;
		19'b1101101110100101100: color_data = Z;
		19'b1101101110100101101: color_data = Z;
		19'b1101101110100101110: color_data = Z;
		19'b1101101110100101111: color_data = Z;
		19'b1101101110100110000: color_data = Z;
		19'b1101101110100110001: color_data = Z;
		19'b1101101110100110010: color_data = Z;
		19'b1101101110100110011: color_data = Z;
		19'b1101101110100110100: color_data = Z;
		19'b1101101110100110101: color_data = Z;
		19'b1101101110100110110: color_data = Z;
		19'b1101101110100110111: color_data = Z;
		19'b1101101110100111000: color_data = Z;
		19'b1101101110100111001: color_data = Z;
		19'b1101101110100111010: color_data = Z;
		19'b1101101110100111011: color_data = Z;
		19'b1101101110100111100: color_data = Z;
		19'b1101101110100111101: color_data = Z;
		19'b1101101110100111110: color_data = Z;
		19'b1101101110100111111: color_data = Z;
		19'b1101101110101000000: color_data = Z;
		19'b1101101110101000001: color_data = Z;
		19'b1101101110101000010: color_data = Z;
		19'b1101101110101000011: color_data = Z;
		19'b1101101110101000100: color_data = Z;
		19'b1101101110101000101: color_data = Z;
		19'b1101101110101000110: color_data = Z;
		19'b1101101110101000111: color_data = Z;
		19'b1101101110101001000: color_data = Z;
		19'b1101101110101001001: color_data = Z;
		19'b1101101110101001010: color_data = Z;
		19'b1101101110101001011: color_data = Z;
		19'b1101101110101001100: color_data = Z;
		19'b1101101110101001101: color_data = Z;
		19'b1101101110101001110: color_data = Z;
		19'b1101101110101001111: color_data = Z;
		19'b1101101110101010000: color_data = Z;
		19'b1101101110101010001: color_data = Z;
		19'b1101101110101010010: color_data = Z;
		19'b1101101110101010011: color_data = Z;
		19'b1101101110101010100: color_data = Z;
		19'b1101101110101010101: color_data = Z;
		19'b1101101110101010110: color_data = Z;
		19'b1101101110101010111: color_data = Z;
		19'b1101101110101011000: color_data = Z;
		19'b1101101110101011001: color_data = Z;
		19'b1101101110101011010: color_data = Z;
		19'b1101101110101011011: color_data = Z;
		19'b1101101110101011100: color_data = Z;
		19'b1101101110101011101: color_data = Z;
		19'b1101101110101011110: color_data = Z;
		19'b1101101110101011111: color_data = Z;
		19'b1101101110101100000: color_data = Z;
		19'b1101101110101100001: color_data = Z;
		19'b1101101110101100010: color_data = Z;
		19'b1101101110101100011: color_data = Z;
		19'b1101101110101100100: color_data = Z;
		19'b1101101110101100101: color_data = Z;
		19'b1101101110101100110: color_data = Z;
		19'b1101101110101100111: color_data = Z;
		19'b1101101110101101000: color_data = Z;
		19'b1101101110101101001: color_data = Z;
		19'b1101101110101101010: color_data = Z;
		19'b1101101110101101011: color_data = Z;
		19'b1101101110101101100: color_data = Z;
		19'b1101101110101101101: color_data = Z;
		19'b1101101110101101110: color_data = Z;
		19'b1101101110101101111: color_data = Z;
		19'b1101101110101110000: color_data = Z;
		19'b1101101110101110001: color_data = Z;
		19'b1101101110101110010: color_data = Z;
		19'b1101110000100011011: color_data = Z;
		19'b1101110000100011100: color_data = Z;
		19'b1101110000100100101: color_data = Z;
		19'b1101110000100100110: color_data = Z;
		19'b1101110000100100111: color_data = Z;
		19'b1101110000100101000: color_data = Z;
		19'b1101110000100101001: color_data = Z;
		19'b1101110000100101010: color_data = Z;
		19'b1101110000100101011: color_data = Z;
		19'b1101110000100101100: color_data = Z;
		19'b1101110000100101101: color_data = Z;
		19'b1101110000100101110: color_data = Z;
		19'b1101110000100101111: color_data = Z;
		19'b1101110000100110000: color_data = Z;
		19'b1101110000100110001: color_data = Z;
		19'b1101110000100110010: color_data = Z;
		19'b1101110000100110011: color_data = Z;
		19'b1101110000100110100: color_data = Z;
		19'b1101110000100110101: color_data = Z;
		19'b1101110000100110110: color_data = Z;
		19'b1101110000100110111: color_data = Z;
		19'b1101110000100111000: color_data = Z;
		19'b1101110000100111001: color_data = Z;
		19'b1101110000100111010: color_data = Z;
		19'b1101110000100111011: color_data = Z;
		19'b1101110000100111100: color_data = Z;
		19'b1101110000100111101: color_data = Z;
		19'b1101110000100111110: color_data = Z;
		19'b1101110000100111111: color_data = Z;
		19'b1101110000101000000: color_data = Z;
		19'b1101110000101000001: color_data = Z;
		19'b1101110000101000010: color_data = Z;
		19'b1101110000101000011: color_data = Z;
		19'b1101110000101000100: color_data = Z;
		19'b1101110000101000101: color_data = Z;
		19'b1101110000101000110: color_data = Z;
		19'b1101110000101000111: color_data = Z;
		19'b1101110000101001000: color_data = Z;
		19'b1101110000101001001: color_data = Z;
		19'b1101110000101001010: color_data = Z;
		19'b1101110000101001011: color_data = Z;
		19'b1101110000101001100: color_data = Z;
		19'b1101110000101001101: color_data = Z;
		19'b1101110000101001110: color_data = Z;
		19'b1101110000101001111: color_data = Z;
		19'b1101110000101010000: color_data = Z;
		19'b1101110000101010001: color_data = Z;
		19'b1101110000101010010: color_data = Z;
		19'b1101110000101010011: color_data = Z;
		19'b1101110000101010100: color_data = Z;
		19'b1101110000101010101: color_data = Z;
		19'b1101110000101010110: color_data = Z;
		19'b1101110000101010111: color_data = Z;
		19'b1101110000101011000: color_data = Z;
		19'b1101110000101011001: color_data = Z;
		19'b1101110000101011010: color_data = Z;
		19'b1101110000101011011: color_data = Z;
		19'b1101110000101011100: color_data = Z;
		19'b1101110000101011101: color_data = Z;
		19'b1101110000101011110: color_data = Z;
		19'b1101110000101011111: color_data = Z;
		19'b1101110000101100000: color_data = Z;
		19'b1101110000101100001: color_data = Z;
		19'b1101110000101100010: color_data = Z;
		19'b1101110000101100011: color_data = Z;
		19'b1101110000101100100: color_data = Z;
		19'b1101110000101100101: color_data = Z;
		19'b1101110000101100110: color_data = Z;
		19'b1101110000101100111: color_data = Z;
		19'b1101110000101101000: color_data = Z;
		19'b1101110000101101001: color_data = Z;
		19'b1101110000101101010: color_data = Z;
		19'b1101110000101101011: color_data = Z;
		19'b1101110000101101100: color_data = Z;
		19'b1101110000101101101: color_data = Z;
		19'b1101110000101101110: color_data = Z;
		19'b1101110000101101111: color_data = Z;
		19'b1101110000101110000: color_data = Z;
		19'b1101110000101110001: color_data = Z;
		19'b1101110000101110111: color_data = Z;
		19'b1101110010100011100: color_data = Z;
		19'b1101110010100100101: color_data = Z;
		19'b1101110010100100110: color_data = Z;
		19'b1101110010100100111: color_data = Z;
		19'b1101110010100101000: color_data = Z;
		19'b1101110010100101001: color_data = Z;
		19'b1101110010100101010: color_data = Z;
		19'b1101110010100101011: color_data = Z;
		19'b1101110010100101100: color_data = Z;
		19'b1101110010100101101: color_data = Z;
		19'b1101110010100101110: color_data = Z;
		19'b1101110010100101111: color_data = Z;
		19'b1101110010100110000: color_data = Z;
		19'b1101110010100110001: color_data = Z;
		19'b1101110010100110010: color_data = Z;
		19'b1101110010100110011: color_data = Z;
		19'b1101110010100110100: color_data = Z;
		19'b1101110010100110101: color_data = Z;
		19'b1101110010100110110: color_data = Z;
		19'b1101110010100110111: color_data = Z;
		19'b1101110010100111000: color_data = Z;
		19'b1101110010100111001: color_data = Z;
		19'b1101110010100111010: color_data = Z;
		19'b1101110010100111011: color_data = Z;
		19'b1101110010100111100: color_data = Z;
		19'b1101110010100111101: color_data = Z;
		19'b1101110010100111110: color_data = Z;
		19'b1101110010100111111: color_data = Z;
		19'b1101110010101000000: color_data = Z;
		19'b1101110010101000001: color_data = Z;
		19'b1101110010101000010: color_data = Z;
		19'b1101110010101000011: color_data = Z;
		19'b1101110010101000100: color_data = Z;
		19'b1101110010101000101: color_data = Z;
		19'b1101110010101000110: color_data = Z;
		19'b1101110010101000111: color_data = Z;
		19'b1101110010101001000: color_data = Z;
		19'b1101110010101001001: color_data = Z;
		19'b1101110010101001010: color_data = Z;
		19'b1101110010101001011: color_data = Z;
		19'b1101110010101001100: color_data = Z;
		19'b1101110010101001101: color_data = Z;
		19'b1101110010101001110: color_data = Z;
		19'b1101110010101001111: color_data = Z;
		19'b1101110010101010000: color_data = Z;
		19'b1101110010101010001: color_data = Z;
		19'b1101110010101010010: color_data = Z;
		19'b1101110010101010011: color_data = Z;
		19'b1101110010101010100: color_data = Z;
		19'b1101110010101010101: color_data = Z;
		19'b1101110010101010110: color_data = Z;
		19'b1101110010101010111: color_data = Z;
		19'b1101110010101011000: color_data = Z;
		19'b1101110010101011001: color_data = Z;
		19'b1101110010101011010: color_data = Z;
		19'b1101110010101011011: color_data = Z;
		19'b1101110010101011100: color_data = Z;
		19'b1101110010101011101: color_data = Z;
		19'b1101110010101011110: color_data = Z;
		19'b1101110010101011111: color_data = Z;
		19'b1101110010101100000: color_data = Z;
		19'b1101110010101100001: color_data = Z;
		19'b1101110010101100010: color_data = Z;
		19'b1101110010101100011: color_data = Z;
		19'b1101110010101100100: color_data = Z;
		19'b1101110010101100101: color_data = Z;
		19'b1101110010101100110: color_data = Z;
		19'b1101110010101100111: color_data = Z;
		19'b1101110010101101000: color_data = Z;
		19'b1101110010101101001: color_data = Z;
		19'b1101110010101101010: color_data = Z;
		19'b1101110010101101011: color_data = Z;
		19'b1101110010101101100: color_data = Z;
		19'b1101110010101101101: color_data = Z;
		19'b1101110010101101110: color_data = Z;
		19'b1101110010101101111: color_data = Z;
		19'b1101110010101110000: color_data = Z;
		19'b1101110010101110001: color_data = Z;
		19'b1101110010101110101: color_data = Z;
		19'b1101110010101110110: color_data = Z;
		19'b1101110010101110111: color_data = Z;
		19'b1101110100100011100: color_data = Z;
		19'b1101110100100100101: color_data = Z;
		19'b1101110100100100110: color_data = Z;
		19'b1101110100100100111: color_data = Z;
		19'b1101110100100101000: color_data = Z;
		19'b1101110100100101001: color_data = Z;
		19'b1101110100100101010: color_data = Z;
		19'b1101110100100101011: color_data = Z;
		19'b1101110100100101100: color_data = Z;
		19'b1101110100100101101: color_data = Z;
		19'b1101110100100101110: color_data = Z;
		19'b1101110100100101111: color_data = Z;
		19'b1101110100100110000: color_data = Z;
		19'b1101110100100110001: color_data = Z;
		19'b1101110100100110010: color_data = Z;
		19'b1101110100100110011: color_data = Z;
		19'b1101110100100110100: color_data = Z;
		19'b1101110100100110101: color_data = Z;
		19'b1101110100100110110: color_data = Z;
		19'b1101110100100110111: color_data = Z;
		19'b1101110100100111000: color_data = Z;
		19'b1101110100100111001: color_data = Z;
		19'b1101110100100111010: color_data = Z;
		19'b1101110100100111011: color_data = Z;
		19'b1101110100100111100: color_data = Z;
		19'b1101110100100111101: color_data = Z;
		19'b1101110100100111110: color_data = Z;
		19'b1101110100100111111: color_data = Z;
		19'b1101110100101000000: color_data = Z;
		19'b1101110100101000001: color_data = Z;
		19'b1101110100101000010: color_data = Z;
		19'b1101110100101000011: color_data = Z;
		19'b1101110100101000100: color_data = Z;
		19'b1101110100101000101: color_data = Z;
		19'b1101110100101000110: color_data = Z;
		19'b1101110100101000111: color_data = Z;
		19'b1101110100101001000: color_data = Z;
		19'b1101110100101001001: color_data = Z;
		19'b1101110100101001010: color_data = Z;
		19'b1101110100101001011: color_data = Z;
		19'b1101110100101001100: color_data = Z;
		19'b1101110100101001101: color_data = Z;
		19'b1101110100101001110: color_data = Z;
		19'b1101110100101001111: color_data = Z;
		19'b1101110100101010000: color_data = Z;
		19'b1101110100101010001: color_data = Z;
		19'b1101110100101010010: color_data = Z;
		19'b1101110100101010011: color_data = Z;
		19'b1101110100101010100: color_data = Z;
		19'b1101110100101010101: color_data = Z;
		19'b1101110100101010110: color_data = Z;
		19'b1101110100101010111: color_data = Z;
		19'b1101110100101011000: color_data = Z;
		19'b1101110100101011001: color_data = Z;
		19'b1101110100101011010: color_data = Z;
		19'b1101110100101011011: color_data = Z;
		19'b1101110100101011100: color_data = Z;
		19'b1101110100101011101: color_data = Z;
		19'b1101110100101011110: color_data = Z;
		19'b1101110100101011111: color_data = Z;
		19'b1101110100101100000: color_data = Z;
		19'b1101110100101100001: color_data = Z;
		19'b1101110100101100010: color_data = Z;
		19'b1101110100101100011: color_data = Z;
		19'b1101110100101100100: color_data = Z;
		19'b1101110100101100101: color_data = Z;
		19'b1101110100101100110: color_data = Z;
		19'b1101110100101100111: color_data = Z;
		19'b1101110100101101000: color_data = Z;
		19'b1101110100101101001: color_data = Z;
		19'b1101110100101101010: color_data = Z;
		19'b1101110100101101011: color_data = Z;
		19'b1101110100101101100: color_data = Z;
		19'b1101110100101101101: color_data = Z;
		19'b1101110100101101110: color_data = Z;
		19'b1101110100101101111: color_data = Z;
		19'b1101110100101110000: color_data = Z;
		19'b1101110100101110001: color_data = Z;
		19'b1101110100101110100: color_data = Z;
		19'b1101110100101110101: color_data = Z;
		19'b1101110100101110110: color_data = Z;
		19'b1101110100101110111: color_data = Z;
		19'b1101110110100011100: color_data = Z;
		19'b1101110110100100101: color_data = Z;
		19'b1101110110100100110: color_data = Z;
		19'b1101110110100100111: color_data = Z;
		19'b1101110110100101000: color_data = Z;
		19'b1101110110100101001: color_data = Z;
		19'b1101110110100101010: color_data = Z;
		19'b1101110110100101011: color_data = Z;
		19'b1101110110100101100: color_data = Z;
		19'b1101110110100101101: color_data = Z;
		19'b1101110110100101110: color_data = Z;
		19'b1101110110100101111: color_data = Z;
		19'b1101110110100110000: color_data = Z;
		19'b1101110110100110001: color_data = Z;
		19'b1101110110100110010: color_data = Z;
		19'b1101110110100110011: color_data = Z;
		19'b1101110110100110100: color_data = Z;
		19'b1101110110100110101: color_data = Z;
		19'b1101110110100110110: color_data = Z;
		19'b1101110110100110111: color_data = Z;
		19'b1101110110100111000: color_data = Z;
		19'b1101110110100111001: color_data = Z;
		19'b1101110110100111010: color_data = Z;
		19'b1101110110100111011: color_data = Z;
		19'b1101110110100111100: color_data = Z;
		19'b1101110110100111101: color_data = Z;
		19'b1101110110100111110: color_data = Z;
		19'b1101110110100111111: color_data = Z;
		19'b1101110110101000000: color_data = Z;
		19'b1101110110101000001: color_data = Z;
		19'b1101110110101000010: color_data = Z;
		19'b1101110110101000011: color_data = Z;
		19'b1101110110101000100: color_data = Z;
		19'b1101110110101000101: color_data = Z;
		19'b1101110110101000110: color_data = Z;
		19'b1101110110101000111: color_data = Z;
		19'b1101110110101001000: color_data = Z;
		19'b1101110110101001001: color_data = Z;
		19'b1101110110101001010: color_data = Z;
		19'b1101110110101001011: color_data = Z;
		19'b1101110110101001100: color_data = Z;
		19'b1101110110101001101: color_data = Z;
		19'b1101110110101001110: color_data = Z;
		19'b1101110110101001111: color_data = Z;
		19'b1101110110101010000: color_data = Z;
		19'b1101110110101010001: color_data = Z;
		19'b1101110110101010010: color_data = Z;
		19'b1101110110101010011: color_data = Z;
		19'b1101110110101010100: color_data = Z;
		19'b1101110110101010101: color_data = Z;
		19'b1101110110101010110: color_data = Z;
		19'b1101110110101010111: color_data = Z;
		19'b1101110110101011000: color_data = Z;
		19'b1101110110101011001: color_data = Z;
		19'b1101110110101011010: color_data = Z;
		19'b1101110110101011011: color_data = Z;
		19'b1101110110101011100: color_data = Z;
		19'b1101110110101011101: color_data = Z;
		19'b1101110110101011110: color_data = Z;
		19'b1101110110101011111: color_data = Z;
		19'b1101110110101100000: color_data = Z;
		19'b1101110110101100001: color_data = Z;
		19'b1101110110101100010: color_data = Z;
		19'b1101110110101100011: color_data = Z;
		19'b1101110110101100100: color_data = Z;
		19'b1101110110101100101: color_data = Z;
		19'b1101110110101100110: color_data = Z;
		19'b1101110110101100111: color_data = Z;
		19'b1101110110101101000: color_data = Z;
		19'b1101110110101101001: color_data = Z;
		19'b1101110110101101010: color_data = Z;
		19'b1101110110101101011: color_data = Z;
		19'b1101110110101101100: color_data = Z;
		19'b1101110110101101101: color_data = Z;
		19'b1101110110101101110: color_data = Z;
		19'b1101110110101101111: color_data = Z;
		19'b1101110110101110000: color_data = Z;
		19'b1101110110101110001: color_data = Z;
		19'b1101110110101110100: color_data = Z;
		19'b1101110110101110101: color_data = Z;
		19'b1101110110101110110: color_data = Z;
		19'b1101110110101110111: color_data = Z;
		19'b1101111000100100101: color_data = Z;
		19'b1101111000100100110: color_data = Z;
		19'b1101111000100100111: color_data = Z;
		19'b1101111000100101000: color_data = Z;
		19'b1101111000100101001: color_data = Z;
		19'b1101111000100101010: color_data = Z;
		19'b1101111000100101011: color_data = Z;
		19'b1101111000100101100: color_data = Z;
		19'b1101111000100101101: color_data = Z;
		19'b1101111000100101110: color_data = Z;
		19'b1101111000100101111: color_data = Z;
		19'b1101111000100110000: color_data = Z;
		19'b1101111000100110001: color_data = Z;
		19'b1101111000100110010: color_data = Z;
		19'b1101111000100110011: color_data = Z;
		19'b1101111000100110100: color_data = Z;
		19'b1101111000100110101: color_data = Z;
		19'b1101111000100110110: color_data = Z;
		19'b1101111000100110111: color_data = Z;
		19'b1101111000100111000: color_data = Z;
		19'b1101111000100111001: color_data = Z;
		19'b1101111000100111010: color_data = Z;
		19'b1101111000100111011: color_data = Z;
		19'b1101111000100111100: color_data = Z;
		19'b1101111000100111101: color_data = Z;
		19'b1101111000100111110: color_data = Z;
		19'b1101111000100111111: color_data = Z;
		19'b1101111000101000000: color_data = Z;
		19'b1101111000101000001: color_data = Z;
		19'b1101111000101000010: color_data = Z;
		19'b1101111000101000011: color_data = Z;
		19'b1101111000101000100: color_data = Z;
		19'b1101111000101000101: color_data = Z;
		19'b1101111000101000110: color_data = Z;
		19'b1101111000101000111: color_data = Z;
		19'b1101111000101001000: color_data = Z;
		19'b1101111000101001001: color_data = Z;
		19'b1101111000101001010: color_data = Z;
		19'b1101111000101001011: color_data = Z;
		19'b1101111000101001100: color_data = Z;
		19'b1101111000101001101: color_data = Z;
		19'b1101111000101001110: color_data = Z;
		19'b1101111000101001111: color_data = Z;
		19'b1101111000101010000: color_data = Z;
		19'b1101111000101010001: color_data = Z;
		19'b1101111000101010010: color_data = Z;
		19'b1101111000101010011: color_data = Z;
		19'b1101111000101010100: color_data = Z;
		19'b1101111000101010101: color_data = Z;
		19'b1101111000101010110: color_data = Z;
		19'b1101111000101010111: color_data = Z;
		19'b1101111000101011000: color_data = Z;
		19'b1101111000101011001: color_data = Z;
		19'b1101111000101011010: color_data = Z;
		19'b1101111000101011011: color_data = Z;
		19'b1101111000101011100: color_data = Z;
		19'b1101111000101011101: color_data = Z;
		19'b1101111000101011110: color_data = Z;
		19'b1101111000101011111: color_data = Z;
		19'b1101111000101100000: color_data = Z;
		19'b1101111000101100001: color_data = Z;
		19'b1101111000101100010: color_data = Z;
		19'b1101111000101100011: color_data = Z;
		19'b1101111000101100100: color_data = Z;
		19'b1101111000101100101: color_data = Z;
		19'b1101111000101100110: color_data = Z;
		19'b1101111000101100111: color_data = Z;
		19'b1101111000101101000: color_data = Z;
		19'b1101111000101101001: color_data = Z;
		19'b1101111000101101010: color_data = Z;
		19'b1101111000101101011: color_data = Z;
		19'b1101111000101101100: color_data = Z;
		19'b1101111000101101101: color_data = Z;
		19'b1101111000101101110: color_data = Z;
		19'b1101111000101101111: color_data = Z;
		19'b1101111000101110000: color_data = Z;
		19'b1101111000101110100: color_data = Z;
		19'b1101111000101110101: color_data = Z;
		19'b1101111000101110110: color_data = Z;
		19'b1101111000101110111: color_data = Z;
		19'b1101111010100100101: color_data = Z;
		19'b1101111010100100110: color_data = Z;
		19'b1101111010100100111: color_data = Z;
		19'b1101111010100101000: color_data = Z;
		19'b1101111010100101001: color_data = Z;
		19'b1101111010100101010: color_data = Z;
		19'b1101111010100101011: color_data = Z;
		19'b1101111010100101100: color_data = Z;
		19'b1101111010100101101: color_data = Z;
		19'b1101111010100101110: color_data = Z;
		19'b1101111010100101111: color_data = Z;
		19'b1101111010100110000: color_data = Z;
		19'b1101111010100110001: color_data = Z;
		19'b1101111010100110010: color_data = Z;
		19'b1101111010100110011: color_data = Z;
		19'b1101111010100110100: color_data = Z;
		19'b1101111010100110101: color_data = Z;
		19'b1101111010100110110: color_data = Z;
		19'b1101111010100110111: color_data = Z;
		19'b1101111010100111000: color_data = Z;
		19'b1101111010100111001: color_data = Z;
		19'b1101111010100111010: color_data = Z;
		19'b1101111010100111011: color_data = Z;
		19'b1101111010100111100: color_data = Z;
		19'b1101111010100111101: color_data = Z;
		19'b1101111010100111110: color_data = Z;
		19'b1101111010100111111: color_data = Z;
		19'b1101111010101000000: color_data = Z;
		19'b1101111010101000001: color_data = Z;
		19'b1101111010101000010: color_data = Z;
		19'b1101111010101000011: color_data = Z;
		19'b1101111010101000100: color_data = Z;
		19'b1101111010101000101: color_data = Z;
		19'b1101111010101000110: color_data = Z;
		19'b1101111010101000111: color_data = Z;
		19'b1101111010101001000: color_data = Z;
		19'b1101111010101001001: color_data = Z;
		19'b1101111010101001010: color_data = Z;
		19'b1101111010101001011: color_data = Z;
		19'b1101111010101001100: color_data = Z;
		19'b1101111010101001101: color_data = Z;
		19'b1101111010101001110: color_data = Z;
		19'b1101111010101001111: color_data = Z;
		19'b1101111010101010000: color_data = Z;
		19'b1101111010101010001: color_data = Z;
		19'b1101111010101010010: color_data = Z;
		19'b1101111010101010011: color_data = Z;
		19'b1101111010101010100: color_data = Z;
		19'b1101111010101010101: color_data = Z;
		19'b1101111010101010110: color_data = Z;
		19'b1101111010101010111: color_data = Z;
		19'b1101111010101011000: color_data = Z;
		19'b1101111010101011001: color_data = Z;
		19'b1101111010101011010: color_data = Z;
		19'b1101111010101011011: color_data = Z;
		19'b1101111010101011100: color_data = Z;
		19'b1101111010101011101: color_data = Z;
		19'b1101111010101011110: color_data = Z;
		19'b1101111010101011111: color_data = Z;
		19'b1101111010101100000: color_data = Z;
		19'b1101111010101100001: color_data = Z;
		19'b1101111010101100010: color_data = Z;
		19'b1101111010101100011: color_data = Z;
		19'b1101111010101100100: color_data = Z;
		19'b1101111010101100101: color_data = Z;
		19'b1101111010101100110: color_data = Z;
		19'b1101111010101100111: color_data = Z;
		19'b1101111010101101000: color_data = Z;
		19'b1101111010101101001: color_data = Z;
		19'b1101111010101101010: color_data = Z;
		19'b1101111010101101011: color_data = Z;
		19'b1101111010101101100: color_data = Z;
		19'b1101111010101101101: color_data = Z;
		19'b1101111010101101110: color_data = Z;
		19'b1101111010101101111: color_data = Z;
		19'b1101111010101110000: color_data = Z;
		19'b1101111010101110010: color_data = Z;
		19'b1101111010101110011: color_data = Z;
		19'b1101111010101110100: color_data = Z;
		19'b1101111010101110101: color_data = Z;
		19'b1101111010101110110: color_data = Z;
		19'b1101111010101110111: color_data = Z;
		19'b1101111100100100110: color_data = Z;
		19'b1101111100100100111: color_data = Z;
		19'b1101111100100101000: color_data = Z;
		19'b1101111100100101001: color_data = Z;
		19'b1101111100100101010: color_data = Z;
		19'b1101111100100101011: color_data = Z;
		19'b1101111100100101100: color_data = Z;
		19'b1101111100100101101: color_data = Z;
		19'b1101111100100101110: color_data = Z;
		19'b1101111100100101111: color_data = Z;
		19'b1101111100100110000: color_data = Z;
		19'b1101111100100110001: color_data = Z;
		19'b1101111100100110010: color_data = Z;
		19'b1101111100100110011: color_data = Z;
		19'b1101111100100110100: color_data = Z;
		19'b1101111100100110101: color_data = Z;
		19'b1101111100100110110: color_data = Z;
		19'b1101111100100110111: color_data = Z;
		19'b1101111100100111000: color_data = Z;
		19'b1101111100100111001: color_data = Z;
		19'b1101111100100111010: color_data = Z;
		19'b1101111100100111011: color_data = Z;
		19'b1101111100100111100: color_data = Z;
		19'b1101111100100111101: color_data = Z;
		19'b1101111100100111110: color_data = Z;
		19'b1101111100100111111: color_data = Z;
		19'b1101111100101000000: color_data = Z;
		19'b1101111100101000001: color_data = Z;
		19'b1101111100101000010: color_data = Z;
		19'b1101111100101000011: color_data = Z;
		19'b1101111100101000100: color_data = Z;
		19'b1101111100101000101: color_data = Z;
		19'b1101111100101000110: color_data = Z;
		19'b1101111100101000111: color_data = Z;
		19'b1101111100101001000: color_data = Z;
		19'b1101111100101001001: color_data = Z;
		19'b1101111100101001010: color_data = Z;
		19'b1101111100101001011: color_data = Z;
		19'b1101111100101001100: color_data = Z;
		19'b1101111100101001101: color_data = Z;
		19'b1101111100101001110: color_data = Z;
		19'b1101111100101001111: color_data = Z;
		19'b1101111100101010000: color_data = Z;
		19'b1101111100101010001: color_data = Z;
		19'b1101111100101010010: color_data = Z;
		19'b1101111100101010011: color_data = Z;
		19'b1101111100101010100: color_data = Z;
		19'b1101111100101010101: color_data = Z;
		19'b1101111100101010110: color_data = Z;
		19'b1101111100101010111: color_data = Z;
		19'b1101111100101011000: color_data = Z;
		19'b1101111100101011001: color_data = Z;
		19'b1101111100101011010: color_data = Z;
		19'b1101111100101011011: color_data = Z;
		19'b1101111100101011100: color_data = Z;
		19'b1101111100101011101: color_data = Z;
		19'b1101111100101011110: color_data = Z;
		19'b1101111100101011111: color_data = Z;
		19'b1101111100101100000: color_data = Z;
		19'b1101111100101100001: color_data = Z;
		19'b1101111100101100010: color_data = Z;
		19'b1101111100101100011: color_data = Z;
		19'b1101111100101100100: color_data = Z;
		19'b1101111100101100101: color_data = Z;
		19'b1101111100101100110: color_data = Z;
		19'b1101111100101100111: color_data = Z;
		19'b1101111100101101000: color_data = Z;
		19'b1101111100101101001: color_data = Z;
		19'b1101111100101101010: color_data = Z;
		19'b1101111100101101011: color_data = Z;
		19'b1101111100101101100: color_data = Z;
		19'b1101111100101101101: color_data = Z;
		19'b1101111100101101110: color_data = Z;
		19'b1101111100101101111: color_data = Z;
		19'b1101111100101110000: color_data = Z;
		19'b1101111100101110001: color_data = Z;
		19'b1101111100101110010: color_data = Z;
		19'b1101111100101110011: color_data = Z;
		19'b1101111100101110100: color_data = Z;
		19'b1101111100101110101: color_data = Z;
		19'b1101111100101110110: color_data = Z;
		19'b1101111100101110111: color_data = Z;
		19'b1101111110100100110: color_data = Z;
		19'b1101111110100100111: color_data = Z;
		19'b1101111110100101000: color_data = Z;
		19'b1101111110100101001: color_data = Z;
		19'b1101111110100101010: color_data = Z;
		19'b1101111110100101011: color_data = Z;
		19'b1101111110100101100: color_data = Z;
		19'b1101111110100101101: color_data = Z;
		19'b1101111110100101110: color_data = Z;
		19'b1101111110100101111: color_data = Z;
		19'b1101111110100110000: color_data = Z;
		19'b1101111110100110001: color_data = Z;
		19'b1101111110100110010: color_data = Z;
		19'b1101111110100110011: color_data = Z;
		19'b1101111110100110100: color_data = Z;
		19'b1101111110100110101: color_data = Z;
		19'b1101111110100110110: color_data = Z;
		19'b1101111110100110111: color_data = Z;
		19'b1101111110100111000: color_data = Z;
		19'b1101111110100111001: color_data = Z;
		19'b1101111110100111010: color_data = Z;
		19'b1101111110100111011: color_data = Z;
		19'b1101111110100111100: color_data = Z;
		19'b1101111110100111101: color_data = Z;
		19'b1101111110100111110: color_data = Z;
		19'b1101111110100111111: color_data = Z;
		19'b1101111110101000000: color_data = Z;
		19'b1101111110101000001: color_data = Z;
		19'b1101111110101000010: color_data = Z;
		19'b1101111110101000011: color_data = Z;
		19'b1101111110101000100: color_data = Z;
		19'b1101111110101000101: color_data = Z;
		19'b1101111110101000110: color_data = Z;
		19'b1101111110101000111: color_data = Z;
		19'b1101111110101001000: color_data = Z;
		19'b1101111110101001001: color_data = Z;
		19'b1101111110101001010: color_data = Z;
		19'b1101111110101001011: color_data = Z;
		19'b1101111110101001100: color_data = Z;
		19'b1101111110101001101: color_data = Z;
		19'b1101111110101001110: color_data = Z;
		19'b1101111110101001111: color_data = Z;
		19'b1101111110101010000: color_data = Z;
		19'b1101111110101010001: color_data = Z;
		19'b1101111110101010010: color_data = Z;
		19'b1101111110101010011: color_data = Z;
		19'b1101111110101010100: color_data = Z;
		19'b1101111110101010101: color_data = Z;
		19'b1101111110101010110: color_data = Z;
		19'b1101111110101010111: color_data = Z;
		19'b1101111110101011000: color_data = Z;
		19'b1101111110101011001: color_data = Z;
		19'b1101111110101011010: color_data = Z;
		19'b1101111110101011011: color_data = Z;
		19'b1101111110101011100: color_data = Z;
		19'b1101111110101011101: color_data = Z;
		19'b1101111110101011110: color_data = Z;
		19'b1101111110101011111: color_data = Z;
		19'b1101111110101100000: color_data = Z;
		19'b1101111110101100001: color_data = Z;
		19'b1101111110101100010: color_data = Z;
		19'b1101111110101100011: color_data = Z;
		19'b1101111110101100100: color_data = Z;
		19'b1101111110101100101: color_data = Z;
		19'b1101111110101100110: color_data = Z;
		19'b1101111110101100111: color_data = Z;
		19'b1101111110101101000: color_data = Z;
		19'b1101111110101101001: color_data = Z;
		19'b1101111110101101010: color_data = Z;
		19'b1101111110101101011: color_data = Z;
		19'b1101111110101101100: color_data = Z;
		19'b1101111110101101101: color_data = Z;
		19'b1101111110101101110: color_data = Z;
		19'b1101111110101101111: color_data = Z;
		19'b1101111110101110000: color_data = Z;
		19'b1101111110101110001: color_data = Z;
		19'b1101111110101110010: color_data = Z;
		19'b1101111110101110011: color_data = Z;
		19'b1101111110101110100: color_data = Z;
		19'b1101111110101110101: color_data = Z;
		19'b1101111110101110110: color_data = Z;
		19'b1101111110101110111: color_data = Z;
		19'b1110000000100100110: color_data = Z;
		19'b1110000000100100111: color_data = Z;
		19'b1110000000100101000: color_data = Z;
		19'b1110000000100101001: color_data = Z;
		19'b1110000000100101010: color_data = Z;
		19'b1110000000100101011: color_data = Z;
		19'b1110000000100101100: color_data = Z;
		19'b1110000000100101101: color_data = Z;
		19'b1110000000100101110: color_data = Z;
		19'b1110000000100101111: color_data = Z;
		19'b1110000000100110000: color_data = Z;
		19'b1110000000100110001: color_data = Z;
		19'b1110000000100110010: color_data = Z;
		19'b1110000000100110011: color_data = Z;
		19'b1110000000100110100: color_data = Z;
		19'b1110000000100110101: color_data = Z;
		19'b1110000000100110110: color_data = Z;
		19'b1110000000100110111: color_data = Z;
		19'b1110000000100111000: color_data = Z;
		19'b1110000000100111001: color_data = Z;
		19'b1110000000100111010: color_data = Z;
		19'b1110000000100111011: color_data = Z;
		19'b1110000000100111100: color_data = Z;
		19'b1110000000100111101: color_data = Z;
		19'b1110000000100111110: color_data = Z;
		19'b1110000000100111111: color_data = Z;
		19'b1110000000101000000: color_data = Z;
		19'b1110000000101000001: color_data = Z;
		19'b1110000000101000010: color_data = Z;
		19'b1110000000101000011: color_data = Z;
		19'b1110000000101000100: color_data = Z;
		19'b1110000000101000101: color_data = Z;
		19'b1110000000101000110: color_data = Z;
		19'b1110000000101000111: color_data = Z;
		19'b1110000000101001000: color_data = Z;
		19'b1110000000101001001: color_data = Z;
		19'b1110000000101001010: color_data = Z;
		19'b1110000000101001011: color_data = Z;
		19'b1110000000101001100: color_data = Z;
		19'b1110000000101001101: color_data = Z;
		19'b1110000000101001110: color_data = Z;
		19'b1110000000101001111: color_data = Z;
		19'b1110000000101010000: color_data = Z;
		19'b1110000000101010001: color_data = Z;
		19'b1110000000101010010: color_data = Z;
		19'b1110000000101010011: color_data = Z;
		19'b1110000000101010100: color_data = Z;
		19'b1110000000101010101: color_data = Z;
		19'b1110000000101010110: color_data = Z;
		19'b1110000000101010111: color_data = Z;
		19'b1110000000101011000: color_data = Z;
		19'b1110000000101011001: color_data = Z;
		19'b1110000000101011010: color_data = Z;
		19'b1110000000101011011: color_data = Z;
		19'b1110000000101011100: color_data = Z;
		19'b1110000000101011101: color_data = Z;
		19'b1110000000101011110: color_data = Z;
		19'b1110000000101011111: color_data = Z;
		19'b1110000000101100000: color_data = Z;
		19'b1110000000101100001: color_data = Z;
		19'b1110000000101100010: color_data = Z;
		19'b1110000000101100011: color_data = Z;
		19'b1110000000101100100: color_data = Z;
		19'b1110000000101100101: color_data = Z;
		19'b1110000000101100110: color_data = Z;
		19'b1110000000101100111: color_data = Z;
		19'b1110000000101101000: color_data = Z;
		19'b1110000000101101001: color_data = Z;
		19'b1110000000101101010: color_data = Z;
		19'b1110000000101101011: color_data = Z;
		19'b1110000000101101100: color_data = Z;
		19'b1110000000101101101: color_data = Z;
		19'b1110000000101101110: color_data = Z;
		19'b1110000000101101111: color_data = Z;
		19'b1110000000101110000: color_data = Z;
		19'b1110000000101110001: color_data = Z;
		19'b1110000000101110010: color_data = Z;
		19'b1110000000101110011: color_data = Z;
		19'b1110000000101110100: color_data = Z;
		19'b1110000000101110101: color_data = Z;
		19'b1110000000101110110: color_data = Z;
		19'b1110000000101110111: color_data = Z;
		19'b1110000010100100110: color_data = Z;
		19'b1110000010100100111: color_data = Z;
		19'b1110000010100101000: color_data = Z;
		19'b1110000010100101001: color_data = Z;
		19'b1110000010100101010: color_data = Z;
		19'b1110000010100101011: color_data = Z;
		19'b1110000010100101100: color_data = Z;
		19'b1110000010100101101: color_data = Z;
		19'b1110000010100101110: color_data = Z;
		19'b1110000010100101111: color_data = Z;
		19'b1110000010100110000: color_data = Z;
		19'b1110000010100110001: color_data = Z;
		19'b1110000010100110010: color_data = Z;
		19'b1110000010100110011: color_data = Z;
		19'b1110000010100110100: color_data = Z;
		19'b1110000010100110101: color_data = Z;
		19'b1110000010100110110: color_data = Z;
		19'b1110000010100110111: color_data = Z;
		19'b1110000010100111000: color_data = Z;
		19'b1110000010100111001: color_data = Z;
		19'b1110000010100111010: color_data = Z;
		19'b1110000010100111011: color_data = Z;
		19'b1110000010100111100: color_data = Z;
		19'b1110000010100111101: color_data = Z;
		19'b1110000010100111110: color_data = Z;
		19'b1110000010100111111: color_data = Z;
		19'b1110000010101000000: color_data = Z;
		19'b1110000010101000001: color_data = Z;
		19'b1110000010101000010: color_data = Z;
		19'b1110000010101000011: color_data = Z;
		19'b1110000010101000100: color_data = Z;
		19'b1110000010101000101: color_data = Z;
		19'b1110000010101000110: color_data = Z;
		19'b1110000010101000111: color_data = Z;
		19'b1110000010101001000: color_data = Z;
		19'b1110000010101001001: color_data = Z;
		19'b1110000010101001010: color_data = Z;
		19'b1110000010101001011: color_data = Z;
		19'b1110000010101001100: color_data = Z;
		19'b1110000010101001101: color_data = Z;
		19'b1110000010101001110: color_data = Z;
		19'b1110000010101001111: color_data = Z;
		19'b1110000010101010000: color_data = Z;
		19'b1110000010101010001: color_data = Z;
		19'b1110000010101010010: color_data = Z;
		19'b1110000010101010011: color_data = Z;
		19'b1110000010101010100: color_data = Z;
		19'b1110000010101010101: color_data = Z;
		19'b1110000010101010110: color_data = Z;
		19'b1110000010101010111: color_data = Z;
		19'b1110000010101011000: color_data = Z;
		19'b1110000010101011001: color_data = Z;
		19'b1110000010101011010: color_data = Z;
		19'b1110000010101011011: color_data = Z;
		19'b1110000010101011100: color_data = Z;
		19'b1110000010101011101: color_data = Z;
		19'b1110000010101011110: color_data = Z;
		19'b1110000010101011111: color_data = Z;
		19'b1110000010101100000: color_data = Z;
		19'b1110000010101100001: color_data = Z;
		19'b1110000010101100010: color_data = Z;
		19'b1110000010101100011: color_data = Z;
		19'b1110000010101100100: color_data = Z;
		19'b1110000010101100101: color_data = Z;
		19'b1110000010101100110: color_data = Z;
		19'b1110000010101100111: color_data = Z;
		19'b1110000010101101000: color_data = Z;
		19'b1110000010101101001: color_data = Z;
		19'b1110000010101101010: color_data = Z;
		19'b1110000010101101011: color_data = Z;
		19'b1110000010101101100: color_data = Z;
		19'b1110000010101101101: color_data = Z;
		19'b1110000010101101110: color_data = Z;
		19'b1110000010101101111: color_data = Z;
		19'b1110000010101110000: color_data = Z;
		19'b1110000010101110001: color_data = Z;
		19'b1110000010101110010: color_data = Z;
		19'b1110000010101110011: color_data = Z;
		19'b1110000010101110100: color_data = Z;
		19'b1110000010101110101: color_data = Z;
		19'b1110000010101110110: color_data = Z;
		19'b1110000010101110111: color_data = Z;
		19'b1110000100100100110: color_data = Z;
		19'b1110000100100100111: color_data = Z;
		19'b1110000100100101000: color_data = Z;
		19'b1110000100100101001: color_data = Z;
		19'b1110000100100101010: color_data = Z;
		19'b1110000100100101011: color_data = Z;
		19'b1110000100100101100: color_data = Z;
		19'b1110000100100101101: color_data = Z;
		19'b1110000100100101110: color_data = Z;
		19'b1110000100100101111: color_data = Z;
		19'b1110000100100110000: color_data = Z;
		19'b1110000100100110001: color_data = Z;
		19'b1110000100100110010: color_data = Z;
		19'b1110000100100110011: color_data = Z;
		19'b1110000100100110100: color_data = Z;
		19'b1110000100100110101: color_data = Z;
		19'b1110000100100110110: color_data = Z;
		19'b1110000100100110111: color_data = Z;
		19'b1110000100100111000: color_data = Z;
		19'b1110000100100111001: color_data = Z;
		19'b1110000100100111010: color_data = Z;
		19'b1110000100100111011: color_data = Z;
		19'b1110000100100111100: color_data = Z;
		19'b1110000100100111101: color_data = Z;
		19'b1110000100100111110: color_data = Z;
		19'b1110000100100111111: color_data = Z;
		19'b1110000100101000000: color_data = Z;
		19'b1110000100101000001: color_data = Z;
		19'b1110000100101000010: color_data = Z;
		19'b1110000100101000011: color_data = Z;
		19'b1110000100101000100: color_data = Z;
		19'b1110000100101000101: color_data = Z;
		19'b1110000100101000110: color_data = Z;
		19'b1110000100101000111: color_data = Z;
		19'b1110000100101001000: color_data = Z;
		19'b1110000100101001001: color_data = Z;
		19'b1110000100101001010: color_data = Z;
		19'b1110000100101001011: color_data = Z;
		19'b1110000100101001100: color_data = Z;
		19'b1110000100101001101: color_data = Z;
		19'b1110000100101001110: color_data = Z;
		19'b1110000100101001111: color_data = Z;
		19'b1110000100101010000: color_data = Z;
		19'b1110000100101010001: color_data = Z;
		19'b1110000100101010010: color_data = Z;
		19'b1110000100101010011: color_data = Z;
		19'b1110000100101010100: color_data = Z;
		19'b1110000100101010101: color_data = Z;
		19'b1110000100101010110: color_data = Z;
		19'b1110000100101010111: color_data = Z;
		19'b1110000100101011000: color_data = Z;
		19'b1110000100101011001: color_data = Z;
		19'b1110000100101011010: color_data = Z;
		19'b1110000100101011011: color_data = Z;
		19'b1110000100101011100: color_data = Z;
		19'b1110000100101011101: color_data = Z;
		19'b1110000100101011110: color_data = Z;
		19'b1110000100101011111: color_data = Z;
		19'b1110000100101100000: color_data = Z;
		19'b1110000100101100001: color_data = Z;
		19'b1110000100101100010: color_data = Z;
		19'b1110000100101100011: color_data = Z;
		19'b1110000100101100100: color_data = Z;
		19'b1110000100101100101: color_data = Z;
		19'b1110000100101100110: color_data = Z;
		19'b1110000100101100111: color_data = Z;
		19'b1110000100101101000: color_data = Z;
		19'b1110000100101101001: color_data = Z;
		19'b1110000100101101010: color_data = Z;
		19'b1110000100101101011: color_data = Z;
		19'b1110000100101101100: color_data = Z;
		19'b1110000100101101101: color_data = Z;
		19'b1110000100101101110: color_data = Z;
		19'b1110000100101101111: color_data = Z;
		19'b1110000100101110000: color_data = Z;
		19'b1110000100101110001: color_data = Z;
		19'b1110000100101110010: color_data = Z;
		19'b1110000100101110011: color_data = Z;
		19'b1110000100101110100: color_data = Z;
		19'b1110000100101110101: color_data = Z;
		19'b1110000100101110110: color_data = Z;
		19'b1110000100101110111: color_data = Z;
		19'b1110000110100100110: color_data = Z;
		19'b1110000110100100111: color_data = Z;
		19'b1110000110100101000: color_data = Z;
		19'b1110000110100101001: color_data = Z;
		19'b1110000110100101010: color_data = Z;
		19'b1110000110100101011: color_data = Z;
		19'b1110000110100101100: color_data = Z;
		19'b1110000110100101101: color_data = Z;
		19'b1110000110100101110: color_data = Z;
		19'b1110000110100101111: color_data = Z;
		19'b1110000110100110000: color_data = Z;
		19'b1110000110100110001: color_data = Z;
		19'b1110000110100110010: color_data = Z;
		19'b1110000110100110011: color_data = Z;
		19'b1110000110100110100: color_data = Z;
		19'b1110000110100110101: color_data = Z;
		19'b1110000110100110110: color_data = Z;
		19'b1110000110100110111: color_data = Z;
		19'b1110000110100111000: color_data = Z;
		19'b1110000110100111001: color_data = Z;
		19'b1110000110100111010: color_data = Z;
		19'b1110000110100111011: color_data = Z;
		19'b1110000110100111100: color_data = Z;
		19'b1110000110100111101: color_data = Z;
		19'b1110000110100111110: color_data = Z;
		19'b1110000110100111111: color_data = Z;
		19'b1110000110101000000: color_data = Z;
		19'b1110000110101000001: color_data = Z;
		19'b1110000110101000010: color_data = Z;
		19'b1110000110101000011: color_data = Z;
		19'b1110000110101000100: color_data = Z;
		19'b1110000110101000101: color_data = Z;
		19'b1110000110101000110: color_data = Z;
		19'b1110000110101000111: color_data = Z;
		19'b1110000110101001000: color_data = Z;
		19'b1110000110101001001: color_data = Z;
		19'b1110000110101001010: color_data = Z;
		19'b1110000110101001011: color_data = Z;
		19'b1110000110101001100: color_data = Z;
		19'b1110000110101001101: color_data = Z;
		19'b1110000110101001110: color_data = Z;
		19'b1110000110101001111: color_data = Z;
		19'b1110000110101010000: color_data = Z;
		19'b1110000110101010001: color_data = Z;
		19'b1110000110101010010: color_data = Z;
		19'b1110000110101010011: color_data = Z;
		19'b1110000110101010100: color_data = Z;
		19'b1110000110101010101: color_data = Z;
		19'b1110000110101010110: color_data = Z;
		19'b1110000110101010111: color_data = Z;
		19'b1110000110101011000: color_data = Z;
		19'b1110000110101011001: color_data = Z;
		19'b1110000110101011010: color_data = Z;
		19'b1110000110101011011: color_data = Z;
		19'b1110000110101011100: color_data = Z;
		19'b1110000110101011101: color_data = Z;
		19'b1110000110101011110: color_data = Z;
		19'b1110000110101011111: color_data = Z;
		19'b1110000110101100000: color_data = Z;
		19'b1110000110101100001: color_data = Z;
		19'b1110000110101100010: color_data = Z;
		19'b1110000110101100011: color_data = Z;
		19'b1110000110101100100: color_data = Z;
		19'b1110000110101100101: color_data = Z;
		19'b1110000110101100110: color_data = Z;
		19'b1110000110101100111: color_data = Z;
		19'b1110000110101101000: color_data = Z;
		19'b1110000110101101001: color_data = Z;
		19'b1110000110101101010: color_data = Z;
		19'b1110000110101101011: color_data = Z;
		19'b1110000110101101100: color_data = Z;
		19'b1110000110101101101: color_data = Z;
		19'b1110000110101101110: color_data = Z;
		19'b1110000110101101111: color_data = Z;
		19'b1110000110101110000: color_data = Z;
		19'b1110000110101110001: color_data = Z;
		19'b1110000110101110010: color_data = Z;
		19'b1110000110101110011: color_data = Z;
		19'b1110000110101110100: color_data = Z;
		19'b1110000110101110101: color_data = Z;
		19'b1110000110101110110: color_data = Z;
		19'b1110000110101110111: color_data = Z;
		19'b1110001000100011111: color_data = Z;
		19'b1110001000100100110: color_data = Z;
		19'b1110001000100100111: color_data = Z;
		19'b1110001000100101000: color_data = Z;
		19'b1110001000100101001: color_data = Z;
		19'b1110001000100101010: color_data = Z;
		19'b1110001000100101011: color_data = Z;
		19'b1110001000100101100: color_data = Z;
		19'b1110001000100101101: color_data = Z;
		19'b1110001000100101110: color_data = Z;
		19'b1110001000100101111: color_data = Z;
		19'b1110001000100110000: color_data = Z;
		19'b1110001000100110001: color_data = Z;
		19'b1110001000100110010: color_data = Z;
		19'b1110001000100110011: color_data = Z;
		19'b1110001000100110100: color_data = Z;
		19'b1110001000100110101: color_data = Z;
		19'b1110001000100110110: color_data = Z;
		19'b1110001000100110111: color_data = Z;
		19'b1110001000100111000: color_data = Z;
		19'b1110001000100111001: color_data = Z;
		19'b1110001000100111010: color_data = Z;
		19'b1110001000100111011: color_data = Z;
		19'b1110001000100111100: color_data = Z;
		19'b1110001000100111101: color_data = Z;
		19'b1110001000100111110: color_data = Z;
		19'b1110001000100111111: color_data = Z;
		19'b1110001000101000000: color_data = Z;
		19'b1110001000101000001: color_data = Z;
		19'b1110001000101000010: color_data = Z;
		19'b1110001000101000011: color_data = Z;
		19'b1110001000101000100: color_data = Z;
		19'b1110001000101000101: color_data = Z;
		19'b1110001000101000110: color_data = Z;
		19'b1110001000101000111: color_data = Z;
		19'b1110001000101001000: color_data = Z;
		19'b1110001000101001001: color_data = Z;
		19'b1110001000101001010: color_data = Z;
		19'b1110001000101001011: color_data = Z;
		19'b1110001000101001100: color_data = Z;
		19'b1110001000101001101: color_data = Z;
		19'b1110001000101001110: color_data = Z;
		19'b1110001000101001111: color_data = Z;
		19'b1110001000101010000: color_data = Z;
		19'b1110001000101010001: color_data = Z;
		19'b1110001000101010010: color_data = Z;
		19'b1110001000101010011: color_data = Z;
		19'b1110001000101010100: color_data = Z;
		19'b1110001000101010101: color_data = Z;
		19'b1110001000101010110: color_data = Z;
		19'b1110001000101010111: color_data = Z;
		19'b1110001000101011000: color_data = Z;
		19'b1110001000101011001: color_data = Z;
		19'b1110001000101011010: color_data = Z;
		19'b1110001000101011011: color_data = Z;
		19'b1110001000101011100: color_data = Z;
		19'b1110001000101011101: color_data = Z;
		19'b1110001000101011110: color_data = Z;
		19'b1110001000101011111: color_data = Z;
		19'b1110001000101100000: color_data = Z;
		19'b1110001000101100001: color_data = Z;
		19'b1110001000101100010: color_data = Z;
		19'b1110001000101100011: color_data = Z;
		19'b1110001000101100100: color_data = Z;
		19'b1110001000101100101: color_data = Z;
		19'b1110001000101100110: color_data = Z;
		19'b1110001000101100111: color_data = Z;
		19'b1110001000101101000: color_data = Z;
		19'b1110001000101101001: color_data = Z;
		19'b1110001000101101010: color_data = Z;
		19'b1110001000101101011: color_data = Z;
		19'b1110001000101101100: color_data = Z;
		19'b1110001000101101101: color_data = Z;
		19'b1110001000101101110: color_data = Z;
		19'b1110001000101101111: color_data = Z;
		19'b1110001000101110000: color_data = Z;
		19'b1110001000101110001: color_data = Z;
		19'b1110001000101110010: color_data = Z;
		19'b1110001000101110011: color_data = Z;
		19'b1110001000101110100: color_data = Z;
		19'b1110001000101110101: color_data = Z;
		19'b1110001000101110110: color_data = Z;
		19'b1110001010100011111: color_data = Z;
		19'b1110001010100100110: color_data = Z;
		19'b1110001010100100111: color_data = Z;
		19'b1110001010100101000: color_data = Z;
		19'b1110001010100101001: color_data = Z;
		19'b1110001010100101010: color_data = Z;
		19'b1110001010100101011: color_data = Z;
		19'b1110001010100101100: color_data = Z;
		19'b1110001010100101101: color_data = Z;
		19'b1110001010100101110: color_data = Z;
		19'b1110001010100101111: color_data = Z;
		19'b1110001010100110000: color_data = Z;
		19'b1110001010100110001: color_data = Z;
		19'b1110001010100110010: color_data = Z;
		19'b1110001010100110011: color_data = Z;
		19'b1110001010100110100: color_data = Z;
		19'b1110001010100110101: color_data = Z;
		19'b1110001010100110110: color_data = Z;
		19'b1110001010100110111: color_data = Z;
		19'b1110001010100111000: color_data = Z;
		19'b1110001010100111001: color_data = Z;
		19'b1110001010100111010: color_data = Z;
		19'b1110001010100111011: color_data = Z;
		19'b1110001010100111100: color_data = Z;
		19'b1110001010100111101: color_data = Z;
		19'b1110001010100111110: color_data = Z;
		19'b1110001010100111111: color_data = Z;
		19'b1110001010101000000: color_data = Z;
		19'b1110001010101000001: color_data = Z;
		19'b1110001010101000010: color_data = Z;
		19'b1110001010101000011: color_data = Z;
		19'b1110001010101000100: color_data = Z;
		19'b1110001010101000101: color_data = Z;
		19'b1110001010101000110: color_data = Z;
		19'b1110001010101000111: color_data = Z;
		19'b1110001010101001000: color_data = Z;
		19'b1110001010101001001: color_data = Z;
		19'b1110001010101001010: color_data = Z;
		19'b1110001010101001011: color_data = Z;
		19'b1110001010101001100: color_data = Z;
		19'b1110001010101001101: color_data = Z;
		19'b1110001010101001110: color_data = Z;
		19'b1110001010101001111: color_data = Z;
		19'b1110001010101010000: color_data = Z;
		19'b1110001010101010001: color_data = Z;
		19'b1110001010101010010: color_data = Z;
		19'b1110001010101010011: color_data = Z;
		19'b1110001010101010100: color_data = Z;
		19'b1110001010101010101: color_data = Z;
		19'b1110001010101010110: color_data = Z;
		19'b1110001010101010111: color_data = Z;
		19'b1110001010101011000: color_data = Z;
		19'b1110001010101011001: color_data = Z;
		19'b1110001010101011010: color_data = Z;
		19'b1110001010101011011: color_data = Z;
		19'b1110001010101011100: color_data = Z;
		19'b1110001010101011101: color_data = Z;
		19'b1110001010101011110: color_data = Z;
		19'b1110001010101011111: color_data = Z;
		19'b1110001010101100000: color_data = Z;
		19'b1110001010101100001: color_data = Z;
		19'b1110001010101100010: color_data = Z;
		19'b1110001010101100011: color_data = Z;
		19'b1110001010101100100: color_data = Z;
		19'b1110001010101100101: color_data = Z;
		19'b1110001010101100110: color_data = Z;
		19'b1110001010101100111: color_data = Z;
		19'b1110001010101101000: color_data = Z;
		19'b1110001010101101001: color_data = Z;
		19'b1110001010101101010: color_data = Z;
		19'b1110001010101101011: color_data = Z;
		19'b1110001010101101100: color_data = Z;
		19'b1110001010101101101: color_data = Z;
		19'b1110001010101101110: color_data = Z;
		19'b1110001010101101111: color_data = Z;
		19'b1110001010101110000: color_data = Z;
		19'b1110001010101110001: color_data = Z;
		19'b1110001010101110010: color_data = Z;
		19'b1110001010101110011: color_data = Z;
		19'b1110001010101110100: color_data = Z;
		19'b1110001010101110101: color_data = Z;
		19'b1110001010101110110: color_data = Z;
		19'b1110001100100100110: color_data = Z;
		19'b1110001100100100111: color_data = Z;
		19'b1110001100100101000: color_data = Z;
		19'b1110001100100101001: color_data = Z;
		19'b1110001100100101010: color_data = Z;
		19'b1110001100100101011: color_data = Z;
		19'b1110001100100101100: color_data = Z;
		19'b1110001100100101101: color_data = Z;
		19'b1110001100100101110: color_data = Z;
		19'b1110001100100101111: color_data = Z;
		19'b1110001100100110000: color_data = Z;
		19'b1110001100100110001: color_data = Z;
		19'b1110001100100110010: color_data = Z;
		19'b1110001100100110011: color_data = Z;
		19'b1110001100100110100: color_data = Z;
		19'b1110001100100110101: color_data = Z;
		19'b1110001100100110110: color_data = Z;
		19'b1110001100100110111: color_data = Z;
		19'b1110001100100111000: color_data = Z;
		19'b1110001100100111001: color_data = Z;
		19'b1110001100100111010: color_data = Z;
		19'b1110001100100111011: color_data = Z;
		19'b1110001100100111100: color_data = Z;
		19'b1110001100100111101: color_data = Z;
		19'b1110001100100111110: color_data = Z;
		19'b1110001100100111111: color_data = Z;
		19'b1110001100101000000: color_data = Z;
		19'b1110001100101000001: color_data = Z;
		19'b1110001100101000010: color_data = Z;
		19'b1110001100101000011: color_data = Z;
		19'b1110001100101000100: color_data = Z;
		19'b1110001100101000101: color_data = Z;
		19'b1110001100101000110: color_data = Z;
		19'b1110001100101000111: color_data = Z;
		19'b1110001100101001000: color_data = Z;
		19'b1110001100101001001: color_data = Z;
		19'b1110001100101001010: color_data = Z;
		19'b1110001100101001011: color_data = Z;
		19'b1110001100101001100: color_data = Z;
		19'b1110001100101001101: color_data = Z;
		19'b1110001100101001110: color_data = Z;
		19'b1110001100101001111: color_data = Z;
		19'b1110001100101010000: color_data = Z;
		19'b1110001100101010001: color_data = Z;
		19'b1110001100101010010: color_data = Z;
		19'b1110001100101010011: color_data = Z;
		19'b1110001100101010100: color_data = Z;
		19'b1110001100101010101: color_data = Z;
		19'b1110001100101010110: color_data = Z;
		19'b1110001100101010111: color_data = Z;
		19'b1110001100101011000: color_data = Z;
		19'b1110001100101011001: color_data = Z;
		19'b1110001100101011010: color_data = Z;
		19'b1110001100101011011: color_data = Z;
		19'b1110001100101011100: color_data = Z;
		19'b1110001100101011101: color_data = Z;
		19'b1110001100101011110: color_data = Z;
		19'b1110001100101011111: color_data = Z;
		19'b1110001100101100000: color_data = Z;
		19'b1110001100101100001: color_data = Z;
		19'b1110001100101100010: color_data = Z;
		19'b1110001100101100011: color_data = Z;
		19'b1110001100101100100: color_data = Z;
		19'b1110001100101100101: color_data = Z;
		19'b1110001100101100110: color_data = Z;
		19'b1110001100101100111: color_data = Z;
		19'b1110001100101101000: color_data = Z;
		19'b1110001100101101001: color_data = Z;
		19'b1110001100101101010: color_data = Z;
		19'b1110001100101101011: color_data = Z;
		19'b1110001100101101100: color_data = Z;
		19'b1110001100101101101: color_data = Z;
		19'b1110001100101101110: color_data = Z;
		19'b1110001100101101111: color_data = Z;
		19'b1110001100101110000: color_data = Z;
		19'b1110001100101110001: color_data = Z;
		19'b1110001100101110010: color_data = Z;
		19'b1110001100101110011: color_data = Z;
		19'b1110001100101110100: color_data = Z;
		19'b1110001100101110101: color_data = Z;
		19'b1110001100101110110: color_data = Z;
		19'b1110001110100100000: color_data = Z;
		19'b1110001110100100110: color_data = Z;
		19'b1110001110100100111: color_data = Z;
		19'b1110001110100101000: color_data = Z;
		19'b1110001110100101001: color_data = Z;
		19'b1110001110100101010: color_data = Z;
		19'b1110001110100101011: color_data = Z;
		19'b1110001110100101100: color_data = Z;
		19'b1110001110100101101: color_data = Z;
		19'b1110001110100101110: color_data = Z;
		19'b1110001110100101111: color_data = Z;
		19'b1110001110100110000: color_data = Z;
		19'b1110001110100110001: color_data = Z;
		19'b1110001110100110010: color_data = Z;
		19'b1110001110100110011: color_data = Z;
		19'b1110001110100110100: color_data = Z;
		19'b1110001110100110101: color_data = Z;
		19'b1110001110100110110: color_data = Z;
		19'b1110001110100110111: color_data = Z;
		19'b1110001110100111000: color_data = Z;
		19'b1110001110100111001: color_data = Z;
		19'b1110001110100111010: color_data = Z;
		19'b1110001110100111011: color_data = Z;
		19'b1110001110100111100: color_data = Z;
		19'b1110001110100111101: color_data = Z;
		19'b1110001110100111110: color_data = Z;
		19'b1110001110100111111: color_data = Z;
		19'b1110001110101000000: color_data = Z;
		19'b1110001110101000001: color_data = Z;
		19'b1110001110101000010: color_data = Z;
		19'b1110001110101000011: color_data = Z;
		19'b1110001110101000100: color_data = Z;
		19'b1110001110101000101: color_data = Z;
		19'b1110001110101000110: color_data = Z;
		19'b1110001110101000111: color_data = Z;
		19'b1110001110101001000: color_data = Z;
		19'b1110001110101001001: color_data = Z;
		19'b1110001110101001010: color_data = Z;
		19'b1110001110101001011: color_data = Z;
		19'b1110001110101001100: color_data = Z;
		19'b1110001110101001101: color_data = Z;
		19'b1110001110101001110: color_data = Z;
		19'b1110001110101001111: color_data = Z;
		19'b1110001110101010000: color_data = Z;
		19'b1110001110101010001: color_data = Z;
		19'b1110001110101010010: color_data = Z;
		19'b1110001110101010011: color_data = Z;
		19'b1110001110101010100: color_data = Z;
		19'b1110001110101010101: color_data = Z;
		19'b1110001110101010110: color_data = Z;
		19'b1110001110101010111: color_data = Z;
		19'b1110001110101011000: color_data = Z;
		19'b1110001110101011001: color_data = Z;
		19'b1110001110101011010: color_data = Z;
		19'b1110001110101011011: color_data = Z;
		19'b1110001110101011100: color_data = Z;
		19'b1110001110101011101: color_data = Z;
		19'b1110001110101011110: color_data = Z;
		19'b1110001110101011111: color_data = Z;
		19'b1110001110101100000: color_data = Z;
		19'b1110001110101100001: color_data = Z;
		19'b1110001110101100010: color_data = Z;
		19'b1110001110101100011: color_data = Z;
		19'b1110001110101100100: color_data = Z;
		19'b1110001110101100101: color_data = Z;
		19'b1110001110101100110: color_data = Z;
		19'b1110001110101100111: color_data = Z;
		19'b1110001110101101000: color_data = Z;
		19'b1110001110101101001: color_data = Z;
		19'b1110001110101101010: color_data = Z;
		19'b1110001110101101011: color_data = Z;
		19'b1110001110101101100: color_data = Z;
		19'b1110001110101101101: color_data = Z;
		19'b1110001110101101110: color_data = Z;
		19'b1110001110101101111: color_data = Z;
		19'b1110001110101110000: color_data = Z;
		19'b1110001110101110001: color_data = Z;
		19'b1110001110101110010: color_data = Z;
		19'b1110001110101110011: color_data = Z;
		19'b1110001110101110100: color_data = Z;
		19'b1110001110101110101: color_data = Z;
		19'b1110001110101110110: color_data = Z;
		19'b1110010000100100000: color_data = Z;
		19'b1110010000100100110: color_data = Z;
		19'b1110010000100100111: color_data = Z;
		19'b1110010000100101000: color_data = Z;
		19'b1110010000100101001: color_data = Z;
		19'b1110010000100101010: color_data = Z;
		19'b1110010000100101011: color_data = Z;
		19'b1110010000100101100: color_data = Z;
		19'b1110010000100101101: color_data = Z;
		19'b1110010000100101110: color_data = Z;
		19'b1110010000100101111: color_data = Z;
		19'b1110010000100110000: color_data = Z;
		19'b1110010000100110001: color_data = Z;
		19'b1110010000100110010: color_data = Z;
		19'b1110010000100110011: color_data = Z;
		19'b1110010000100110100: color_data = Z;
		19'b1110010000100110101: color_data = Z;
		19'b1110010000100110110: color_data = Z;
		19'b1110010000100110111: color_data = Z;
		19'b1110010000100111000: color_data = Z;
		19'b1110010000100111001: color_data = Z;
		19'b1110010000100111010: color_data = Z;
		19'b1110010000100111011: color_data = Z;
		19'b1110010000100111100: color_data = Z;
		19'b1110010000100111101: color_data = Z;
		19'b1110010000100111110: color_data = Z;
		19'b1110010000100111111: color_data = Z;
		19'b1110010000101000000: color_data = Z;
		19'b1110010000101000001: color_data = Z;
		19'b1110010000101000010: color_data = Z;
		19'b1110010000101000011: color_data = Z;
		19'b1110010000101000100: color_data = Z;
		19'b1110010000101000101: color_data = Z;
		19'b1110010000101000110: color_data = Z;
		19'b1110010000101000111: color_data = Z;
		19'b1110010000101001000: color_data = Z;
		19'b1110010000101001001: color_data = Z;
		19'b1110010000101001010: color_data = Z;
		19'b1110010000101001011: color_data = Z;
		19'b1110010000101001100: color_data = Z;
		19'b1110010000101001101: color_data = Z;
		19'b1110010000101001110: color_data = Z;
		19'b1110010000101001111: color_data = Z;
		19'b1110010000101010000: color_data = Z;
		19'b1110010000101010001: color_data = Z;
		19'b1110010000101010010: color_data = Z;
		19'b1110010000101010011: color_data = Z;
		19'b1110010000101010100: color_data = Z;
		19'b1110010000101010101: color_data = Z;
		19'b1110010000101010110: color_data = Z;
		19'b1110010000101010111: color_data = Z;
		19'b1110010000101011000: color_data = Z;
		19'b1110010000101011001: color_data = Z;
		19'b1110010000101011010: color_data = Z;
		19'b1110010000101011011: color_data = Z;
		19'b1110010000101011100: color_data = Z;
		19'b1110010000101011101: color_data = Z;
		19'b1110010000101011110: color_data = Z;
		19'b1110010000101011111: color_data = Z;
		19'b1110010000101100000: color_data = Z;
		19'b1110010000101100001: color_data = Z;
		19'b1110010000101100010: color_data = Z;
		19'b1110010000101100011: color_data = Z;
		19'b1110010000101100100: color_data = Z;
		19'b1110010000101100101: color_data = Z;
		19'b1110010000101100110: color_data = Z;
		19'b1110010000101100111: color_data = Z;
		19'b1110010000101101000: color_data = Z;
		19'b1110010000101101001: color_data = Z;
		19'b1110010000101101010: color_data = Z;
		19'b1110010000101101011: color_data = Z;
		19'b1110010000101101100: color_data = Z;
		19'b1110010000101101101: color_data = Z;
		19'b1110010000101101110: color_data = Z;
		19'b1110010000101101111: color_data = Z;
		19'b1110010000101110000: color_data = Z;
		19'b1110010000101110001: color_data = Z;
		19'b1110010000101110010: color_data = Z;
		19'b1110010000101110011: color_data = Z;
		19'b1110010000101110100: color_data = Z;
		19'b1110010000101110101: color_data = Z;
		19'b1110010000101110110: color_data = Z;
		19'b1110010010100100110: color_data = Z;
		19'b1110010010100100111: color_data = Z;
		19'b1110010010100101000: color_data = Z;
		19'b1110010010100101001: color_data = Z;
		19'b1110010010100101010: color_data = Z;
		19'b1110010010100101011: color_data = Z;
		19'b1110010010100101100: color_data = Z;
		19'b1110010010100101101: color_data = Z;
		19'b1110010010100101110: color_data = Z;
		19'b1110010010100101111: color_data = Z;
		19'b1110010010100110000: color_data = Z;
		19'b1110010010100110001: color_data = Z;
		19'b1110010010100110010: color_data = Z;
		19'b1110010010100110011: color_data = Z;
		19'b1110010010100110100: color_data = Z;
		19'b1110010010100110101: color_data = Z;
		19'b1110010010100110110: color_data = Z;
		19'b1110010010100110111: color_data = Z;
		19'b1110010010100111000: color_data = Z;
		19'b1110010010100111001: color_data = Z;
		19'b1110010010100111010: color_data = Z;
		19'b1110010010100111011: color_data = Z;
		19'b1110010010100111100: color_data = Z;
		19'b1110010010100111101: color_data = Z;
		19'b1110010010100111110: color_data = Z;
		19'b1110010010100111111: color_data = Z;
		19'b1110010010101000000: color_data = Z;
		19'b1110010010101000001: color_data = Z;
		19'b1110010010101000010: color_data = Z;
		19'b1110010010101000011: color_data = Z;
		19'b1110010010101000100: color_data = Z;
		19'b1110010010101000101: color_data = Z;
		19'b1110010010101000110: color_data = Z;
		19'b1110010010101000111: color_data = Z;
		19'b1110010010101001000: color_data = Z;
		19'b1110010010101001001: color_data = Z;
		19'b1110010010101001010: color_data = Z;
		19'b1110010010101001011: color_data = Z;
		19'b1110010010101001100: color_data = Z;
		19'b1110010010101001101: color_data = Z;
		19'b1110010010101001110: color_data = Z;
		19'b1110010010101001111: color_data = Z;
		19'b1110010010101010000: color_data = Z;
		19'b1110010010101010001: color_data = Z;
		19'b1110010010101010010: color_data = Z;
		19'b1110010010101010011: color_data = Z;
		19'b1110010010101010100: color_data = Z;
		19'b1110010010101010101: color_data = Z;
		19'b1110010010101010110: color_data = Z;
		19'b1110010010101010111: color_data = Z;
		19'b1110010010101011000: color_data = Z;
		19'b1110010010101011001: color_data = Z;
		19'b1110010010101011010: color_data = Z;
		19'b1110010010101011011: color_data = Z;
		19'b1110010010101011100: color_data = Z;
		19'b1110010010101011101: color_data = Z;
		19'b1110010010101011110: color_data = Z;
		19'b1110010010101011111: color_data = Z;
		19'b1110010010101100000: color_data = Z;
		19'b1110010010101100001: color_data = Z;
		19'b1110010010101100010: color_data = Z;
		19'b1110010010101100011: color_data = Z;
		19'b1110010010101100100: color_data = Z;
		19'b1110010010101100101: color_data = Z;
		19'b1110010010101100110: color_data = Z;
		19'b1110010010101100111: color_data = Z;
		19'b1110010010101101000: color_data = Z;
		19'b1110010010101101001: color_data = Z;
		19'b1110010010101101010: color_data = Z;
		19'b1110010010101101011: color_data = Z;
		19'b1110010010101101100: color_data = Z;
		19'b1110010010101101101: color_data = Z;
		19'b1110010010101101110: color_data = Z;
		19'b1110010010101101111: color_data = Z;
		19'b1110010010101110000: color_data = Z;
		19'b1110010010101110001: color_data = Z;
		19'b1110010010101110010: color_data = Z;
		19'b1110010010101110011: color_data = Z;
		19'b1110010010101110100: color_data = Z;
		19'b1110010010101110101: color_data = Z;
		19'b1110010010101110110: color_data = Z;
		19'b1110010010101110111: color_data = Z;
		19'b1110010100100100110: color_data = Z;
		19'b1110010100100100111: color_data = Z;
		19'b1110010100100101000: color_data = Z;
		19'b1110010100100101001: color_data = Z;
		19'b1110010100100101010: color_data = Z;
		19'b1110010100100101011: color_data = Z;
		19'b1110010100100101100: color_data = Z;
		19'b1110010100100101101: color_data = Z;
		19'b1110010100100101110: color_data = Z;
		19'b1110010100100101111: color_data = Z;
		19'b1110010100100110000: color_data = Z;
		19'b1110010100100110001: color_data = Z;
		19'b1110010100100110010: color_data = Z;
		19'b1110010100100110011: color_data = Z;
		19'b1110010100100110100: color_data = Z;
		19'b1110010100100110101: color_data = Z;
		19'b1110010100100110110: color_data = Z;
		19'b1110010100100110111: color_data = Z;
		19'b1110010100100111000: color_data = Z;
		19'b1110010100100111001: color_data = Z;
		19'b1110010100100111010: color_data = Z;
		19'b1110010100100111011: color_data = Z;
		19'b1110010100100111100: color_data = Z;
		19'b1110010100100111101: color_data = Z;
		19'b1110010100100111110: color_data = Z;
		19'b1110010100100111111: color_data = Z;
		19'b1110010100101000000: color_data = Z;
		19'b1110010100101000001: color_data = Z;
		19'b1110010100101000010: color_data = Z;
		19'b1110010100101000011: color_data = Z;
		19'b1110010100101000100: color_data = Z;
		19'b1110010100101000101: color_data = Z;
		19'b1110010100101000110: color_data = Z;
		19'b1110010100101000111: color_data = Z;
		19'b1110010100101001000: color_data = Z;
		19'b1110010100101001001: color_data = Z;
		19'b1110010100101001010: color_data = Z;
		19'b1110010100101001011: color_data = Z;
		19'b1110010100101001100: color_data = Z;
		19'b1110010100101001101: color_data = Z;
		19'b1110010100101001110: color_data = Z;
		19'b1110010100101001111: color_data = Z;
		19'b1110010100101010000: color_data = Z;
		19'b1110010100101010001: color_data = Z;
		19'b1110010100101010010: color_data = Z;
		19'b1110010100101010011: color_data = Z;
		19'b1110010100101010100: color_data = Z;
		19'b1110010100101010101: color_data = Z;
		19'b1110010100101010110: color_data = Z;
		19'b1110010100101010111: color_data = Z;
		19'b1110010100101011000: color_data = Z;
		19'b1110010100101011001: color_data = Z;
		19'b1110010100101011010: color_data = Z;
		19'b1110010100101011011: color_data = Z;
		19'b1110010100101011100: color_data = Z;
		19'b1110010100101011101: color_data = Z;
		19'b1110010100101011110: color_data = Z;
		19'b1110010100101011111: color_data = Z;
		19'b1110010100101100000: color_data = Z;
		19'b1110010100101100001: color_data = Z;
		19'b1110010100101100010: color_data = Z;
		19'b1110010100101100011: color_data = Z;
		19'b1110010100101100100: color_data = Z;
		19'b1110010100101100101: color_data = Z;
		19'b1110010100101100110: color_data = Z;
		19'b1110010100101100111: color_data = Z;
		19'b1110010100101101000: color_data = Z;
		19'b1110010100101101001: color_data = Z;
		19'b1110010100101101010: color_data = Z;
		19'b1110010100101101011: color_data = Z;
		19'b1110010100101101100: color_data = Z;
		19'b1110010100101101101: color_data = Z;
		19'b1110010100101101110: color_data = Z;
		19'b1110010100101101111: color_data = Z;
		19'b1110010100101110000: color_data = Z;
		19'b1110010100101110001: color_data = Z;
		19'b1110010100101110010: color_data = Z;
		19'b1110010100101110011: color_data = Z;
		19'b1110010100101110100: color_data = Z;
		19'b1110010100101110101: color_data = Z;
		19'b1110010100101110110: color_data = Z;
		19'b1110010100101110111: color_data = Z;
		19'b1110010110100100110: color_data = Z;
		19'b1110010110100100111: color_data = Z;
		19'b1110010110100101000: color_data = Z;
		19'b1110010110100101001: color_data = Z;
		19'b1110010110100101010: color_data = Z;
		19'b1110010110100101011: color_data = Z;
		19'b1110010110100101100: color_data = Z;
		19'b1110010110100101101: color_data = Z;
		19'b1110010110100101110: color_data = Z;
		19'b1110010110100101111: color_data = Z;
		19'b1110010110100110000: color_data = Z;
		19'b1110010110100110001: color_data = Z;
		19'b1110010110100110010: color_data = Z;
		19'b1110010110100110011: color_data = Z;
		19'b1110010110100110100: color_data = Z;
		19'b1110010110100110101: color_data = Z;
		19'b1110010110100110110: color_data = Z;
		19'b1110010110100110111: color_data = Z;
		19'b1110010110100111000: color_data = Z;
		19'b1110010110100111001: color_data = Z;
		19'b1110010110100111010: color_data = Z;
		19'b1110010110100111011: color_data = Z;
		19'b1110010110100111100: color_data = Z;
		19'b1110010110100111101: color_data = Z;
		19'b1110010110100111110: color_data = Z;
		19'b1110010110100111111: color_data = Z;
		19'b1110010110101000000: color_data = Z;
		19'b1110010110101000001: color_data = Z;
		19'b1110010110101000010: color_data = Z;
		19'b1110010110101000011: color_data = Z;
		19'b1110010110101000100: color_data = Z;
		19'b1110010110101000101: color_data = Z;
		19'b1110010110101000110: color_data = Z;
		19'b1110010110101000111: color_data = Z;
		19'b1110010110101001000: color_data = Z;
		19'b1110010110101001001: color_data = Z;
		19'b1110010110101001010: color_data = Z;
		19'b1110010110101001011: color_data = Z;
		19'b1110010110101001100: color_data = Z;
		19'b1110010110101001101: color_data = Z;
		19'b1110010110101001110: color_data = Z;
		19'b1110010110101001111: color_data = Z;
		19'b1110010110101010000: color_data = Z;
		19'b1110010110101010001: color_data = Z;
		19'b1110010110101010010: color_data = Z;
		19'b1110010110101010011: color_data = Z;
		19'b1110010110101010100: color_data = Z;
		19'b1110010110101010101: color_data = Z;
		19'b1110010110101010110: color_data = Z;
		19'b1110010110101010111: color_data = Z;
		19'b1110010110101011000: color_data = Z;
		19'b1110010110101011001: color_data = Z;
		19'b1110010110101011010: color_data = Z;
		19'b1110010110101011011: color_data = Z;
		19'b1110010110101011100: color_data = Z;
		19'b1110010110101011101: color_data = Z;
		19'b1110010110101011110: color_data = Z;
		19'b1110010110101011111: color_data = Z;
		19'b1110010110101100000: color_data = Z;
		19'b1110010110101100001: color_data = Z;
		19'b1110010110101100010: color_data = Z;
		19'b1110010110101100011: color_data = Z;
		19'b1110010110101100100: color_data = Z;
		19'b1110010110101100101: color_data = Z;
		19'b1110010110101100110: color_data = Z;
		19'b1110010110101100111: color_data = Z;
		19'b1110010110101101000: color_data = Z;
		19'b1110010110101101001: color_data = Z;
		19'b1110010110101101010: color_data = Z;
		19'b1110010110101101011: color_data = Z;
		19'b1110010110101101100: color_data = Z;
		19'b1110010110101101101: color_data = Z;
		19'b1110010110101101110: color_data = Z;
		19'b1110010110101101111: color_data = Z;
		19'b1110010110101110000: color_data = Z;
		19'b1110010110101110001: color_data = Z;
		19'b1110010110101110010: color_data = Z;
		19'b1110010110101110011: color_data = Z;
		19'b1110010110101110100: color_data = Z;
		19'b1110010110101110101: color_data = Z;
		19'b1110010110101110110: color_data = Z;
		19'b1110010110101110111: color_data = Z;
		19'b1110011000100100111: color_data = Z;
		19'b1110011000100101000: color_data = Z;
		19'b1110011000100101001: color_data = Z;
		19'b1110011000100101010: color_data = Z;
		19'b1110011000100101011: color_data = Z;
		19'b1110011000100101100: color_data = Z;
		19'b1110011000100101101: color_data = Z;
		19'b1110011000100101110: color_data = Z;
		19'b1110011000100101111: color_data = Z;
		19'b1110011000100110000: color_data = Z;
		19'b1110011000100110001: color_data = Z;
		19'b1110011000100110010: color_data = Z;
		19'b1110011000100110011: color_data = Z;
		19'b1110011000100110100: color_data = Z;
		19'b1110011000100110101: color_data = Z;
		19'b1110011000100110110: color_data = Z;
		19'b1110011000100110111: color_data = Z;
		19'b1110011000100111000: color_data = Z;
		19'b1110011000100111001: color_data = Z;
		19'b1110011000100111010: color_data = Z;
		19'b1110011000100111011: color_data = Z;
		19'b1110011000100111100: color_data = Z;
		19'b1110011000100111101: color_data = Z;
		19'b1110011000100111110: color_data = Z;
		19'b1110011000100111111: color_data = Z;
		19'b1110011000101000000: color_data = Z;
		19'b1110011000101000001: color_data = Z;
		19'b1110011000101000010: color_data = Z;
		19'b1110011000101000011: color_data = Z;
		19'b1110011000101000100: color_data = Z;
		19'b1110011000101000101: color_data = Z;
		19'b1110011000101000110: color_data = Z;
		19'b1110011000101000111: color_data = Z;
		19'b1110011000101001000: color_data = Z;
		19'b1110011000101001001: color_data = Z;
		19'b1110011000101001010: color_data = Z;
		19'b1110011000101001011: color_data = Z;
		19'b1110011000101001100: color_data = Z;
		19'b1110011000101001101: color_data = Z;
		19'b1110011000101001110: color_data = Z;
		19'b1110011000101001111: color_data = Z;
		19'b1110011000101010000: color_data = Z;
		19'b1110011000101010001: color_data = Z;
		19'b1110011000101010010: color_data = Z;
		19'b1110011000101010011: color_data = Z;
		19'b1110011000101010100: color_data = Z;
		19'b1110011000101010101: color_data = Z;
		19'b1110011000101010110: color_data = Z;
		19'b1110011000101010111: color_data = Z;
		19'b1110011000101011000: color_data = Z;
		19'b1110011000101011001: color_data = Z;
		19'b1110011000101011010: color_data = Z;
		19'b1110011000101011011: color_data = Z;
		19'b1110011000101011100: color_data = Z;
		19'b1110011000101011101: color_data = Z;
		19'b1110011000101011110: color_data = Z;
		19'b1110011000101011111: color_data = Z;
		19'b1110011000101100000: color_data = Z;
		19'b1110011000101100001: color_data = Z;
		19'b1110011000101100010: color_data = Z;
		19'b1110011000101100011: color_data = Z;
		19'b1110011000101100100: color_data = Z;
		19'b1110011000101100101: color_data = Z;
		19'b1110011000101100110: color_data = Z;
		19'b1110011000101100111: color_data = Z;
		19'b1110011000101101000: color_data = Z;
		19'b1110011000101101001: color_data = Z;
		19'b1110011000101101010: color_data = Z;
		19'b1110011000101101011: color_data = Z;
		19'b1110011000101101100: color_data = Z;
		19'b1110011000101101101: color_data = Z;
		19'b1110011000101101110: color_data = Z;
		19'b1110011000101101111: color_data = Z;
		19'b1110011000101110000: color_data = Z;
		19'b1110011000101110001: color_data = Z;
		19'b1110011000101110010: color_data = Z;
		19'b1110011000101110011: color_data = Z;
		19'b1110011000101110100: color_data = Z;
		19'b1110011000101110101: color_data = Z;
		19'b1110011000101110110: color_data = Z;
		19'b1110011000101110111: color_data = Z;
		19'b1110011010100100110: color_data = Z;
		19'b1110011010100100111: color_data = Z;
		19'b1110011010100101000: color_data = Z;
		19'b1110011010100101001: color_data = Z;
		19'b1110011010100101010: color_data = Z;
		19'b1110011010100101011: color_data = Z;
		19'b1110011010100101100: color_data = Z;
		19'b1110011010100101101: color_data = Z;
		19'b1110011010100101110: color_data = Z;
		19'b1110011010100101111: color_data = Z;
		19'b1110011010100110000: color_data = Z;
		19'b1110011010100110001: color_data = Z;
		19'b1110011010100110010: color_data = Z;
		19'b1110011010100110011: color_data = Z;
		19'b1110011010100110100: color_data = Z;
		19'b1110011010100110101: color_data = Z;
		19'b1110011010100110110: color_data = Z;
		19'b1110011010100110111: color_data = Z;
		19'b1110011010100111000: color_data = Z;
		19'b1110011010100111001: color_data = Z;
		19'b1110011010100111010: color_data = Z;
		19'b1110011010100111011: color_data = Z;
		19'b1110011010100111100: color_data = Z;
		19'b1110011010100111101: color_data = Z;
		19'b1110011010100111110: color_data = Z;
		19'b1110011010100111111: color_data = Z;
		19'b1110011010101000000: color_data = Z;
		19'b1110011010101000001: color_data = Z;
		19'b1110011010101000010: color_data = Z;
		19'b1110011010101000011: color_data = Z;
		19'b1110011010101000100: color_data = Z;
		19'b1110011010101000101: color_data = Z;
		19'b1110011010101000110: color_data = Z;
		19'b1110011010101000111: color_data = Z;
		19'b1110011010101001000: color_data = Z;
		19'b1110011010101001001: color_data = Z;
		19'b1110011010101001010: color_data = Z;
		19'b1110011010101001011: color_data = Z;
		19'b1110011010101001100: color_data = Z;
		19'b1110011010101001101: color_data = Z;
		19'b1110011010101001110: color_data = Z;
		19'b1110011010101001111: color_data = Z;
		19'b1110011010101010000: color_data = Z;
		19'b1110011010101010001: color_data = Z;
		19'b1110011010101010010: color_data = Z;
		19'b1110011010101010011: color_data = Z;
		19'b1110011010101010100: color_data = Z;
		19'b1110011010101010101: color_data = Z;
		19'b1110011010101010110: color_data = Z;
		19'b1110011010101010111: color_data = Z;
		19'b1110011010101011000: color_data = Z;
		19'b1110011010101011001: color_data = Z;
		19'b1110011010101011010: color_data = Z;
		19'b1110011010101011011: color_data = Z;
		19'b1110011010101011100: color_data = Z;
		19'b1110011010101011101: color_data = Z;
		19'b1110011010101011110: color_data = Z;
		19'b1110011010101011111: color_data = Z;
		19'b1110011010101100000: color_data = Z;
		19'b1110011010101100001: color_data = Z;
		19'b1110011010101100010: color_data = Z;
		19'b1110011010101100011: color_data = Z;
		19'b1110011010101100100: color_data = Z;
		19'b1110011010101100101: color_data = Z;
		19'b1110011010101100110: color_data = Z;
		19'b1110011010101100111: color_data = Z;
		19'b1110011010101101000: color_data = Z;
		19'b1110011010101101001: color_data = Z;
		19'b1110011010101101010: color_data = Z;
		19'b1110011010101101011: color_data = Z;
		19'b1110011010101101100: color_data = Z;
		19'b1110011010101101101: color_data = Z;
		19'b1110011010101101110: color_data = Z;
		19'b1110011010101101111: color_data = Z;
		19'b1110011010101110000: color_data = Z;
		19'b1110011010101110001: color_data = Z;
		19'b1110011010101110010: color_data = Z;
		19'b1110011010101110011: color_data = Z;
		19'b1110011010101110100: color_data = Z;
		19'b1110011010101110101: color_data = Z;
		19'b1110011010101110110: color_data = Z;
		19'b1110011010101110111: color_data = Z;
		19'b1110011100100100110: color_data = Z;
		19'b1110011100100100111: color_data = Z;
		19'b1110011100100101000: color_data = Z;
		19'b1110011100100101001: color_data = Z;
		19'b1110011100100101010: color_data = Z;
		19'b1110011100100101011: color_data = Z;
		19'b1110011100100101100: color_data = Z;
		19'b1110011100100101101: color_data = Z;
		19'b1110011100100101110: color_data = Z;
		19'b1110011100100101111: color_data = Z;
		19'b1110011100100110000: color_data = Z;
		19'b1110011100100110001: color_data = Z;
		19'b1110011100100110010: color_data = Z;
		19'b1110011100100110011: color_data = Z;
		19'b1110011100100110100: color_data = Z;
		19'b1110011100100110101: color_data = Z;
		19'b1110011100100110110: color_data = Z;
		19'b1110011100100110111: color_data = Z;
		19'b1110011100100111000: color_data = Z;
		19'b1110011100100111001: color_data = Z;
		19'b1110011100100111010: color_data = Z;
		19'b1110011100100111011: color_data = Z;
		19'b1110011100100111100: color_data = Z;
		19'b1110011100100111101: color_data = Z;
		19'b1110011100100111110: color_data = Z;
		19'b1110011100100111111: color_data = Z;
		19'b1110011100101000000: color_data = Z;
		19'b1110011100101000001: color_data = Z;
		19'b1110011100101000010: color_data = Z;
		19'b1110011100101000011: color_data = Z;
		19'b1110011100101000100: color_data = Z;
		19'b1110011100101000101: color_data = Z;
		19'b1110011100101000110: color_data = Z;
		19'b1110011100101000111: color_data = Z;
		19'b1110011100101001000: color_data = Z;
		19'b1110011100101001001: color_data = Z;
		19'b1110011100101001010: color_data = Z;
		19'b1110011100101001011: color_data = Z;
		19'b1110011100101001100: color_data = Z;
		19'b1110011100101001101: color_data = Z;
		19'b1110011100101001110: color_data = Z;
		19'b1110011100101001111: color_data = Z;
		19'b1110011100101010000: color_data = Z;
		19'b1110011100101010001: color_data = Z;
		19'b1110011100101010010: color_data = Z;
		19'b1110011100101010011: color_data = Z;
		19'b1110011100101010100: color_data = Z;
		19'b1110011100101010101: color_data = Z;
		19'b1110011100101010110: color_data = Z;
		19'b1110011100101010111: color_data = Z;
		19'b1110011100101011000: color_data = Z;
		19'b1110011100101011001: color_data = Z;
		19'b1110011100101011010: color_data = Z;
		19'b1110011100101011011: color_data = Z;
		19'b1110011100101011100: color_data = Z;
		19'b1110011100101011101: color_data = Z;
		19'b1110011100101011110: color_data = Z;
		19'b1110011100101011111: color_data = Z;
		19'b1110011100101100000: color_data = Z;
		19'b1110011100101100001: color_data = Z;
		19'b1110011100101100010: color_data = Z;
		19'b1110011100101100011: color_data = Z;
		19'b1110011100101100100: color_data = Z;
		19'b1110011100101100101: color_data = Z;
		19'b1110011100101100110: color_data = Z;
		19'b1110011100101100111: color_data = Z;
		19'b1110011100101101000: color_data = Z;
		19'b1110011100101101001: color_data = Z;
		19'b1110011100101101010: color_data = Z;
		19'b1110011100101101011: color_data = Z;
		19'b1110011100101101100: color_data = Z;
		19'b1110011100101101101: color_data = Z;
		19'b1110011100101101110: color_data = Z;
		19'b1110011100101101111: color_data = Z;
		19'b1110011100101110000: color_data = Z;
		19'b1110011100101110001: color_data = Z;
		19'b1110011100101110010: color_data = Z;
		19'b1110011100101110011: color_data = Z;
		19'b1110011100101110100: color_data = Z;
		19'b1110011100101110101: color_data = Z;
		19'b1110011100101110110: color_data = Z;
		19'b1110011110100100111: color_data = Z;
		19'b1110011110100101000: color_data = Z;
		19'b1110011110100101001: color_data = Z;
		19'b1110011110100101010: color_data = Z;
		19'b1110011110100101011: color_data = Z;
		19'b1110011110100101100: color_data = Z;
		19'b1110011110100101101: color_data = Z;
		19'b1110011110100101110: color_data = Z;
		19'b1110011110100101111: color_data = Z;
		19'b1110011110100110000: color_data = Z;
		19'b1110011110100110001: color_data = Z;
		19'b1110011110100110010: color_data = Z;
		19'b1110011110100110011: color_data = Z;
		19'b1110011110100110100: color_data = Z;
		19'b1110011110100110101: color_data = Z;
		19'b1110011110100110110: color_data = Z;
		19'b1110011110100110111: color_data = Z;
		19'b1110011110100111000: color_data = Z;
		19'b1110011110100111001: color_data = Z;
		19'b1110011110100111010: color_data = Z;
		19'b1110011110100111011: color_data = Z;
		19'b1110011110100111100: color_data = Z;
		19'b1110011110100111101: color_data = Z;
		19'b1110011110100111110: color_data = Z;
		19'b1110011110100111111: color_data = Z;
		19'b1110011110101000000: color_data = Z;
		19'b1110011110101000001: color_data = Z;
		19'b1110011110101000010: color_data = Z;
		19'b1110011110101000011: color_data = Z;
		19'b1110011110101000100: color_data = Z;
		19'b1110011110101000101: color_data = Z;
		19'b1110011110101000110: color_data = Z;
		19'b1110011110101000111: color_data = Z;
		19'b1110011110101001000: color_data = Z;
		19'b1110011110101001001: color_data = Z;
		19'b1110011110101001010: color_data = Z;
		19'b1110011110101001011: color_data = Z;
		19'b1110011110101001100: color_data = Z;
		19'b1110011110101001101: color_data = Z;
		19'b1110011110101001110: color_data = Z;
		19'b1110011110101001111: color_data = Z;
		19'b1110011110101010000: color_data = Z;
		19'b1110011110101010001: color_data = Z;
		19'b1110011110101010010: color_data = Z;
		19'b1110011110101010011: color_data = Z;
		19'b1110011110101010100: color_data = Z;
		19'b1110011110101010101: color_data = Z;
		19'b1110011110101010110: color_data = Z;
		19'b1110011110101010111: color_data = Z;
		19'b1110011110101011000: color_data = Z;
		19'b1110011110101011001: color_data = Z;
		19'b1110011110101011010: color_data = Z;
		19'b1110011110101011011: color_data = Z;
		19'b1110011110101011100: color_data = Z;
		19'b1110011110101011101: color_data = Z;
		19'b1110011110101011110: color_data = Z;
		19'b1110011110101011111: color_data = Z;
		19'b1110011110101100000: color_data = Z;
		19'b1110011110101100001: color_data = Z;
		19'b1110011110101100010: color_data = Z;
		19'b1110011110101100011: color_data = Z;
		19'b1110011110101100100: color_data = Z;
		19'b1110011110101100101: color_data = Z;
		19'b1110011110101100110: color_data = Z;
		19'b1110011110101100111: color_data = Z;
		19'b1110011110101101000: color_data = Z;
		19'b1110011110101101001: color_data = Z;
		19'b1110011110101101010: color_data = Z;
		19'b1110011110101101011: color_data = Z;
		19'b1110011110101101100: color_data = Z;
		19'b1110011110101101101: color_data = Z;
		19'b1110011110101101110: color_data = Z;
		19'b1110011110101101111: color_data = Z;
		19'b1110011110101110000: color_data = Z;
		19'b1110011110101110001: color_data = Z;
		19'b1110011110101110010: color_data = Z;
		19'b1110011110101110011: color_data = Z;
		19'b1110011110101110100: color_data = Z;
		19'b1110011110101110101: color_data = Z;
		19'b1110011110101110110: color_data = Z;
		19'b1110100000100101000: color_data = Z;
		19'b1110100000100101001: color_data = Z;
		19'b1110100000100101010: color_data = Z;
		19'b1110100000100101011: color_data = Z;
		19'b1110100000100101100: color_data = Z;
		19'b1110100000100101101: color_data = Z;
		19'b1110100000100101110: color_data = Z;
		19'b1110100000100101111: color_data = Z;
		19'b1110100000100110000: color_data = Z;
		19'b1110100000100110001: color_data = Z;
		19'b1110100000100110010: color_data = Z;
		19'b1110100000100110011: color_data = Z;
		19'b1110100000100110100: color_data = Z;
		19'b1110100000100110101: color_data = Z;
		19'b1110100000100110110: color_data = Z;
		19'b1110100000100110111: color_data = Z;
		19'b1110100000100111000: color_data = Z;
		19'b1110100000100111001: color_data = Z;
		19'b1110100000100111010: color_data = Z;
		19'b1110100000100111011: color_data = Z;
		19'b1110100000100111100: color_data = Z;
		19'b1110100000100111101: color_data = Z;
		19'b1110100000100111110: color_data = Z;
		19'b1110100000100111111: color_data = Z;
		19'b1110100000101000000: color_data = Z;
		19'b1110100000101000001: color_data = Z;
		19'b1110100000101000010: color_data = Z;
		19'b1110100000101000011: color_data = Z;
		19'b1110100000101000100: color_data = Z;
		19'b1110100000101000101: color_data = Z;
		19'b1110100000101000110: color_data = Z;
		19'b1110100000101000111: color_data = Z;
		19'b1110100000101001000: color_data = Z;
		19'b1110100000101001001: color_data = Z;
		19'b1110100000101001010: color_data = Z;
		19'b1110100000101001011: color_data = Z;
		19'b1110100000101001100: color_data = Z;
		19'b1110100000101001101: color_data = Z;
		19'b1110100000101001110: color_data = Z;
		19'b1110100000101001111: color_data = Z;
		19'b1110100000101010000: color_data = Z;
		19'b1110100000101010001: color_data = Z;
		19'b1110100000101010010: color_data = Z;
		19'b1110100000101010011: color_data = Z;
		19'b1110100000101010100: color_data = Z;
		19'b1110100000101010101: color_data = Z;
		19'b1110100000101010110: color_data = Z;
		19'b1110100000101010111: color_data = Z;
		19'b1110100000101011000: color_data = Z;
		19'b1110100000101011001: color_data = Z;
		19'b1110100000101011010: color_data = Z;
		19'b1110100000101011011: color_data = Z;
		19'b1110100000101011100: color_data = Z;
		19'b1110100000101011101: color_data = Z;
		19'b1110100000101011110: color_data = Z;
		19'b1110100000101011111: color_data = Z;
		19'b1110100000101100000: color_data = Z;
		19'b1110100000101100001: color_data = Z;
		19'b1110100000101100010: color_data = Z;
		19'b1110100000101100011: color_data = Z;
		19'b1110100000101100100: color_data = Z;
		19'b1110100000101100101: color_data = Z;
		19'b1110100000101100110: color_data = Z;
		19'b1110100000101100111: color_data = Z;
		19'b1110100000101101000: color_data = Z;
		19'b1110100000101101001: color_data = Z;
		19'b1110100000101101010: color_data = Z;
		19'b1110100000101101011: color_data = Z;
		19'b1110100000101101100: color_data = Z;
		19'b1110100000101101101: color_data = Z;
		19'b1110100000101101110: color_data = Z;
		19'b1110100000101101111: color_data = Z;
		19'b1110100000101110000: color_data = Z;
		19'b1110100000101110001: color_data = Z;
		19'b1110100000101110010: color_data = Z;
		19'b1110100000101110011: color_data = Z;
		19'b1110100000101110100: color_data = Z;
		19'b1110100000101110101: color_data = Z;
		19'b1110100000101110110: color_data = Z;
		19'b1110100010100101001: color_data = Z;
		19'b1110100010100101010: color_data = Z;
		19'b1110100010100101011: color_data = Z;
		19'b1110100010100101100: color_data = Z;
		19'b1110100010100101101: color_data = Z;
		19'b1110100010100101110: color_data = Z;
		19'b1110100010100101111: color_data = Z;
		19'b1110100010100110000: color_data = Z;
		19'b1110100010100110001: color_data = Z;
		19'b1110100010100110010: color_data = Z;
		19'b1110100010100110011: color_data = Z;
		19'b1110100010100110100: color_data = Z;
		19'b1110100010100110101: color_data = Z;
		19'b1110100010100110110: color_data = Z;
		19'b1110100010100110111: color_data = Z;
		19'b1110100010100111000: color_data = Z;
		19'b1110100010100111001: color_data = Z;
		19'b1110100010100111010: color_data = Z;
		19'b1110100010100111011: color_data = Z;
		19'b1110100010100111100: color_data = Z;
		19'b1110100010100111101: color_data = Z;
		19'b1110100010100111110: color_data = Z;
		19'b1110100010100111111: color_data = Z;
		19'b1110100010101000000: color_data = Z;
		19'b1110100010101000001: color_data = Z;
		19'b1110100010101000010: color_data = Z;
		19'b1110100010101000011: color_data = Z;
		19'b1110100010101000100: color_data = Z;
		19'b1110100010101000101: color_data = Z;
		19'b1110100010101000110: color_data = Z;
		19'b1110100010101000111: color_data = Z;
		19'b1110100010101001000: color_data = Z;
		19'b1110100010101001001: color_data = Z;
		19'b1110100010101001010: color_data = Z;
		19'b1110100010101001011: color_data = Z;
		19'b1110100010101001100: color_data = Z;
		19'b1110100010101001101: color_data = Z;
		19'b1110100010101001110: color_data = Z;
		19'b1110100010101001111: color_data = Z;
		19'b1110100010101010000: color_data = Z;
		19'b1110100010101010001: color_data = Z;
		19'b1110100010101010010: color_data = Z;
		19'b1110100010101010011: color_data = Z;
		19'b1110100010101010100: color_data = Z;
		19'b1110100010101010101: color_data = Z;
		19'b1110100010101010110: color_data = Z;
		19'b1110100010101010111: color_data = Z;
		19'b1110100010101011000: color_data = Z;
		19'b1110100010101011001: color_data = Z;
		19'b1110100010101011010: color_data = Z;
		19'b1110100010101011011: color_data = Z;
		19'b1110100010101011100: color_data = Z;
		19'b1110100010101011101: color_data = Z;
		19'b1110100010101011110: color_data = Z;
		19'b1110100010101011111: color_data = Z;
		19'b1110100010101100000: color_data = Z;
		19'b1110100010101100001: color_data = Z;
		19'b1110100010101100010: color_data = Z;
		19'b1110100010101100011: color_data = Z;
		19'b1110100010101100100: color_data = Z;
		19'b1110100010101100101: color_data = Z;
		19'b1110100010101100110: color_data = Z;
		19'b1110100010101100111: color_data = Z;
		19'b1110100010101101000: color_data = Z;
		19'b1110100010101101001: color_data = Z;
		19'b1110100010101101010: color_data = Z;
		19'b1110100010101101011: color_data = Z;
		19'b1110100010101101100: color_data = Z;
		19'b1110100010101101101: color_data = Z;
		19'b1110100010101101110: color_data = Z;
		19'b1110100010101101111: color_data = Z;
		19'b1110100010101110000: color_data = Z;
		19'b1110100010101110001: color_data = Z;
		19'b1110100010101110010: color_data = Z;
		19'b1110100010101110011: color_data = Z;
		19'b1110100010101110100: color_data = Z;
		19'b1110100010101110101: color_data = Z;
		19'b1110100010101110110: color_data = Z;
		19'b1110100100100101001: color_data = Z;
		19'b1110100100100101010: color_data = Z;
		19'b1110100100100101011: color_data = Z;
		19'b1110100100100101100: color_data = Z;
		19'b1110100100100101101: color_data = Z;
		19'b1110100100100101110: color_data = Z;
		19'b1110100100100101111: color_data = Z;
		19'b1110100100100110000: color_data = Z;
		19'b1110100100100110001: color_data = Z;
		19'b1110100100100110010: color_data = Z;
		19'b1110100100100110011: color_data = Z;
		19'b1110100100100110100: color_data = Z;
		19'b1110100100100110101: color_data = Z;
		19'b1110100100100110110: color_data = Z;
		19'b1110100100100110111: color_data = Z;
		19'b1110100100100111000: color_data = Z;
		19'b1110100100100111001: color_data = Z;
		19'b1110100100100111010: color_data = Z;
		19'b1110100100100111011: color_data = Z;
		19'b1110100100100111100: color_data = Z;
		19'b1110100100100111101: color_data = Z;
		19'b1110100100100111110: color_data = Z;
		19'b1110100100100111111: color_data = Z;
		19'b1110100100101000000: color_data = Z;
		19'b1110100100101000001: color_data = Z;
		19'b1110100100101000010: color_data = Z;
		19'b1110100100101000011: color_data = Z;
		19'b1110100100101000100: color_data = Z;
		19'b1110100100101000101: color_data = Z;
		19'b1110100100101000110: color_data = Z;
		19'b1110100100101000111: color_data = Z;
		19'b1110100100101001000: color_data = Z;
		19'b1110100100101001001: color_data = Z;
		19'b1110100100101001010: color_data = Z;
		19'b1110100100101001011: color_data = Z;
		19'b1110100100101001100: color_data = Z;
		19'b1110100100101001101: color_data = Z;
		19'b1110100100101001110: color_data = Z;
		19'b1110100100101001111: color_data = Z;
		19'b1110100100101010000: color_data = Z;
		19'b1110100100101010001: color_data = Z;
		19'b1110100100101010010: color_data = Z;
		19'b1110100100101010011: color_data = Z;
		19'b1110100100101010100: color_data = Z;
		19'b1110100100101010101: color_data = Z;
		19'b1110100100101010110: color_data = Z;
		19'b1110100100101010111: color_data = Z;
		19'b1110100100101011000: color_data = Z;
		19'b1110100100101011001: color_data = Z;
		19'b1110100100101011010: color_data = Z;
		19'b1110100100101011011: color_data = Z;
		19'b1110100100101011100: color_data = Z;
		19'b1110100100101011101: color_data = Z;
		19'b1110100100101011110: color_data = Z;
		19'b1110100100101011111: color_data = Z;
		19'b1110100100101100000: color_data = Z;
		19'b1110100100101100001: color_data = Z;
		19'b1110100100101100010: color_data = Z;
		19'b1110100100101100011: color_data = Z;
		19'b1110100100101100100: color_data = Z;
		19'b1110100100101100101: color_data = Z;
		19'b1110100100101100110: color_data = Z;
		19'b1110100100101100111: color_data = Z;
		19'b1110100100101101000: color_data = Z;
		19'b1110100100101101001: color_data = Z;
		19'b1110100100101101010: color_data = Z;
		19'b1110100100101101011: color_data = Z;
		19'b1110100100101101100: color_data = Z;
		19'b1110100100101101101: color_data = Z;
		19'b1110100100101101110: color_data = Z;
		19'b1110100100101101111: color_data = Z;
		19'b1110100100101110000: color_data = Z;
		19'b1110100100101110001: color_data = Z;
		19'b1110100100101110010: color_data = Z;
		19'b1110100100101110011: color_data = Z;
		19'b1110100100101110100: color_data = Z;
		19'b1110100100101110101: color_data = Z;
		19'b1110100110100101010: color_data = Z;
		19'b1110100110100101011: color_data = Z;
		19'b1110100110100101100: color_data = Z;
		19'b1110100110100101101: color_data = Z;
		19'b1110100110100101110: color_data = Z;
		19'b1110100110100101111: color_data = Z;
		19'b1110100110100110000: color_data = Z;
		19'b1110100110100110001: color_data = Z;
		19'b1110100110100110010: color_data = Z;
		19'b1110100110100110011: color_data = Z;
		19'b1110100110100110100: color_data = Z;
		19'b1110100110100110101: color_data = Z;
		19'b1110100110100110110: color_data = Z;
		19'b1110100110100110111: color_data = Z;
		19'b1110100110100111000: color_data = Z;
		19'b1110100110100111001: color_data = Z;
		19'b1110100110100111010: color_data = Z;
		19'b1110100110100111011: color_data = Z;
		19'b1110100110100111100: color_data = Z;
		19'b1110100110100111101: color_data = Z;
		19'b1110100110100111110: color_data = Z;
		19'b1110100110100111111: color_data = Z;
		19'b1110100110101000000: color_data = Z;
		19'b1110100110101000001: color_data = Z;
		19'b1110100110101000010: color_data = Z;
		19'b1110100110101000011: color_data = Z;
		19'b1110100110101000100: color_data = Z;
		19'b1110100110101000101: color_data = Z;
		19'b1110100110101000110: color_data = Z;
		19'b1110100110101000111: color_data = Z;
		19'b1110100110101001000: color_data = Z;
		19'b1110100110101001001: color_data = Z;
		19'b1110100110101001010: color_data = Z;
		19'b1110100110101001011: color_data = Z;
		19'b1110100110101001100: color_data = Z;
		19'b1110100110101001101: color_data = Z;
		19'b1110100110101001110: color_data = Z;
		19'b1110100110101001111: color_data = Z;
		19'b1110100110101010000: color_data = Z;
		19'b1110100110101010001: color_data = Z;
		19'b1110100110101010010: color_data = Z;
		19'b1110100110101010011: color_data = Z;
		19'b1110100110101010100: color_data = Z;
		19'b1110100110101010101: color_data = Z;
		19'b1110100110101010110: color_data = Z;
		19'b1110100110101010111: color_data = Z;
		19'b1110100110101011000: color_data = Z;
		19'b1110100110101011001: color_data = Z;
		19'b1110100110101011010: color_data = Z;
		19'b1110100110101011011: color_data = Z;
		19'b1110100110101011100: color_data = Z;
		19'b1110100110101011101: color_data = Z;
		19'b1110100110101011110: color_data = Z;
		19'b1110100110101011111: color_data = Z;
		19'b1110100110101100000: color_data = Z;
		19'b1110100110101100001: color_data = Z;
		19'b1110100110101100010: color_data = Z;
		19'b1110100110101100011: color_data = Z;
		19'b1110100110101100100: color_data = Z;
		19'b1110100110101100101: color_data = Z;
		19'b1110100110101100110: color_data = Z;
		19'b1110100110101100111: color_data = Z;
		19'b1110100110101101000: color_data = Z;
		19'b1110100110101101001: color_data = Z;
		19'b1110100110101101010: color_data = Z;
		19'b1110100110101101011: color_data = Z;
		19'b1110100110101101100: color_data = Z;
		19'b1110100110101101101: color_data = Z;
		19'b1110100110101101110: color_data = Z;
		19'b1110100110101101111: color_data = Z;
		19'b1110100110101110000: color_data = Z;
		19'b1110100110101110001: color_data = Z;
		19'b1110100110101110010: color_data = Z;
		19'b1110100110101110011: color_data = Z;
		19'b1110100110101110100: color_data = Z;
		19'b1110100110101110101: color_data = Z;
		19'b1110101000100101010: color_data = Z;
		19'b1110101000100101011: color_data = Z;
		19'b1110101000100101100: color_data = Z;
		19'b1110101000100101101: color_data = Z;
		19'b1110101000100101110: color_data = Z;
		19'b1110101000100101111: color_data = Z;
		19'b1110101000100110000: color_data = Z;
		19'b1110101000100110001: color_data = Z;
		19'b1110101000100110010: color_data = Z;
		19'b1110101000100110011: color_data = Z;
		19'b1110101000100110100: color_data = Z;
		19'b1110101000100110101: color_data = Z;
		19'b1110101000100110110: color_data = Z;
		19'b1110101000100110111: color_data = Z;
		19'b1110101000100111000: color_data = Z;
		19'b1110101000100111001: color_data = Z;
		19'b1110101000100111010: color_data = Z;
		19'b1110101000100111011: color_data = Z;
		19'b1110101000100111100: color_data = Z;
		19'b1110101000100111101: color_data = Z;
		19'b1110101000100111110: color_data = Z;
		19'b1110101000100111111: color_data = Z;
		19'b1110101000101000000: color_data = Z;
		19'b1110101000101000001: color_data = Z;
		19'b1110101000101000010: color_data = Z;
		19'b1110101000101000011: color_data = Z;
		19'b1110101000101000100: color_data = Z;
		19'b1110101000101000101: color_data = Z;
		19'b1110101000101000110: color_data = Z;
		19'b1110101000101000111: color_data = Z;
		19'b1110101000101001000: color_data = Z;
		19'b1110101000101001001: color_data = Z;
		19'b1110101000101001010: color_data = Z;
		19'b1110101000101001011: color_data = Z;
		19'b1110101000101001100: color_data = Z;
		19'b1110101000101001101: color_data = Z;
		19'b1110101000101001110: color_data = Z;
		19'b1110101000101001111: color_data = Z;
		19'b1110101000101010000: color_data = Z;
		19'b1110101000101010001: color_data = Z;
		19'b1110101000101010010: color_data = Z;
		19'b1110101000101010011: color_data = Z;
		19'b1110101000101010100: color_data = Z;
		19'b1110101000101010101: color_data = Z;
		19'b1110101000101010110: color_data = Z;
		19'b1110101000101010111: color_data = Z;
		19'b1110101000101011000: color_data = Z;
		19'b1110101000101011001: color_data = Z;
		19'b1110101000101011010: color_data = Z;
		19'b1110101000101011011: color_data = Z;
		19'b1110101000101011100: color_data = Z;
		19'b1110101000101011101: color_data = Z;
		19'b1110101000101011110: color_data = Z;
		19'b1110101000101011111: color_data = Z;
		19'b1110101000101100000: color_data = Z;
		19'b1110101000101100001: color_data = Z;
		19'b1110101000101100010: color_data = Z;
		19'b1110101000101100011: color_data = Z;
		19'b1110101000101100100: color_data = Z;
		19'b1110101000101100101: color_data = Z;
		19'b1110101000101100110: color_data = Z;
		19'b1110101000101100111: color_data = Z;
		19'b1110101000101101000: color_data = Z;
		19'b1110101000101101001: color_data = Z;
		19'b1110101000101101010: color_data = Z;
		19'b1110101000101101011: color_data = Z;
		19'b1110101000101101100: color_data = Z;
		19'b1110101000101101101: color_data = Z;
		19'b1110101000101101110: color_data = Z;
		19'b1110101000101101111: color_data = Z;
		19'b1110101000101110000: color_data = Z;
		19'b1110101000101110001: color_data = Z;
		19'b1110101000101110010: color_data = Z;
		19'b1110101000101110011: color_data = Z;
		19'b1110101000101110100: color_data = Z;
		19'b1110101010100101011: color_data = Z;
		19'b1110101010100101100: color_data = Z;
		19'b1110101010100101101: color_data = Z;
		19'b1110101010100101110: color_data = Z;
		19'b1110101010100101111: color_data = Z;
		19'b1110101010100110000: color_data = Z;
		19'b1110101010100110001: color_data = Z;
		19'b1110101010100110010: color_data = Z;
		19'b1110101010100110011: color_data = Z;
		19'b1110101010100110100: color_data = Z;
		19'b1110101010100110101: color_data = Z;
		19'b1110101010100110110: color_data = Z;
		19'b1110101010100110111: color_data = Z;
		19'b1110101010100111000: color_data = Z;
		19'b1110101010100111001: color_data = Z;
		19'b1110101010100111010: color_data = Z;
		19'b1110101010100111011: color_data = Z;
		19'b1110101010100111100: color_data = Z;
		19'b1110101010100111101: color_data = Z;
		19'b1110101010100111110: color_data = Z;
		19'b1110101010100111111: color_data = Z;
		19'b1110101010101000000: color_data = Z;
		19'b1110101010101000001: color_data = Z;
		19'b1110101010101000010: color_data = Z;
		19'b1110101010101000011: color_data = Z;
		19'b1110101010101000100: color_data = Z;
		19'b1110101010101000101: color_data = Z;
		19'b1110101010101000110: color_data = Z;
		19'b1110101010101000111: color_data = Z;
		19'b1110101010101001000: color_data = Z;
		19'b1110101010101001001: color_data = Z;
		19'b1110101010101001010: color_data = Z;
		19'b1110101010101001011: color_data = Z;
		19'b1110101010101001100: color_data = Z;
		19'b1110101010101001101: color_data = Z;
		19'b1110101010101001110: color_data = Z;
		19'b1110101010101001111: color_data = Z;
		19'b1110101010101010000: color_data = Z;
		19'b1110101010101010001: color_data = Z;
		19'b1110101010101010010: color_data = Z;
		19'b1110101010101010011: color_data = Z;
		19'b1110101010101010100: color_data = Z;
		19'b1110101010101010101: color_data = Z;
		19'b1110101010101010110: color_data = Z;
		19'b1110101010101010111: color_data = Z;
		19'b1110101010101011000: color_data = Z;
		19'b1110101010101011001: color_data = Z;
		19'b1110101010101011010: color_data = Z;
		19'b1110101010101011011: color_data = Z;
		19'b1110101010101011100: color_data = Z;
		19'b1110101010101011101: color_data = Z;
		19'b1110101010101011110: color_data = Z;
		19'b1110101010101011111: color_data = Z;
		19'b1110101010101100000: color_data = Z;
		19'b1110101010101100001: color_data = Z;
		19'b1110101010101100010: color_data = Z;
		19'b1110101010101100011: color_data = Z;
		19'b1110101010101100100: color_data = Z;
		19'b1110101010101100101: color_data = Z;
		19'b1110101010101100110: color_data = Z;
		19'b1110101010101100111: color_data = Z;
		19'b1110101010101101000: color_data = Z;
		19'b1110101010101101001: color_data = Z;
		19'b1110101010101101010: color_data = Z;
		19'b1110101010101101011: color_data = Z;
		19'b1110101010101101100: color_data = Z;
		19'b1110101010101101101: color_data = Z;
		19'b1110101010101101110: color_data = Z;
		19'b1110101010101101111: color_data = Z;
		19'b1110101010101110000: color_data = Z;
		19'b1110101010101110001: color_data = Z;
		19'b1110101010101110010: color_data = Z;
		19'b1110101010101110011: color_data = Z;
		19'b1110101100100101011: color_data = Z;
		19'b1110101100100101100: color_data = Z;
		19'b1110101100100101101: color_data = Z;
		19'b1110101100100101110: color_data = Z;
		19'b1110101100100101111: color_data = Z;
		19'b1110101100100110000: color_data = Z;
		19'b1110101100100110001: color_data = Z;
		19'b1110101100100110010: color_data = Z;
		19'b1110101100100110011: color_data = Z;
		19'b1110101100100110100: color_data = Z;
		19'b1110101100100110101: color_data = Z;
		19'b1110101100100110110: color_data = Z;
		19'b1110101100100110111: color_data = Z;
		19'b1110101100100111000: color_data = Z;
		19'b1110101100100111001: color_data = Z;
		19'b1110101100100111010: color_data = Z;
		19'b1110101100100111011: color_data = Z;
		19'b1110101100100111100: color_data = Z;
		19'b1110101100100111101: color_data = Z;
		19'b1110101100100111110: color_data = Z;
		19'b1110101100100111111: color_data = Z;
		19'b1110101100101000000: color_data = Z;
		19'b1110101100101000001: color_data = Z;
		19'b1110101100101000010: color_data = Z;
		19'b1110101100101000011: color_data = Z;
		19'b1110101100101000100: color_data = Z;
		19'b1110101100101000101: color_data = Z;
		19'b1110101100101000110: color_data = Z;
		19'b1110101100101000111: color_data = Z;
		19'b1110101100101001000: color_data = Z;
		19'b1110101100101001001: color_data = Z;
		19'b1110101100101001010: color_data = Z;
		19'b1110101100101001011: color_data = Z;
		19'b1110101100101001100: color_data = Z;
		19'b1110101100101001101: color_data = Z;
		19'b1110101100101001110: color_data = Z;
		19'b1110101100101001111: color_data = Z;
		19'b1110101100101010000: color_data = Z;
		19'b1110101100101010001: color_data = Z;
		19'b1110101100101010010: color_data = Z;
		19'b1110101100101010011: color_data = Z;
		19'b1110101100101010100: color_data = Z;
		19'b1110101100101010101: color_data = Z;
		19'b1110101100101010110: color_data = Z;
		19'b1110101100101010111: color_data = Z;
		19'b1110101100101011000: color_data = Z;
		19'b1110101100101011001: color_data = Z;
		19'b1110101100101011010: color_data = Z;
		19'b1110101100101011011: color_data = Z;
		19'b1110101100101011100: color_data = Z;
		19'b1110101100101011101: color_data = Z;
		19'b1110101100101011110: color_data = Z;
		19'b1110101100101011111: color_data = Z;
		19'b1110101100101100000: color_data = Z;
		19'b1110101100101100001: color_data = Z;
		19'b1110101100101100010: color_data = Z;
		19'b1110101100101100011: color_data = Z;
		19'b1110101100101100100: color_data = Z;
		19'b1110101100101100101: color_data = Z;
		19'b1110101100101100110: color_data = Z;
		19'b1110101100101100111: color_data = Z;
		19'b1110101100101101000: color_data = Z;
		19'b1110101100101101001: color_data = Z;
		19'b1110101100101101010: color_data = Z;
		19'b1110101100101101011: color_data = Z;
		19'b1110101100101101100: color_data = Z;
		19'b1110101100101101101: color_data = Z;
		19'b1110101100101101110: color_data = Z;
		19'b1110101100101101111: color_data = Z;
		19'b1110101100101110000: color_data = Z;
		19'b1110101100101110001: color_data = Z;
		19'b1110101100101110010: color_data = Z;
		19'b1110101100101110011: color_data = Z;
		19'b1110101110100101100: color_data = Z;
		19'b1110101110100101101: color_data = Z;
		19'b1110101110100101110: color_data = Z;
		19'b1110101110100101111: color_data = Z;
		19'b1110101110100110000: color_data = Z;
		19'b1110101110100110001: color_data = Z;
		19'b1110101110100110010: color_data = Z;
		19'b1110101110100110011: color_data = Z;
		19'b1110101110100110100: color_data = Z;
		19'b1110101110100110101: color_data = Z;
		19'b1110101110100110110: color_data = Z;
		19'b1110101110100110111: color_data = Z;
		19'b1110101110100111000: color_data = Z;
		19'b1110101110100111001: color_data = Z;
		19'b1110101110100111010: color_data = Z;
		19'b1110101110100111011: color_data = Z;
		19'b1110101110100111100: color_data = Z;
		19'b1110101110100111101: color_data = Z;
		19'b1110101110100111110: color_data = Z;
		19'b1110101110100111111: color_data = Z;
		19'b1110101110101000000: color_data = Z;
		19'b1110101110101000001: color_data = Z;
		19'b1110101110101000010: color_data = Z;
		19'b1110101110101000011: color_data = Z;
		19'b1110101110101000100: color_data = Z;
		19'b1110101110101000101: color_data = Z;
		19'b1110101110101000110: color_data = Z;
		19'b1110101110101000111: color_data = Z;
		19'b1110101110101001000: color_data = Z;
		19'b1110101110101001001: color_data = Z;
		19'b1110101110101001010: color_data = Z;
		19'b1110101110101001011: color_data = Z;
		19'b1110101110101001100: color_data = Z;
		19'b1110101110101001101: color_data = Z;
		19'b1110101110101001110: color_data = Z;
		19'b1110101110101001111: color_data = Z;
		19'b1110101110101010000: color_data = Z;
		19'b1110101110101010001: color_data = Z;
		19'b1110101110101010010: color_data = Z;
		19'b1110101110101010011: color_data = Z;
		19'b1110101110101010100: color_data = Z;
		19'b1110101110101010101: color_data = Z;
		19'b1110101110101010110: color_data = Z;
		19'b1110101110101010111: color_data = Z;
		19'b1110101110101011000: color_data = Z;
		19'b1110101110101011001: color_data = Z;
		19'b1110101110101011010: color_data = Z;
		19'b1110101110101011011: color_data = Z;
		19'b1110101110101011100: color_data = Z;
		19'b1110101110101011101: color_data = Z;
		19'b1110101110101011110: color_data = Z;
		19'b1110101110101011111: color_data = Z;
		19'b1110101110101100000: color_data = Z;
		19'b1110101110101100001: color_data = Z;
		19'b1110101110101100010: color_data = Z;
		19'b1110101110101100011: color_data = Z;
		19'b1110101110101100100: color_data = Z;
		19'b1110101110101100101: color_data = Z;
		19'b1110101110101100110: color_data = Z;
		19'b1110101110101100111: color_data = Z;
		19'b1110101110101101000: color_data = Z;
		19'b1110101110101101001: color_data = Z;
		19'b1110101110101101010: color_data = Z;
		19'b1110101110101101011: color_data = Z;
		19'b1110101110101101100: color_data = Z;
		19'b1110101110101101101: color_data = Z;
		19'b1110101110101101110: color_data = Z;
		19'b1110101110101101111: color_data = Z;
		19'b1110101110101110000: color_data = Z;
		19'b1110101110101110001: color_data = Z;
		19'b1110101110101110010: color_data = Z;
		19'b1110101110101110011: color_data = Z;
		19'b1110110000100101101: color_data = Z;
		19'b1110110000100101110: color_data = Z;
		19'b1110110000100101111: color_data = Z;
		19'b1110110000100110000: color_data = Z;
		19'b1110110000100110001: color_data = Z;
		19'b1110110000100110010: color_data = Z;
		19'b1110110000100110011: color_data = Z;
		19'b1110110000100110100: color_data = Z;
		19'b1110110000100110101: color_data = Z;
		19'b1110110000100110110: color_data = Z;
		19'b1110110000100110111: color_data = Z;
		19'b1110110000100111000: color_data = Z;
		19'b1110110000100111001: color_data = Z;
		19'b1110110000100111010: color_data = Z;
		19'b1110110000100111011: color_data = Z;
		19'b1110110000100111100: color_data = Z;
		19'b1110110000100111101: color_data = Z;
		19'b1110110000100111110: color_data = Z;
		19'b1110110000100111111: color_data = Z;
		19'b1110110000101000000: color_data = Z;
		19'b1110110000101000001: color_data = Z;
		19'b1110110000101000010: color_data = Z;
		19'b1110110000101000011: color_data = Z;
		19'b1110110000101000100: color_data = Z;
		19'b1110110000101000101: color_data = Z;
		19'b1110110000101000110: color_data = Z;
		19'b1110110000101000111: color_data = Z;
		19'b1110110000101001000: color_data = Z;
		19'b1110110000101001001: color_data = Z;
		19'b1110110000101001010: color_data = Z;
		19'b1110110000101001011: color_data = Z;
		19'b1110110000101001100: color_data = Z;
		19'b1110110000101001101: color_data = Z;
		19'b1110110000101001110: color_data = Z;
		19'b1110110000101001111: color_data = Z;
		19'b1110110000101010000: color_data = Z;
		19'b1110110000101010001: color_data = Z;
		19'b1110110000101010010: color_data = Z;
		19'b1110110000101010011: color_data = Z;
		19'b1110110000101010100: color_data = Z;
		19'b1110110000101010101: color_data = Z;
		19'b1110110000101010110: color_data = Z;
		19'b1110110000101010111: color_data = Z;
		19'b1110110000101011000: color_data = Z;
		19'b1110110000101011001: color_data = Z;
		19'b1110110000101011010: color_data = Z;
		19'b1110110000101011011: color_data = Z;
		19'b1110110000101011100: color_data = Z;
		19'b1110110000101011101: color_data = Z;
		19'b1110110000101011110: color_data = Z;
		19'b1110110000101011111: color_data = Z;
		19'b1110110000101100000: color_data = Z;
		19'b1110110000101100001: color_data = Z;
		19'b1110110000101100010: color_data = Z;
		19'b1110110000101100011: color_data = Z;
		19'b1110110000101100100: color_data = Z;
		19'b1110110000101100101: color_data = Z;
		19'b1110110000101100110: color_data = Z;
		19'b1110110000101100111: color_data = Z;
		19'b1110110000101101000: color_data = Z;
		19'b1110110000101101001: color_data = Z;
		19'b1110110000101101010: color_data = Z;
		19'b1110110000101101011: color_data = Z;
		19'b1110110000101101100: color_data = Z;
		19'b1110110000101101101: color_data = Z;
		19'b1110110000101101110: color_data = Z;
		19'b1110110000101101111: color_data = Z;
		19'b1110110000101110000: color_data = Z;
		19'b1110110000101110001: color_data = Z;
		19'b1110110000101110010: color_data = Z;
		19'b1110110010100101101: color_data = Z;
		19'b1110110010100101110: color_data = Z;
		19'b1110110010100101111: color_data = Z;
		19'b1110110010100110000: color_data = Z;
		19'b1110110010100110001: color_data = Z;
		19'b1110110010100110010: color_data = Z;
		19'b1110110010100110011: color_data = Z;
		19'b1110110010100110100: color_data = Z;
		19'b1110110010100110101: color_data = Z;
		19'b1110110010100110110: color_data = Z;
		19'b1110110010100110111: color_data = Z;
		19'b1110110010100111000: color_data = Z;
		19'b1110110010100111001: color_data = Z;
		19'b1110110010100111010: color_data = Z;
		19'b1110110010100111011: color_data = Z;
		19'b1110110010100111100: color_data = Z;
		19'b1110110010100111101: color_data = Z;
		19'b1110110010100111110: color_data = Z;
		19'b1110110010100111111: color_data = Z;
		19'b1110110010101000000: color_data = Z;
		19'b1110110010101000001: color_data = Z;
		19'b1110110010101000010: color_data = Z;
		19'b1110110010101000011: color_data = Z;
		19'b1110110010101000100: color_data = Z;
		19'b1110110010101000101: color_data = Z;
		19'b1110110010101000110: color_data = Z;
		19'b1110110010101000111: color_data = Z;
		19'b1110110010101001000: color_data = Z;
		19'b1110110010101001001: color_data = Z;
		19'b1110110010101001010: color_data = Z;
		19'b1110110010101001011: color_data = Z;
		19'b1110110010101001100: color_data = Z;
		19'b1110110010101001101: color_data = Z;
		19'b1110110010101001110: color_data = Z;
		19'b1110110010101001111: color_data = Z;
		19'b1110110010101010000: color_data = Z;
		19'b1110110010101010001: color_data = Z;
		19'b1110110010101010010: color_data = Z;
		19'b1110110010101010011: color_data = Z;
		19'b1110110010101010100: color_data = Z;
		19'b1110110010101010101: color_data = Z;
		19'b1110110010101010110: color_data = Z;
		19'b1110110010101010111: color_data = Z;
		19'b1110110010101011000: color_data = Z;
		19'b1110110010101011001: color_data = Z;
		19'b1110110010101011010: color_data = Z;
		19'b1110110010101011011: color_data = Z;
		19'b1110110010101011100: color_data = Z;
		19'b1110110010101011101: color_data = Z;
		19'b1110110010101011110: color_data = Z;
		19'b1110110010101011111: color_data = Z;
		19'b1110110010101100000: color_data = Z;
		19'b1110110010101100001: color_data = Z;
		19'b1110110010101100010: color_data = Z;
		19'b1110110010101100011: color_data = Z;
		19'b1110110010101100100: color_data = Z;
		19'b1110110010101100101: color_data = Z;
		19'b1110110010101100110: color_data = Z;
		19'b1110110010101100111: color_data = Z;
		19'b1110110010101101000: color_data = Z;
		19'b1110110010101101001: color_data = Z;
		19'b1110110010101101010: color_data = Z;
		19'b1110110010101101011: color_data = Z;
		19'b1110110010101101100: color_data = Z;
		19'b1110110010101101101: color_data = Z;
		19'b1110110010101101110: color_data = Z;
		19'b1110110010101101111: color_data = Z;
		19'b1110110010101110000: color_data = Z;
		19'b1110110010101110001: color_data = Z;
		19'b1110110100100101110: color_data = Z;
		19'b1110110100100101111: color_data = Z;
		19'b1110110100100110000: color_data = Z;
		19'b1110110100100110001: color_data = Z;
		19'b1110110100100110010: color_data = Z;
		19'b1110110100100110011: color_data = Z;
		19'b1110110100100110100: color_data = Z;
		19'b1110110100100110101: color_data = Z;
		19'b1110110100100110110: color_data = Z;
		19'b1110110100100110111: color_data = Z;
		19'b1110110100100111000: color_data = Z;
		19'b1110110100100111001: color_data = Z;
		19'b1110110100100111010: color_data = Z;
		19'b1110110100100111011: color_data = Z;
		19'b1110110100100111100: color_data = Z;
		19'b1110110100100111101: color_data = Z;
		19'b1110110100100111110: color_data = Z;
		19'b1110110100100111111: color_data = Z;
		19'b1110110100101000000: color_data = Z;
		19'b1110110100101000001: color_data = Z;
		19'b1110110100101000010: color_data = Z;
		19'b1110110100101000011: color_data = Z;
		19'b1110110100101000100: color_data = Z;
		19'b1110110100101000101: color_data = Z;
		19'b1110110100101000110: color_data = Z;
		19'b1110110100101000111: color_data = Z;
		19'b1110110100101001000: color_data = Z;
		19'b1110110100101001001: color_data = Z;
		19'b1110110100101001010: color_data = Z;
		19'b1110110100101001011: color_data = Z;
		19'b1110110100101001100: color_data = Z;
		19'b1110110100101001101: color_data = Z;
		19'b1110110100101001110: color_data = Z;
		19'b1110110100101001111: color_data = Z;
		19'b1110110100101010000: color_data = Z;
		19'b1110110100101010001: color_data = Z;
		19'b1110110100101010010: color_data = Z;
		19'b1110110100101010011: color_data = Z;
		19'b1110110100101010100: color_data = Z;
		19'b1110110100101010101: color_data = Z;
		19'b1110110100101010110: color_data = Z;
		19'b1110110100101010111: color_data = Z;
		19'b1110110100101011000: color_data = Z;
		19'b1110110100101011001: color_data = Z;
		19'b1110110100101011010: color_data = Z;
		19'b1110110100101011011: color_data = Z;
		19'b1110110100101011100: color_data = Z;
		19'b1110110100101011101: color_data = Z;
		19'b1110110100101011110: color_data = Z;
		19'b1110110100101011111: color_data = Z;
		19'b1110110100101100000: color_data = Z;
		19'b1110110100101100001: color_data = Z;
		19'b1110110100101100010: color_data = Z;
		19'b1110110100101100011: color_data = Z;
		19'b1110110100101100100: color_data = Z;
		19'b1110110100101100101: color_data = Z;
		19'b1110110100101100110: color_data = Z;
		19'b1110110100101100111: color_data = Z;
		19'b1110110100101101000: color_data = Z;
		19'b1110110100101101001: color_data = Z;
		19'b1110110100101101010: color_data = Z;
		19'b1110110100101101011: color_data = Z;
		19'b1110110100101101100: color_data = Z;
		19'b1110110100101101101: color_data = Z;
		19'b1110110100101101110: color_data = Z;
		19'b1110110100101101111: color_data = Z;
		19'b1110110100101110000: color_data = Z;
		19'b1110110110100101111: color_data = Z;
		19'b1110110110100110000: color_data = Z;
		19'b1110110110100110001: color_data = Z;
		19'b1110110110100110010: color_data = Z;
		19'b1110110110100110011: color_data = Z;
		19'b1110110110100110100: color_data = Z;
		19'b1110110110100110101: color_data = Z;
		19'b1110110110100110110: color_data = Z;
		19'b1110110110100110111: color_data = Z;
		19'b1110110110100111000: color_data = Z;
		19'b1110110110100111001: color_data = Z;
		19'b1110110110100111010: color_data = Z;
		19'b1110110110100111011: color_data = Z;
		19'b1110110110100111100: color_data = Z;
		19'b1110110110100111101: color_data = Z;
		19'b1110110110100111110: color_data = Z;
		19'b1110110110100111111: color_data = Z;
		19'b1110110110101000000: color_data = Z;
		19'b1110110110101000001: color_data = Z;
		19'b1110110110101000010: color_data = Z;
		19'b1110110110101000011: color_data = Z;
		19'b1110110110101000100: color_data = Z;
		19'b1110110110101000101: color_data = Z;
		19'b1110110110101000110: color_data = Z;
		19'b1110110110101000111: color_data = Z;
		19'b1110110110101001000: color_data = Z;
		19'b1110110110101001001: color_data = Z;
		19'b1110110110101001010: color_data = Z;
		19'b1110110110101001011: color_data = Z;
		19'b1110110110101001100: color_data = Z;
		19'b1110110110101001101: color_data = Z;
		19'b1110110110101001110: color_data = Z;
		19'b1110110110101001111: color_data = Z;
		19'b1110110110101010000: color_data = Z;
		19'b1110110110101010001: color_data = Z;
		19'b1110110110101010010: color_data = Z;
		19'b1110110110101010011: color_data = Z;
		19'b1110110110101010100: color_data = Z;
		19'b1110110110101010101: color_data = Z;
		19'b1110110110101010110: color_data = Z;
		19'b1110110110101010111: color_data = Z;
		19'b1110110110101011000: color_data = Z;
		19'b1110110110101011001: color_data = Z;
		19'b1110110110101011010: color_data = Z;
		19'b1110110110101011011: color_data = Z;
		19'b1110110110101011100: color_data = Z;
		19'b1110110110101011101: color_data = Z;
		19'b1110110110101011110: color_data = Z;
		19'b1110110110101011111: color_data = Z;
		19'b1110110110101100000: color_data = Z;
		19'b1110110110101100001: color_data = Z;
		19'b1110110110101100010: color_data = Z;
		19'b1110110110101100011: color_data = Z;
		19'b1110110110101100100: color_data = Z;
		19'b1110110110101100101: color_data = Z;
		19'b1110110110101100110: color_data = Z;
		19'b1110110110101100111: color_data = Z;
		19'b1110110110101101000: color_data = Z;
		19'b1110110110101101001: color_data = Z;
		19'b1110110110101101010: color_data = Z;
		19'b1110110110101101011: color_data = Z;
		19'b1110110110101101100: color_data = Z;
		19'b1110110110101101101: color_data = Z;
		19'b1110110110101101110: color_data = Z;
		19'b1110110110101101111: color_data = Z;
		19'b1110111000100110000: color_data = Z;
		19'b1110111000100110001: color_data = Z;
		19'b1110111000100110010: color_data = Z;
		19'b1110111000100110011: color_data = Z;
		19'b1110111000100110100: color_data = Z;
		19'b1110111000100110101: color_data = Z;
		19'b1110111000100110110: color_data = Z;
		19'b1110111000100110111: color_data = Z;
		19'b1110111000100111000: color_data = Z;
		19'b1110111000100111001: color_data = Z;
		19'b1110111000100111010: color_data = Z;
		19'b1110111000100111011: color_data = Z;
		19'b1110111000100111100: color_data = Z;
		19'b1110111000100111101: color_data = Z;
		19'b1110111000100111110: color_data = Z;
		19'b1110111000100111111: color_data = Z;
		19'b1110111000101000000: color_data = Z;
		19'b1110111000101000001: color_data = Z;
		19'b1110111000101000010: color_data = Z;
		19'b1110111000101000011: color_data = Z;
		19'b1110111000101000100: color_data = Z;
		19'b1110111000101000101: color_data = Z;
		19'b1110111000101000110: color_data = Z;
		19'b1110111000101000111: color_data = Z;
		19'b1110111000101001000: color_data = Z;
		19'b1110111000101001001: color_data = Z;
		19'b1110111000101001010: color_data = Z;
		19'b1110111000101001011: color_data = Z;
		19'b1110111000101001100: color_data = Z;
		19'b1110111000101001101: color_data = Z;
		19'b1110111000101001110: color_data = Z;
		19'b1110111000101001111: color_data = Z;
		19'b1110111000101010000: color_data = Z;
		19'b1110111000101010001: color_data = Z;
		19'b1110111000101010010: color_data = Z;
		19'b1110111000101010011: color_data = Z;
		19'b1110111000101010100: color_data = Z;
		19'b1110111000101010101: color_data = Z;
		19'b1110111000101010110: color_data = Z;
		19'b1110111000101010111: color_data = Z;
		19'b1110111000101011000: color_data = Z;
		19'b1110111000101011001: color_data = Z;
		19'b1110111000101011010: color_data = Z;
		19'b1110111000101011011: color_data = Z;
		19'b1110111000101011100: color_data = Z;
		19'b1110111000101011101: color_data = Z;
		19'b1110111000101011110: color_data = Z;
		19'b1110111000101011111: color_data = Z;
		19'b1110111000101100000: color_data = Z;
		19'b1110111000101100001: color_data = Z;
		19'b1110111000101100010: color_data = Z;
		19'b1110111000101100011: color_data = Z;
		19'b1110111000101100100: color_data = Z;
		19'b1110111000101100101: color_data = Z;
		19'b1110111000101100110: color_data = Z;
		19'b1110111000101100111: color_data = Z;
		19'b1110111000101101000: color_data = Z;
		19'b1110111000101101001: color_data = Z;
		19'b1110111000101101010: color_data = Z;
		19'b1110111000101101011: color_data = Z;
		19'b1110111000101101100: color_data = Z;
		19'b1110111000101101101: color_data = Z;
		19'b1110111000101101110: color_data = Z;
		19'b1110111010100110001: color_data = Z;
		19'b1110111010100110010: color_data = Z;
		19'b1110111010100110011: color_data = Z;
		19'b1110111010100110100: color_data = Z;
		19'b1110111010100110101: color_data = Z;
		19'b1110111010100110110: color_data = Z;
		19'b1110111010100110111: color_data = Z;
		19'b1110111010100111000: color_data = Z;
		19'b1110111010100111001: color_data = Z;
		19'b1110111010100111010: color_data = Z;
		19'b1110111010100111011: color_data = Z;
		19'b1110111010100111100: color_data = Z;
		19'b1110111010100111101: color_data = Z;
		19'b1110111010100111110: color_data = Z;
		19'b1110111010100111111: color_data = Z;
		19'b1110111010101000000: color_data = Z;
		19'b1110111010101000001: color_data = Z;
		19'b1110111010101000010: color_data = Z;
		19'b1110111010101000011: color_data = Z;
		19'b1110111010101000100: color_data = Z;
		19'b1110111010101000101: color_data = Z;
		19'b1110111010101000110: color_data = Z;
		19'b1110111010101000111: color_data = Z;
		19'b1110111010101001000: color_data = Z;
		19'b1110111010101001001: color_data = Z;
		19'b1110111010101001010: color_data = Z;
		19'b1110111010101001011: color_data = Z;
		19'b1110111010101001100: color_data = Z;
		19'b1110111010101001101: color_data = Z;
		19'b1110111010101001110: color_data = Z;
		19'b1110111010101001111: color_data = Z;
		19'b1110111010101010000: color_data = Z;
		19'b1110111010101010001: color_data = Z;
		19'b1110111010101010010: color_data = Z;
		19'b1110111010101010011: color_data = Z;
		19'b1110111010101010100: color_data = Z;
		19'b1110111010101010101: color_data = Z;
		19'b1110111010101010110: color_data = Z;
		19'b1110111010101010111: color_data = Z;
		19'b1110111010101011000: color_data = Z;
		19'b1110111010101011001: color_data = Z;
		19'b1110111010101011010: color_data = Z;
		19'b1110111010101011011: color_data = Z;
		19'b1110111010101011100: color_data = Z;
		19'b1110111010101011101: color_data = Z;
		19'b1110111010101011110: color_data = Z;
		19'b1110111010101011111: color_data = Z;
		19'b1110111010101100000: color_data = Z;
		19'b1110111010101100001: color_data = Z;
		19'b1110111010101100010: color_data = Z;
		19'b1110111010101100011: color_data = Z;
		19'b1110111010101100100: color_data = Z;
		19'b1110111010101100101: color_data = Z;
		19'b1110111010101100110: color_data = Z;
		19'b1110111010101100111: color_data = Z;
		19'b1110111010101101000: color_data = Z;
		19'b1110111010101101001: color_data = Z;
		19'b1110111010101101010: color_data = Z;
		19'b1110111010101101011: color_data = Z;
		19'b1110111010101101100: color_data = Z;
		19'b1110111010101101101: color_data = Z;
		19'b1110111010101101110: color_data = Z;
		19'b1110111100100110010: color_data = Z;
		19'b1110111100100110011: color_data = Z;
		19'b1110111100100110100: color_data = Z;
		19'b1110111100100110101: color_data = Z;
		19'b1110111100100110110: color_data = Z;
		19'b1110111100100110111: color_data = Z;
		19'b1110111100100111000: color_data = Z;
		19'b1110111100100111001: color_data = Z;
		19'b1110111100100111010: color_data = Z;
		19'b1110111100100111011: color_data = Z;
		19'b1110111100100111100: color_data = Z;
		19'b1110111100100111101: color_data = Z;
		19'b1110111100100111110: color_data = Z;
		19'b1110111100100111111: color_data = Z;
		19'b1110111100101000000: color_data = Z;
		19'b1110111100101000001: color_data = Z;
		19'b1110111100101000010: color_data = Z;
		19'b1110111100101000011: color_data = Z;
		19'b1110111100101000100: color_data = Z;
		19'b1110111100101000101: color_data = Z;
		19'b1110111100101000110: color_data = Z;
		19'b1110111100101000111: color_data = Z;
		19'b1110111100101001000: color_data = Z;
		19'b1110111100101001001: color_data = Z;
		19'b1110111100101001010: color_data = Z;
		19'b1110111100101001011: color_data = Z;
		19'b1110111100101001100: color_data = Z;
		19'b1110111100101001101: color_data = Z;
		19'b1110111100101001110: color_data = Z;
		19'b1110111100101001111: color_data = Z;
		19'b1110111100101010000: color_data = Z;
		19'b1110111100101010001: color_data = Z;
		19'b1110111100101010010: color_data = Z;
		19'b1110111100101010011: color_data = Z;
		19'b1110111100101010100: color_data = Z;
		19'b1110111100101010101: color_data = Z;
		19'b1110111100101010110: color_data = Z;
		19'b1110111100101010111: color_data = Z;
		19'b1110111100101011000: color_data = Z;
		19'b1110111100101011001: color_data = Z;
		19'b1110111100101011010: color_data = Z;
		19'b1110111100101011011: color_data = Z;
		19'b1110111100101011100: color_data = Z;
		19'b1110111100101011101: color_data = Z;
		19'b1110111100101011110: color_data = Z;
		19'b1110111100101011111: color_data = Z;
		19'b1110111100101100000: color_data = Z;
		19'b1110111100101100001: color_data = Z;
		19'b1110111100101100010: color_data = Z;
		19'b1110111100101100011: color_data = Z;
		19'b1110111100101100100: color_data = Z;
		19'b1110111100101100101: color_data = Z;
		19'b1110111100101100110: color_data = Z;
		19'b1110111100101100111: color_data = Z;
		19'b1110111100101101000: color_data = Z;
		19'b1110111100101101001: color_data = Z;
		19'b1110111100101101010: color_data = Z;
		19'b1110111100101101011: color_data = Z;
		19'b1110111100101101100: color_data = Z;
		19'b1110111100101101101: color_data = Z;
		19'b1110111110100110011: color_data = Z;
		19'b1110111110100110100: color_data = Z;
		19'b1110111110100110101: color_data = Z;
		19'b1110111110100110110: color_data = Z;
		19'b1110111110100110111: color_data = Z;
		19'b1110111110100111000: color_data = Z;
		19'b1110111110100111001: color_data = Z;
		19'b1110111110100111010: color_data = Z;
		19'b1110111110100111011: color_data = Z;
		19'b1110111110100111100: color_data = Z;
		19'b1110111110100111101: color_data = Z;
		19'b1110111110100111110: color_data = Z;
		19'b1110111110100111111: color_data = Z;
		19'b1110111110101000000: color_data = Z;
		19'b1110111110101000001: color_data = Z;
		19'b1110111110101000010: color_data = Z;
		19'b1110111110101000011: color_data = Z;
		19'b1110111110101000100: color_data = Z;
		19'b1110111110101000101: color_data = Z;
		19'b1110111110101000110: color_data = Z;
		19'b1110111110101000111: color_data = Z;
		19'b1110111110101001000: color_data = Z;
		19'b1110111110101001001: color_data = Z;
		19'b1110111110101001010: color_data = Z;
		19'b1110111110101001011: color_data = Z;
		19'b1110111110101001100: color_data = Z;
		19'b1110111110101001101: color_data = Z;
		19'b1110111110101001110: color_data = Z;
		19'b1110111110101001111: color_data = Z;
		19'b1110111110101010000: color_data = Z;
		19'b1110111110101010001: color_data = Z;
		19'b1110111110101010010: color_data = Z;
		19'b1110111110101010011: color_data = Z;
		19'b1110111110101010100: color_data = Z;
		19'b1110111110101010101: color_data = Z;
		19'b1110111110101010110: color_data = Z;
		19'b1110111110101010111: color_data = Z;
		19'b1110111110101011000: color_data = Z;
		19'b1110111110101011001: color_data = Z;
		19'b1110111110101011010: color_data = Z;
		19'b1110111110101011011: color_data = Z;
		19'b1110111110101011100: color_data = Z;
		19'b1110111110101011101: color_data = Z;
		19'b1110111110101011110: color_data = Z;
		19'b1110111110101011111: color_data = Z;
		19'b1110111110101100000: color_data = Z;
		19'b1110111110101100001: color_data = Z;
		19'b1110111110101100010: color_data = Z;
		19'b1110111110101100011: color_data = Z;
		19'b1110111110101100100: color_data = Z;
		19'b1110111110101100101: color_data = Z;
		19'b1110111110101100110: color_data = Z;
		19'b1110111110101100111: color_data = Z;
		19'b1110111110101101000: color_data = Z;
		19'b1110111110101101001: color_data = Z;
		19'b1110111110101101010: color_data = Z;
		19'b1110111110101101011: color_data = Z;
		19'b1110111110101101100: color_data = Z;
		19'b1110111110101101101: color_data = Z;
		default: color_data = 12'b000000000000;
	endcase
endmodule