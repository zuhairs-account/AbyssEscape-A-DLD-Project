module newNew_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		14'b00000001001100: color_data = 12'b010100000000;
		14'b00000001001101: color_data = 12'b101000000000;
		14'b00000001001110: color_data = 12'b101000000000;
		14'b00000001001111: color_data = 12'b101000000000;
		14'b00000001010000: color_data = 12'b101000000000;
		14'b00000001010001: color_data = 12'b101000000000;
		14'b00000001010010: color_data = 12'b101000000000;
		14'b00000001010011: color_data = 12'b101000000000;
		14'b00000001010100: color_data = 12'b101000000000;
		14'b00000001010101: color_data = 12'b101000000000;
		14'b00000001010110: color_data = 12'b101000000000;
		14'b00000001010111: color_data = 12'b101000000000;
		14'b00000001011000: color_data = 12'b101000000000;
		14'b00000001011001: color_data = 12'b010100000000;
		14'b00000010111100: color_data = 12'b010100000000;
		14'b00000010111101: color_data = 12'b010100000000;
		14'b00000010111110: color_data = 12'b010100000000;
		14'b00000010111111: color_data = 12'b010100000000;
		14'b00000011000001: color_data = 12'b010100000000;
		14'b00000011001101: color_data = 12'b010100000000;
		14'b00000011001110: color_data = 12'b101000000000;
		14'b00000011001111: color_data = 12'b101000000000;
		14'b00000011010000: color_data = 12'b101000000000;
		14'b00000011010001: color_data = 12'b101000000000;
		14'b00000011010010: color_data = 12'b101000000000;
		14'b00000011010011: color_data = 12'b101000000000;
		14'b00000011010100: color_data = 12'b101000000000;
		14'b00000011010101: color_data = 12'b101000000000;
		14'b00000011010110: color_data = 12'b101000000000;
		14'b00000011010111: color_data = 12'b101000000000;
		14'b00000011011000: color_data = 12'b101000000000;
		14'b00000011011001: color_data = 12'b010100000000;
		14'b00000100010010: color_data = 12'b010100000000;
		14'b00000100010011: color_data = 12'b010100000000;
		14'b00000100011000: color_data = 12'b010100000000;
		14'b00000100011001: color_data = 12'b010100000000;
		14'b00000100011010: color_data = 12'b010100000000;
		14'b00000100011011: color_data = 12'b010100000000;
		14'b00000100011100: color_data = 12'b010100000000;
		14'b00000101000001: color_data = 12'b010100000000;
		14'b00000101000010: color_data = 12'b010100000000;
		14'b00000101001111: color_data = 12'b010100000000;
		14'b00000101010000: color_data = 12'b101000000000;
		14'b00000101010001: color_data = 12'b101000000000;
		14'b00000101010010: color_data = 12'b101000000000;
		14'b00000101010011: color_data = 12'b101000000000;
		14'b00000101010100: color_data = 12'b101000000000;
		14'b00000101010101: color_data = 12'b101000000000;
		14'b00000101010110: color_data = 12'b101000000000;
		14'b00000101010111: color_data = 12'b101000000000;
		14'b00000101011000: color_data = 12'b101000000000;
		14'b00000101011001: color_data = 12'b010100000000;
		14'b00000110000011: color_data = 12'b010100000000;
		14'b00000110000100: color_data = 12'b010100000000;
		14'b00000110000101: color_data = 12'b010100000000;
		14'b00000110000110: color_data = 12'b010100000000;
		14'b00000110000111: color_data = 12'b010100000000;
		14'b00000110001000: color_data = 12'b010100000000;
		14'b00000110001001: color_data = 12'b010100000000;
		14'b00000110001010: color_data = 12'b010100000000;
		14'b00000110001011: color_data = 12'b010100000000;
		14'b00000110001100: color_data = 12'b010100000000;
		14'b00000110001101: color_data = 12'b010100000000;
		14'b00000110001110: color_data = 12'b010100000000;
		14'b00000110001111: color_data = 12'b010100000000;
		14'b00000110010000: color_data = 12'b010100000000;
		14'b00000110010001: color_data = 12'b010100000000;
		14'b00000110010010: color_data = 12'b101000000000;
		14'b00000110010011: color_data = 12'b010100000000;
		14'b00000110010100: color_data = 12'b010100000000;
		14'b00000110010101: color_data = 12'b010100000000;
		14'b00000110010110: color_data = 12'b010100000000;
		14'b00000110010111: color_data = 12'b010100000000;
		14'b00000110011000: color_data = 12'b010100000000;
		14'b00000110011001: color_data = 12'b010100000000;
		14'b00000110011010: color_data = 12'b010100000000;
		14'b00000110011011: color_data = 12'b010100000000;
		14'b00000110011100: color_data = 12'b010100000000;
		14'b00000110011101: color_data = 12'b010100000000;
		14'b00000111010000: color_data = 12'b010100000000;
		14'b00000111010001: color_data = 12'b101000000000;
		14'b00000111010010: color_data = 12'b101000000000;
		14'b00000111010011: color_data = 12'b101000000000;
		14'b00000111010100: color_data = 12'b101000000000;
		14'b00000111010101: color_data = 12'b101000000000;
		14'b00000111010110: color_data = 12'b101000000000;
		14'b00000111010111: color_data = 12'b101000000000;
		14'b00000111011000: color_data = 12'b010100000000;
		14'b00000111011111: color_data = 12'b010100000000;
		14'b00000111100000: color_data = 12'b010100000000;
		14'b00001000001000: color_data = 12'b010100000000;
		14'b00001000001001: color_data = 12'b010100000000;
		14'b00001000001010: color_data = 12'b010100000000;
		14'b00001000001011: color_data = 12'b010100000000;
		14'b00001000001100: color_data = 12'b010100000000;
		14'b00001000001101: color_data = 12'b101000000000;
		14'b00001000001110: color_data = 12'b010100000000;
		14'b00001000001111: color_data = 12'b010100000000;
		14'b00001000010000: color_data = 12'b010100000000;
		14'b00001000010001: color_data = 12'b101000000000;
		14'b00001000010010: color_data = 12'b101000000000;
		14'b00001000010011: color_data = 12'b101000000000;
		14'b00001000010100: color_data = 12'b101000000000;
		14'b00001000010101: color_data = 12'b101000000000;
		14'b00001000010110: color_data = 12'b101000000000;
		14'b00001000010111: color_data = 12'b101000000000;
		14'b00001000011000: color_data = 12'b101000000000;
		14'b00001000011001: color_data = 12'b101000000000;
		14'b00001000011010: color_data = 12'b010100000000;
		14'b00001000011011: color_data = 12'b010100000000;
		14'b00001000011100: color_data = 12'b010100000000;
		14'b00001000011101: color_data = 12'b010100000000;
		14'b00001000011110: color_data = 12'b010100000000;
		14'b00001001001111: color_data = 12'b010100000000;
		14'b00001001010000: color_data = 12'b101000000000;
		14'b00001001010001: color_data = 12'b101000000000;
		14'b00001001010010: color_data = 12'b101000000000;
		14'b00001001010011: color_data = 12'b101000000000;
		14'b00001001010100: color_data = 12'b101000000000;
		14'b00001001010101: color_data = 12'b101000000000;
		14'b00001001010110: color_data = 12'b101000000000;
		14'b00001001010111: color_data = 12'b101000000000;
		14'b00001001011000: color_data = 12'b010100000000;
		14'b00001001011101: color_data = 12'b010100000000;
		14'b00001001011110: color_data = 12'b101000000000;
		14'b00001001011111: color_data = 12'b010100000000;
		14'b00001010001000: color_data = 12'b010100000000;
		14'b00001010001001: color_data = 12'b010100000000;
		14'b00001010001010: color_data = 12'b010100000000;
		14'b00001010001011: color_data = 12'b101000000000;
		14'b00001010001100: color_data = 12'b101000000000;
		14'b00001010001101: color_data = 12'b101000000000;
		14'b00001010001110: color_data = 12'b101000000000;
		14'b00001010001111: color_data = 12'b010100000000;
		14'b00001010010000: color_data = 12'b101000000000;
		14'b00001010010001: color_data = 12'b101000000000;
		14'b00001010010010: color_data = 12'b101000000000;
		14'b00001010010011: color_data = 12'b101000000000;
		14'b00001010010100: color_data = 12'b101000000000;
		14'b00001010010101: color_data = 12'b101000000000;
		14'b00001010010110: color_data = 12'b101000000000;
		14'b00001010010111: color_data = 12'b101000000000;
		14'b00001010011000: color_data = 12'b101000000000;
		14'b00001010011001: color_data = 12'b101000000000;
		14'b00001010011010: color_data = 12'b101000000000;
		14'b00001010011011: color_data = 12'b101000000000;
		14'b00001010011100: color_data = 12'b101000000000;
		14'b00001010011101: color_data = 12'b101000000000;
		14'b00001010011110: color_data = 12'b010100000000;
		14'b00001010011111: color_data = 12'b010100000000;
		14'b00001010100000: color_data = 12'b010100000000;
		14'b00001011001110: color_data = 12'b010100000000;
		14'b00001011001111: color_data = 12'b101000000000;
		14'b00001011010000: color_data = 12'b101000000000;
		14'b00001011010001: color_data = 12'b101000000000;
		14'b00001011010010: color_data = 12'b101000000000;
		14'b00001011010011: color_data = 12'b101000000000;
		14'b00001011010100: color_data = 12'b101000000000;
		14'b00001011010101: color_data = 12'b101000000000;
		14'b00001011010110: color_data = 12'b101000000000;
		14'b00001011010111: color_data = 12'b010100000000;
		14'b00001011011011: color_data = 12'b010100000000;
		14'b00001011011100: color_data = 12'b101000000000;
		14'b00001011011101: color_data = 12'b101000000000;
		14'b00001011011110: color_data = 12'b010100000000;
		14'b00001100000111: color_data = 12'b010100000000;
		14'b00001100001000: color_data = 12'b101000000000;
		14'b00001100001001: color_data = 12'b101000000000;
		14'b00001100001010: color_data = 12'b101000000000;
		14'b00001100001011: color_data = 12'b101000000000;
		14'b00001100001100: color_data = 12'b101000000000;
		14'b00001100001101: color_data = 12'b101000000000;
		14'b00001100001110: color_data = 12'b101000000000;
		14'b00001100001111: color_data = 12'b101000000000;
		14'b00001100010000: color_data = 12'b101000000000;
		14'b00001100010001: color_data = 12'b101000000000;
		14'b00001100010010: color_data = 12'b101000000000;
		14'b00001100010011: color_data = 12'b101000000000;
		14'b00001100010100: color_data = 12'b101000000000;
		14'b00001100010101: color_data = 12'b101000000000;
		14'b00001100010110: color_data = 12'b101000000000;
		14'b00001100010111: color_data = 12'b101000000000;
		14'b00001100011000: color_data = 12'b101000000000;
		14'b00001100011001: color_data = 12'b101000000000;
		14'b00001100011010: color_data = 12'b101000000000;
		14'b00001100011011: color_data = 12'b101000000000;
		14'b00001100011100: color_data = 12'b101000000000;
		14'b00001100011101: color_data = 12'b101000000000;
		14'b00001100011110: color_data = 12'b101000000000;
		14'b00001100011111: color_data = 12'b101000000000;
		14'b00001100100000: color_data = 12'b101000000000;
		14'b00001100100001: color_data = 12'b010100000000;
		14'b00001101001101: color_data = 12'b010100000000;
		14'b00001101001110: color_data = 12'b101000000000;
		14'b00001101001111: color_data = 12'b101000000000;
		14'b00001101010000: color_data = 12'b101000000000;
		14'b00001101010001: color_data = 12'b101000000000;
		14'b00001101010010: color_data = 12'b101000000000;
		14'b00001101010011: color_data = 12'b101000000000;
		14'b00001101010100: color_data = 12'b101000000000;
		14'b00001101010101: color_data = 12'b101000000000;
		14'b00001101010110: color_data = 12'b101000000000;
		14'b00001101010111: color_data = 12'b010100000000;
		14'b00001101011010: color_data = 12'b010100000000;
		14'b00001101011011: color_data = 12'b010100000000;
		14'b00001101011100: color_data = 12'b101000000000;
		14'b00001101011101: color_data = 12'b010100000000;
		14'b00001110000110: color_data = 12'b010100000000;
		14'b00001110000111: color_data = 12'b101000000000;
		14'b00001110001000: color_data = 12'b101000000000;
		14'b00001110001001: color_data = 12'b101000000000;
		14'b00001110001010: color_data = 12'b101000000000;
		14'b00001110001011: color_data = 12'b101000000000;
		14'b00001110001100: color_data = 12'b101000000000;
		14'b00001110001101: color_data = 12'b101000000000;
		14'b00001110001110: color_data = 12'b101000000000;
		14'b00001110001111: color_data = 12'b101000000000;
		14'b00001110010000: color_data = 12'b101000000000;
		14'b00001110010001: color_data = 12'b101000000000;
		14'b00001110010010: color_data = 12'b010100000000;
		14'b00001110010011: color_data = 12'b010100000000;
		14'b00001110010100: color_data = 12'b010100000000;
		14'b00001110010101: color_data = 12'b010100000000;
		14'b00001110010110: color_data = 12'b101000000000;
		14'b00001110010111: color_data = 12'b101000000000;
		14'b00001110011000: color_data = 12'b101000000000;
		14'b00001110011001: color_data = 12'b010100000000;
		14'b00001110011010: color_data = 12'b010100000000;
		14'b00001110011011: color_data = 12'b010100000000;
		14'b00001110011100: color_data = 12'b010100000000;
		14'b00001110011101: color_data = 12'b010100000000;
		14'b00001110011110: color_data = 12'b101000000000;
		14'b00001110011111: color_data = 12'b101000000000;
		14'b00001110100000: color_data = 12'b101000000000;
		14'b00001110100001: color_data = 12'b101000000000;
		14'b00001110100010: color_data = 12'b101000000000;
		14'b00001110100011: color_data = 12'b010100000000;
		14'b00001111001110: color_data = 12'b101000000000;
		14'b00001111001111: color_data = 12'b101000000000;
		14'b00001111010000: color_data = 12'b101000000000;
		14'b00001111010001: color_data = 12'b101000000000;
		14'b00001111010010: color_data = 12'b101000000000;
		14'b00001111010011: color_data = 12'b101000000000;
		14'b00001111010100: color_data = 12'b101000000000;
		14'b00001111010101: color_data = 12'b101000000000;
		14'b00001111010110: color_data = 12'b101000000000;
		14'b00001111010111: color_data = 12'b101000000000;
		14'b00001111011000: color_data = 12'b010100000000;
		14'b00001111011001: color_data = 12'b010100000000;
		14'b00001111011010: color_data = 12'b010100000000;
		14'b00001111011011: color_data = 12'b101000000000;
		14'b00001111011100: color_data = 12'b010100000000;
		14'b00010000000101: color_data = 12'b010100000000;
		14'b00010000000110: color_data = 12'b010100000000;
		14'b00010000000111: color_data = 12'b010100000000;
		14'b00010000001000: color_data = 12'b010100000000;
		14'b00010000001001: color_data = 12'b010100000000;
		14'b00010000001010: color_data = 12'b010100000000;
		14'b00010000001011: color_data = 12'b010100000000;
		14'b00010000001100: color_data = 12'b101000000000;
		14'b00010000001101: color_data = 12'b101000000000;
		14'b00010000001110: color_data = 12'b101000000000;
		14'b00010000001111: color_data = 12'b101000000000;
		14'b00010000010000: color_data = 12'b010100000000;
		14'b00010000010001: color_data = 12'b010100000000;
		14'b00010000010111: color_data = 12'b010100000000;
		14'b00010000011000: color_data = 12'b101000000000;
		14'b00010000011001: color_data = 12'b101000000000;
		14'b00010000011010: color_data = 12'b010100000000;
		14'b00010000011011: color_data = 12'b010100000000;
		14'b00010000011111: color_data = 12'b010100000000;
		14'b00010000100000: color_data = 12'b010100000000;
		14'b00010000100001: color_data = 12'b101000000000;
		14'b00010000100010: color_data = 12'b101000000000;
		14'b00010000100011: color_data = 12'b101000000000;
		14'b00010000100100: color_data = 12'b010100000000;
		14'b00010000100101: color_data = 12'b010100000000;
		14'b00010001001110: color_data = 12'b101000000000;
		14'b00010001001111: color_data = 12'b101000000000;
		14'b00010001010000: color_data = 12'b101000000000;
		14'b00010001010001: color_data = 12'b101000000000;
		14'b00010001010010: color_data = 12'b101000000000;
		14'b00010001010011: color_data = 12'b101000000000;
		14'b00010001010100: color_data = 12'b101000000000;
		14'b00010001010101: color_data = 12'b101000000000;
		14'b00010001010110: color_data = 12'b101000000000;
		14'b00010001010111: color_data = 12'b101000000000;
		14'b00010001011000: color_data = 12'b010100000000;
		14'b00010001011001: color_data = 12'b010100000000;
		14'b00010001011010: color_data = 12'b101000000000;
		14'b00010001011011: color_data = 12'b101000000000;
		14'b00010010000101: color_data = 12'b010100000000;
		14'b00010010000110: color_data = 12'b010100000000;
		14'b00010010001001: color_data = 12'b010100000000;
		14'b00010010001010: color_data = 12'b010100000000;
		14'b00010010001011: color_data = 12'b010100000000;
		14'b00010010001100: color_data = 12'b101000000000;
		14'b00010010001101: color_data = 12'b101000000000;
		14'b00010010001110: color_data = 12'b101000000000;
		14'b00010010001111: color_data = 12'b010100000000;
		14'b00010010010111: color_data = 12'b010100000000;
		14'b00010010011000: color_data = 12'b101000000000;
		14'b00010010011001: color_data = 12'b101000000000;
		14'b00010010011010: color_data = 12'b101000000000;
		14'b00010010011011: color_data = 12'b101000000000;
		14'b00010010011100: color_data = 12'b010100000000;
		14'b00010010011101: color_data = 12'b010100000000;
		14'b00010010100010: color_data = 12'b010100000000;
		14'b00010010100011: color_data = 12'b101000000000;
		14'b00010010100100: color_data = 12'b101000000000;
		14'b00010010100101: color_data = 12'b101000000000;
		14'b00010010100110: color_data = 12'b010100000000;
		14'b00010010100111: color_data = 12'b010100000000;
		14'b00010011000110: color_data = 12'b010100000000;
		14'b00010011001110: color_data = 12'b101000000000;
		14'b00010011001111: color_data = 12'b101000000000;
		14'b00010011010000: color_data = 12'b101000000000;
		14'b00010011010001: color_data = 12'b101000000000;
		14'b00010011010010: color_data = 12'b101000000000;
		14'b00010011010011: color_data = 12'b101000000000;
		14'b00010011010100: color_data = 12'b101000000000;
		14'b00010011010101: color_data = 12'b101000000000;
		14'b00010011010110: color_data = 12'b101000000000;
		14'b00010011010111: color_data = 12'b101000000000;
		14'b00010011011000: color_data = 12'b010100000000;
		14'b00010011011001: color_data = 12'b010100000000;
		14'b00010011011010: color_data = 12'b101000000000;
		14'b00010011011011: color_data = 12'b010100000000;
		14'b00010100000100: color_data = 12'b010100000000;
		14'b00010100000101: color_data = 12'b010100000000;
		14'b00010100001001: color_data = 12'b010100000000;
		14'b00010100001010: color_data = 12'b010100000000;
		14'b00010100001011: color_data = 12'b101000000000;
		14'b00010100001100: color_data = 12'b101000000000;
		14'b00010100001101: color_data = 12'b010100000000;
		14'b00010100001110: color_data = 12'b010100000000;
		14'b00010100010100: color_data = 12'b010100000000;
		14'b00010100010101: color_data = 12'b010100000000;
		14'b00010100010110: color_data = 12'b010100000000;
		14'b00010100010111: color_data = 12'b101000000000;
		14'b00010100011000: color_data = 12'b101000000000;
		14'b00010100011001: color_data = 12'b101000000000;
		14'b00010100011010: color_data = 12'b101000000000;
		14'b00010100011011: color_data = 12'b101000000000;
		14'b00010100011100: color_data = 12'b101000000000;
		14'b00010100011101: color_data = 12'b101000000000;
		14'b00010100011110: color_data = 12'b101000000000;
		14'b00010100011111: color_data = 12'b010100000000;
		14'b00010100100100: color_data = 12'b010100000000;
		14'b00010100100101: color_data = 12'b101000000000;
		14'b00010100100110: color_data = 12'b010100000000;
		14'b00010100100111: color_data = 12'b010100000000;
		14'b00010100101000: color_data = 12'b010100000000;
		14'b00010101001101: color_data = 12'b010100000000;
		14'b00010101001110: color_data = 12'b101000000000;
		14'b00010101001111: color_data = 12'b101000000000;
		14'b00010101010000: color_data = 12'b101000000000;
		14'b00010101010001: color_data = 12'b101000000000;
		14'b00010101010010: color_data = 12'b101000000000;
		14'b00010101010011: color_data = 12'b101000000000;
		14'b00010101010100: color_data = 12'b101000000000;
		14'b00010101010101: color_data = 12'b101000000000;
		14'b00010101010110: color_data = 12'b101000000000;
		14'b00010101010111: color_data = 12'b010100000000;
		14'b00010101011000: color_data = 12'b010100000000;
		14'b00010101011001: color_data = 12'b101000000000;
		14'b00010101011010: color_data = 12'b101000000000;
		14'b00010110001000: color_data = 12'b010100000000;
		14'b00010110001001: color_data = 12'b010100000000;
		14'b00010110001010: color_data = 12'b010100000000;
		14'b00010110001011: color_data = 12'b010100000000;
		14'b00010110001100: color_data = 12'b010100000000;
		14'b00010110001101: color_data = 12'b010100000000;
		14'b00010110001110: color_data = 12'b010100000000;
		14'b00010110001111: color_data = 12'b010100000000;
		14'b00010110010000: color_data = 12'b010100000000;
		14'b00010110010001: color_data = 12'b101000000000;
		14'b00010110010010: color_data = 12'b101000000000;
		14'b00010110010011: color_data = 12'b101000000000;
		14'b00010110010100: color_data = 12'b101000000000;
		14'b00010110010101: color_data = 12'b101000000000;
		14'b00010110010110: color_data = 12'b101000000000;
		14'b00010110010111: color_data = 12'b101000000000;
		14'b00010110011000: color_data = 12'b101000000000;
		14'b00010110011001: color_data = 12'b101000000000;
		14'b00010110011010: color_data = 12'b101000000000;
		14'b00010110011011: color_data = 12'b101000000000;
		14'b00010110011100: color_data = 12'b101000000000;
		14'b00010110011101: color_data = 12'b101000000000;
		14'b00010110011110: color_data = 12'b101000000000;
		14'b00010110011111: color_data = 12'b101000000000;
		14'b00010110100000: color_data = 12'b101000000000;
		14'b00010110100001: color_data = 12'b010100000000;
		14'b00010110100010: color_data = 12'b010100000000;
		14'b00010110100110: color_data = 12'b010100000000;
		14'b00010110100111: color_data = 12'b010100000000;
		14'b00010110101000: color_data = 12'b010100000000;
		14'b00010110101001: color_data = 12'b010100000000;
		14'b00010111001101: color_data = 12'b010100000000;
		14'b00010111001110: color_data = 12'b101000000000;
		14'b00010111001111: color_data = 12'b101000000000;
		14'b00010111010000: color_data = 12'b101000000000;
		14'b00010111010001: color_data = 12'b101000000000;
		14'b00010111010010: color_data = 12'b101000000000;
		14'b00010111010011: color_data = 12'b101000000000;
		14'b00010111010100: color_data = 12'b101000000000;
		14'b00010111010101: color_data = 12'b101000000000;
		14'b00010111010110: color_data = 12'b101000000000;
		14'b00010111010111: color_data = 12'b010100000000;
		14'b00010111011000: color_data = 12'b010100000000;
		14'b00010111011001: color_data = 12'b101000000000;
		14'b00010111011010: color_data = 12'b010100000000;
		14'b00011000001000: color_data = 12'b010100000000;
		14'b00011000001100: color_data = 12'b010100000000;
		14'b00011000001101: color_data = 12'b010100000000;
		14'b00011000001110: color_data = 12'b101000000000;
		14'b00011000001111: color_data = 12'b101000000000;
		14'b00011000010000: color_data = 12'b101000000000;
		14'b00011000010001: color_data = 12'b101000000000;
		14'b00011000010010: color_data = 12'b101000000000;
		14'b00011000010011: color_data = 12'b101000000000;
		14'b00011000010100: color_data = 12'b101000000000;
		14'b00011000010101: color_data = 12'b101000000000;
		14'b00011000010110: color_data = 12'b101000000000;
		14'b00011000010111: color_data = 12'b101000000000;
		14'b00011000011000: color_data = 12'b101000000000;
		14'b00011000011001: color_data = 12'b101000000000;
		14'b00011000011010: color_data = 12'b101000000000;
		14'b00011000011011: color_data = 12'b101000000000;
		14'b00011000011100: color_data = 12'b101000000000;
		14'b00011000011101: color_data = 12'b101000000000;
		14'b00011000011110: color_data = 12'b101000000000;
		14'b00011000011111: color_data = 12'b101000000000;
		14'b00011000100000: color_data = 12'b101000000000;
		14'b00011000100001: color_data = 12'b101000000000;
		14'b00011000100010: color_data = 12'b101000000000;
		14'b00011000100011: color_data = 12'b010100000000;
		14'b00011000100100: color_data = 12'b010100000000;
		14'b00011000100111: color_data = 12'b010100000000;
		14'b00011000101000: color_data = 12'b010100000000;
		14'b00011000101001: color_data = 12'b010100000000;
		14'b00011001001101: color_data = 12'b101000000000;
		14'b00011001001110: color_data = 12'b101000000000;
		14'b00011001001111: color_data = 12'b101000000000;
		14'b00011001010000: color_data = 12'b101000000000;
		14'b00011001010001: color_data = 12'b101000000000;
		14'b00011001010010: color_data = 12'b101000000000;
		14'b00011001010011: color_data = 12'b101000000000;
		14'b00011001010100: color_data = 12'b101000000000;
		14'b00011001010101: color_data = 12'b101000000000;
		14'b00011001010110: color_data = 12'b010100000000;
		14'b00011001010111: color_data = 12'b010100000000;
		14'b00011001011000: color_data = 12'b101000000000;
		14'b00011001011001: color_data = 12'b101000000000;
		14'b00011010001101: color_data = 12'b010100000000;
		14'b00011010001110: color_data = 12'b101000000000;
		14'b00011010001111: color_data = 12'b101000000000;
		14'b00011010010000: color_data = 12'b101000000000;
		14'b00011010010001: color_data = 12'b010100000000;
		14'b00011010010010: color_data = 12'b010100000000;
		14'b00011010010011: color_data = 12'b010100000000;
		14'b00011010010100: color_data = 12'b010100000000;
		14'b00011010010101: color_data = 12'b010100000000;
		14'b00011010010110: color_data = 12'b101000000000;
		14'b00011010010111: color_data = 12'b101000000000;
		14'b00011010011000: color_data = 12'b101000000000;
		14'b00011010011001: color_data = 12'b101000000000;
		14'b00011010011010: color_data = 12'b101000000000;
		14'b00011010011011: color_data = 12'b101000000000;
		14'b00011010011100: color_data = 12'b101000000000;
		14'b00011010011101: color_data = 12'b010100000000;
		14'b00011010011110: color_data = 12'b010100000000;
		14'b00011010011111: color_data = 12'b101000000000;
		14'b00011010100000: color_data = 12'b101000000000;
		14'b00011010100001: color_data = 12'b101000000000;
		14'b00011010100010: color_data = 12'b101000000000;
		14'b00011010100011: color_data = 12'b101000000000;
		14'b00011010100100: color_data = 12'b101000000000;
		14'b00011010100101: color_data = 12'b101000000000;
		14'b00011010100110: color_data = 12'b010100000000;
		14'b00011010100111: color_data = 12'b010100000000;
		14'b00011010101000: color_data = 12'b010100000000;
		14'b00011010101001: color_data = 12'b010100000000;
		14'b00011010101010: color_data = 12'b010100000000;
		14'b00011010101011: color_data = 12'b010100000000;
		14'b00011011001101: color_data = 12'b101000000000;
		14'b00011011001110: color_data = 12'b101000000000;
		14'b00011011001111: color_data = 12'b101000000000;
		14'b00011011010000: color_data = 12'b101000000000;
		14'b00011011010001: color_data = 12'b101000000000;
		14'b00011011010010: color_data = 12'b101000000000;
		14'b00011011010011: color_data = 12'b101000000000;
		14'b00011011010100: color_data = 12'b101000000000;
		14'b00011011010101: color_data = 12'b101000000000;
		14'b00011011010110: color_data = 12'b010100000000;
		14'b00011011010111: color_data = 12'b010100000000;
		14'b00011011011000: color_data = 12'b101000000000;
		14'b00011011011001: color_data = 12'b010100000000;
		14'b00011100001100: color_data = 12'b010100000000;
		14'b00011100001101: color_data = 12'b010100000000;
		14'b00011100010011: color_data = 12'b010100000000;
		14'b00011100010100: color_data = 12'b010100000000;
		14'b00011100010101: color_data = 12'b101000000000;
		14'b00011100010110: color_data = 12'b101000000000;
		14'b00011100010111: color_data = 12'b101000000000;
		14'b00011100011000: color_data = 12'b101000000000;
		14'b00011100011001: color_data = 12'b101000000000;
		14'b00011100011010: color_data = 12'b010100000000;
		14'b00011100011011: color_data = 12'b010100000000;
		14'b00011100011111: color_data = 12'b010100000000;
		14'b00011100100000: color_data = 12'b101000000000;
		14'b00011100100001: color_data = 12'b010100000000;
		14'b00011100100010: color_data = 12'b010100000000;
		14'b00011100100011: color_data = 12'b101000000000;
		14'b00011100100100: color_data = 12'b101000000000;
		14'b00011100100101: color_data = 12'b101000000000;
		14'b00011100100110: color_data = 12'b101000000000;
		14'b00011100100111: color_data = 12'b101000000000;
		14'b00011100101000: color_data = 12'b010100000000;
		14'b00011100101001: color_data = 12'b010100000000;
		14'b00011100101010: color_data = 12'b010100000000;
		14'b00011100101011: color_data = 12'b101000000000;
		14'b00011100101100: color_data = 12'b010100000000;
		14'b00011101001100: color_data = 12'b010100000000;
		14'b00011101001101: color_data = 12'b101000000000;
		14'b00011101001110: color_data = 12'b101000000000;
		14'b00011101001111: color_data = 12'b101000000000;
		14'b00011101010000: color_data = 12'b101000000000;
		14'b00011101010001: color_data = 12'b101000000000;
		14'b00011101010010: color_data = 12'b101000000000;
		14'b00011101010011: color_data = 12'b101000000000;
		14'b00011101010100: color_data = 12'b101000000000;
		14'b00011101010101: color_data = 12'b101000000000;
		14'b00011101010110: color_data = 12'b010100000000;
		14'b00011101010111: color_data = 12'b101000000000;
		14'b00011101011000: color_data = 12'b101000000000;
		14'b00011110010010: color_data = 12'b010100000000;
		14'b00011110010011: color_data = 12'b010100000000;
		14'b00011110010100: color_data = 12'b101000000000;
		14'b00011110010101: color_data = 12'b101000000000;
		14'b00011110010110: color_data = 12'b101000000000;
		14'b00011110010111: color_data = 12'b101000000000;
		14'b00011110011000: color_data = 12'b010100000000;
		14'b00011110011001: color_data = 12'b010100000000;
		14'b00011110011110: color_data = 12'b010100000000;
		14'b00011110011111: color_data = 12'b010100000000;
		14'b00011110100000: color_data = 12'b101000000000;
		14'b00011110100001: color_data = 12'b101000000000;
		14'b00011110100010: color_data = 12'b010100000000;
		14'b00011110100100: color_data = 12'b010100000000;
		14'b00011110100101: color_data = 12'b101000000000;
		14'b00011110100110: color_data = 12'b101000000000;
		14'b00011110100111: color_data = 12'b101000000000;
		14'b00011110101000: color_data = 12'b101000000000;
		14'b00011110101001: color_data = 12'b101000000000;
		14'b00011110101010: color_data = 12'b010100000000;
		14'b00011110101011: color_data = 12'b010100000000;
		14'b00011110101100: color_data = 12'b010100000000;
		14'b00011110101101: color_data = 12'b010100000000;
		14'b00011111001101: color_data = 12'b101000000000;
		14'b00011111001110: color_data = 12'b101000000000;
		14'b00011111001111: color_data = 12'b101000000000;
		14'b00011111010000: color_data = 12'b101000000000;
		14'b00011111010001: color_data = 12'b101000000000;
		14'b00011111010010: color_data = 12'b101000000000;
		14'b00011111010011: color_data = 12'b101000000000;
		14'b00011111010100: color_data = 12'b101000000000;
		14'b00011111010101: color_data = 12'b010100000000;
		14'b00011111010110: color_data = 12'b010100000000;
		14'b00011111010111: color_data = 12'b101000000000;
		14'b00011111011000: color_data = 12'b010100000000;
		14'b00100000010000: color_data = 12'b010100000000;
		14'b00100000010001: color_data = 12'b010100000000;
		14'b00100000010010: color_data = 12'b101000000000;
		14'b00100000010011: color_data = 12'b101000000000;
		14'b00100000010100: color_data = 12'b101000000000;
		14'b00100000010101: color_data = 12'b101000000000;
		14'b00100000010110: color_data = 12'b101000000000;
		14'b00100000010111: color_data = 12'b101000000000;
		14'b00100000011000: color_data = 12'b010100000000;
		14'b00100000011001: color_data = 12'b010100000000;
		14'b00100000011010: color_data = 12'b010100000000;
		14'b00100000011011: color_data = 12'b010100000000;
		14'b00100000011100: color_data = 12'b010100000000;
		14'b00100000011101: color_data = 12'b010100000000;
		14'b00100000011110: color_data = 12'b101000000000;
		14'b00100000011111: color_data = 12'b101000000000;
		14'b00100000100000: color_data = 12'b101000000000;
		14'b00100000100001: color_data = 12'b101000000000;
		14'b00100000100010: color_data = 12'b101000000000;
		14'b00100000100011: color_data = 12'b010100000000;
		14'b00100000100100: color_data = 12'b010100000000;
		14'b00100000100101: color_data = 12'b010100000000;
		14'b00100000100110: color_data = 12'b101000000000;
		14'b00100000100111: color_data = 12'b101000000000;
		14'b00100000101000: color_data = 12'b101000000000;
		14'b00100000101001: color_data = 12'b101000000000;
		14'b00100000101010: color_data = 12'b101000000000;
		14'b00100000101011: color_data = 12'b010100000000;
		14'b00100000101100: color_data = 12'b010100000000;
		14'b00100000101101: color_data = 12'b010100000000;
		14'b00100001001101: color_data = 12'b010100000000;
		14'b00100001001110: color_data = 12'b101000000000;
		14'b00100001001111: color_data = 12'b101000000000;
		14'b00100001010000: color_data = 12'b101000000000;
		14'b00100001010001: color_data = 12'b101000000000;
		14'b00100001010010: color_data = 12'b101000000000;
		14'b00100001010011: color_data = 12'b101000000000;
		14'b00100001010100: color_data = 12'b010100000000;
		14'b00100001010101: color_data = 12'b010100000000;
		14'b00100001010110: color_data = 12'b101000000000;
		14'b00100001010111: color_data = 12'b101000000000;
		14'b00100010001110: color_data = 12'b010100000000;
		14'b00100010001111: color_data = 12'b010100000000;
		14'b00100010010000: color_data = 12'b101000000000;
		14'b00100010010001: color_data = 12'b101000000000;
		14'b00100010010010: color_data = 12'b101000000000;
		14'b00100010010011: color_data = 12'b101000000000;
		14'b00100010010100: color_data = 12'b101000000000;
		14'b00100010010101: color_data = 12'b101000000000;
		14'b00100010010110: color_data = 12'b101000000000;
		14'b00100010010111: color_data = 12'b101000000000;
		14'b00100010011000: color_data = 12'b101000000000;
		14'b00100010011001: color_data = 12'b101000000000;
		14'b00100010011010: color_data = 12'b101000000000;
		14'b00100010011011: color_data = 12'b101000000000;
		14'b00100010011100: color_data = 12'b010100000000;
		14'b00100010011101: color_data = 12'b010100000000;
		14'b00100010011110: color_data = 12'b010100000000;
		14'b00100010011111: color_data = 12'b010100000000;
		14'b00100010100000: color_data = 12'b101000000000;
		14'b00100010100001: color_data = 12'b101000000000;
		14'b00100010100010: color_data = 12'b101000000000;
		14'b00100010100011: color_data = 12'b101000000000;
		14'b00100010100100: color_data = 12'b101000000000;
		14'b00100010100101: color_data = 12'b101000000000;
		14'b00100010100110: color_data = 12'b101000000000;
		14'b00100010100111: color_data = 12'b101000000000;
		14'b00100010101000: color_data = 12'b101000000000;
		14'b00100010101001: color_data = 12'b101000000000;
		14'b00100010101010: color_data = 12'b101000000000;
		14'b00100010101011: color_data = 12'b101000000000;
		14'b00100010101100: color_data = 12'b010100000000;
		14'b00100010101101: color_data = 12'b010100000000;
		14'b00100011001101: color_data = 12'b010100000000;
		14'b00100011001110: color_data = 12'b101000000000;
		14'b00100011001111: color_data = 12'b101000000000;
		14'b00100011010000: color_data = 12'b101000000000;
		14'b00100011010001: color_data = 12'b101000000000;
		14'b00100011010010: color_data = 12'b101000000000;
		14'b00100011010011: color_data = 12'b101000000000;
		14'b00100011010100: color_data = 12'b010100000000;
		14'b00100011010101: color_data = 12'b101000000000;
		14'b00100011010110: color_data = 12'b101000000000;
		14'b00100011010111: color_data = 12'b010100000000;
		14'b00100100001101: color_data = 12'b010100000000;
		14'b00100100001110: color_data = 12'b010100000000;
		14'b00100100001111: color_data = 12'b101000000000;
		14'b00100100010000: color_data = 12'b101000000000;
		14'b00100100010001: color_data = 12'b101000000000;
		14'b00100100010010: color_data = 12'b101000000000;
		14'b00100100010011: color_data = 12'b101000000000;
		14'b00100100010100: color_data = 12'b101000000000;
		14'b00100100010101: color_data = 12'b101000000000;
		14'b00100100010110: color_data = 12'b101000000000;
		14'b00100100010111: color_data = 12'b010100000000;
		14'b00100100011000: color_data = 12'b010100000000;
		14'b00100100011001: color_data = 12'b010100000000;
		14'b00100100011010: color_data = 12'b010100000000;
		14'b00100100011011: color_data = 12'b010100000000;
		14'b00100100011111: color_data = 12'b010100000000;
		14'b00100100100000: color_data = 12'b010100000000;
		14'b00100100100001: color_data = 12'b101000000000;
		14'b00100100100010: color_data = 12'b101000000000;
		14'b00100100100011: color_data = 12'b101000000000;
		14'b00100100100100: color_data = 12'b101000000000;
		14'b00100100100101: color_data = 12'b101000000000;
		14'b00100100100110: color_data = 12'b101000000000;
		14'b00100100100111: color_data = 12'b101000000000;
		14'b00100100101000: color_data = 12'b101000000000;
		14'b00100100101001: color_data = 12'b101000000000;
		14'b00100100101010: color_data = 12'b010100000000;
		14'b00100100101011: color_data = 12'b010100000000;
		14'b00100100101100: color_data = 12'b101000000000;
		14'b00100100101101: color_data = 12'b010100000000;
		14'b00100101001100: color_data = 12'b010100000000;
		14'b00100101001101: color_data = 12'b101000000000;
		14'b00100101001110: color_data = 12'b101000000000;
		14'b00100101001111: color_data = 12'b101000000000;
		14'b00100101010000: color_data = 12'b101000000000;
		14'b00100101010001: color_data = 12'b101000000000;
		14'b00100101010010: color_data = 12'b101000000000;
		14'b00100101010011: color_data = 12'b010100000000;
		14'b00100101010100: color_data = 12'b010100000000;
		14'b00100101010101: color_data = 12'b101000000000;
		14'b00100101010110: color_data = 12'b101000000000;
		14'b00100101010111: color_data = 12'b010100000000;
		14'b00100110001100: color_data = 12'b010100000000;
		14'b00100110001101: color_data = 12'b010100000000;
		14'b00100110001110: color_data = 12'b101000000000;
		14'b00100110001111: color_data = 12'b101000000000;
		14'b00100110010000: color_data = 12'b101000000000;
		14'b00100110010001: color_data = 12'b101000000000;
		14'b00100110010010: color_data = 12'b101000000000;
		14'b00100110010011: color_data = 12'b101000000000;
		14'b00100110010100: color_data = 12'b010100000000;
		14'b00100110010101: color_data = 12'b010100000000;
		14'b00100110100000: color_data = 12'b010100000000;
		14'b00100110100001: color_data = 12'b010100000000;
		14'b00100110100010: color_data = 12'b101000000000;
		14'b00100110100011: color_data = 12'b101000000000;
		14'b00100110100100: color_data = 12'b101000000000;
		14'b00100110100101: color_data = 12'b101000000000;
		14'b00100110100110: color_data = 12'b101000000000;
		14'b00100110100111: color_data = 12'b101000000000;
		14'b00100110101000: color_data = 12'b101000000000;
		14'b00100110101001: color_data = 12'b101000000000;
		14'b00100110101010: color_data = 12'b010100000000;
		14'b00100110101011: color_data = 12'b010100000000;
		14'b00100110101100: color_data = 12'b010100000000;
		14'b00100110101101: color_data = 12'b101000000000;
		14'b00100110101110: color_data = 12'b010100000000;
		14'b00100111001100: color_data = 12'b010100000000;
		14'b00100111001101: color_data = 12'b101000000000;
		14'b00100111001110: color_data = 12'b101000000000;
		14'b00100111001111: color_data = 12'b101000000000;
		14'b00100111010000: color_data = 12'b101000000000;
		14'b00100111010001: color_data = 12'b101000000000;
		14'b00100111010010: color_data = 12'b010100000000;
		14'b00100111010011: color_data = 12'b010100000000;
		14'b00100111010100: color_data = 12'b101000000000;
		14'b00100111010101: color_data = 12'b101000000000;
		14'b00100111010110: color_data = 12'b101000000000;
		14'b00101000001011: color_data = 12'b010100000000;
		14'b00101000001100: color_data = 12'b010100000000;
		14'b00101000001101: color_data = 12'b101000000000;
		14'b00101000001110: color_data = 12'b101000000000;
		14'b00101000001111: color_data = 12'b101000000000;
		14'b00101000010000: color_data = 12'b010100000000;
		14'b00101000010001: color_data = 12'b010100000000;
		14'b00101000100000: color_data = 12'b010100000000;
		14'b00101000100001: color_data = 12'b010100000000;
		14'b00101000100010: color_data = 12'b010100000000;
		14'b00101000100011: color_data = 12'b101000000000;
		14'b00101000100100: color_data = 12'b101000000000;
		14'b00101000100101: color_data = 12'b010100000000;
		14'b00101000100110: color_data = 12'b010100000000;
		14'b00101000100111: color_data = 12'b010100000000;
		14'b00101000101000: color_data = 12'b010100000000;
		14'b00101000101001: color_data = 12'b101000000000;
		14'b00101000101010: color_data = 12'b101000000000;
		14'b00101000101011: color_data = 12'b010100000000;
		14'b00101000101101: color_data = 12'b010100000000;
		14'b00101000101110: color_data = 12'b010100000000;
		14'b00101001001100: color_data = 12'b010100000000;
		14'b00101001001101: color_data = 12'b101000000000;
		14'b00101001001110: color_data = 12'b101000000000;
		14'b00101001001111: color_data = 12'b101000000000;
		14'b00101001010000: color_data = 12'b101000000000;
		14'b00101001010001: color_data = 12'b101000000000;
		14'b00101001010010: color_data = 12'b010100000000;
		14'b00101001010011: color_data = 12'b010100000000;
		14'b00101001010100: color_data = 12'b101000000000;
		14'b00101001010101: color_data = 12'b101000000000;
		14'b00101001010110: color_data = 12'b010100000000;
		14'b00101010001001: color_data = 12'b010100000000;
		14'b00101010001010: color_data = 12'b010100000000;
		14'b00101010001011: color_data = 12'b010100000000;
		14'b00101010001100: color_data = 12'b101000000000;
		14'b00101010001101: color_data = 12'b101000000000;
		14'b00101010001110: color_data = 12'b010100000000;
		14'b00101010001111: color_data = 12'b010100000000;
		14'b00101010100001: color_data = 12'b010100000000;
		14'b00101010100010: color_data = 12'b010100000000;
		14'b00101010100011: color_data = 12'b010100000000;
		14'b00101010100100: color_data = 12'b010100000000;
		14'b00101010100101: color_data = 12'b010100000000;
		14'b00101010100110: color_data = 12'b010100000000;
		14'b00101010100111: color_data = 12'b010100000000;
		14'b00101010101000: color_data = 12'b010100000000;
		14'b00101010101001: color_data = 12'b010100000000;
		14'b00101010101010: color_data = 12'b101000000000;
		14'b00101010101011: color_data = 12'b010100000000;
		14'b00101010101110: color_data = 12'b010100000000;
		14'b00101010101111: color_data = 12'b010100000000;
		14'b00101011001100: color_data = 12'b101000000000;
		14'b00101011001101: color_data = 12'b101000000000;
		14'b00101011001110: color_data = 12'b101000000000;
		14'b00101011001111: color_data = 12'b101000000000;
		14'b00101011010000: color_data = 12'b101000000000;
		14'b00101011010001: color_data = 12'b010100000000;
		14'b00101011010010: color_data = 12'b010100000000;
		14'b00101011010011: color_data = 12'b101000000000;
		14'b00101011010100: color_data = 12'b101000000000;
		14'b00101011010101: color_data = 12'b101000000000;
		14'b00101011010111: color_data = 12'b010100000000;
		14'b00101011101001: color_data = 12'b010100000000;
		14'b00101011101010: color_data = 12'b010100000000;
		14'b00101100001000: color_data = 12'b010100000000;
		14'b00101100001001: color_data = 12'b010100000000;
		14'b00101100001010: color_data = 12'b010100000000;
		14'b00101100001011: color_data = 12'b101000000000;
		14'b00101100001100: color_data = 12'b101000000000;
		14'b00101100001101: color_data = 12'b101000000000;
		14'b00101100001110: color_data = 12'b010100000000;
		14'b00101100011101: color_data = 12'b010100000000;
		14'b00101100011110: color_data = 12'b010100000000;
		14'b00101100100011: color_data = 12'b010100000000;
		14'b00101100101000: color_data = 12'b010100000000;
		14'b00101100101001: color_data = 12'b010100000000;
		14'b00101100101010: color_data = 12'b101000000000;
		14'b00101100101011: color_data = 12'b010100000000;
		14'b00101100101111: color_data = 12'b010100000000;
		14'b00101101001011: color_data = 12'b010100000000;
		14'b00101101001100: color_data = 12'b101000000000;
		14'b00101101001101: color_data = 12'b101000000000;
		14'b00101101001110: color_data = 12'b101000000000;
		14'b00101101001111: color_data = 12'b101000000000;
		14'b00101101010000: color_data = 12'b010100000000;
		14'b00101101010001: color_data = 12'b010100000000;
		14'b00101101010010: color_data = 12'b101000000000;
		14'b00101101010011: color_data = 12'b101000000000;
		14'b00101101010100: color_data = 12'b101000000000;
		14'b00101101010101: color_data = 12'b101000000000;
		14'b00101101010110: color_data = 12'b010100000000;
		14'b00101101010111: color_data = 12'b010100000000;
		14'b00101101101001: color_data = 12'b010100000000;
		14'b00101101101010: color_data = 12'b010100000000;
		14'b00101110001000: color_data = 12'b010100000000;
		14'b00101110001001: color_data = 12'b010100000000;
		14'b00101110001010: color_data = 12'b101000000000;
		14'b00101110001011: color_data = 12'b101000000000;
		14'b00101110001100: color_data = 12'b010100000000;
		14'b00101110001101: color_data = 12'b010100000000;
		14'b00101110100000: color_data = 12'b010100000000;
		14'b00101110100001: color_data = 12'b010100000000;
		14'b00101110100111: color_data = 12'b010100000000;
		14'b00101110101000: color_data = 12'b010100000000;
		14'b00101110101001: color_data = 12'b101000000000;
		14'b00101110101010: color_data = 12'b101000000000;
		14'b00101110101011: color_data = 12'b101000000000;
		14'b00101110101100: color_data = 12'b010100000000;
		14'b00101110101111: color_data = 12'b010100000000;
		14'b00101111001010: color_data = 12'b010100000000;
		14'b00101111001011: color_data = 12'b010100000000;
		14'b00101111001100: color_data = 12'b101000000000;
		14'b00101111001101: color_data = 12'b101000000000;
		14'b00101111001110: color_data = 12'b101000000000;
		14'b00101111001111: color_data = 12'b101000000000;
		14'b00101111010000: color_data = 12'b010100000000;
		14'b00101111010001: color_data = 12'b010100000000;
		14'b00101111010010: color_data = 12'b101000000000;
		14'b00101111010011: color_data = 12'b101000000000;
		14'b00101111010100: color_data = 12'b101000000000;
		14'b00101111010101: color_data = 12'b101000000000;
		14'b00101111010110: color_data = 12'b010100000000;
		14'b00101111010111: color_data = 12'b010100000000;
		14'b00101111101000: color_data = 12'b010100000000;
		14'b00101111101001: color_data = 12'b010100000000;
		14'b00110000001000: color_data = 12'b010100000000;
		14'b00110000001001: color_data = 12'b010100000000;
		14'b00110000001010: color_data = 12'b101000000000;
		14'b00110000001011: color_data = 12'b010100000000;
		14'b00110000001100: color_data = 12'b010100000000;
		14'b00110000001101: color_data = 12'b010100000000;
		14'b00110000100000: color_data = 12'b010100000000;
		14'b00110000100001: color_data = 12'b010100000000;
		14'b00110000100111: color_data = 12'b010100000000;
		14'b00110000101000: color_data = 12'b101000000000;
		14'b00110000101001: color_data = 12'b101000000000;
		14'b00110000101010: color_data = 12'b101000000000;
		14'b00110000101011: color_data = 12'b101000000000;
		14'b00110000101100: color_data = 12'b010100000000;
		14'b00110001001001: color_data = 12'b010100000000;
		14'b00110001001010: color_data = 12'b010100000000;
		14'b00110001001011: color_data = 12'b101000000000;
		14'b00110001001100: color_data = 12'b101000000000;
		14'b00110001001101: color_data = 12'b101000000000;
		14'b00110001001110: color_data = 12'b101000000000;
		14'b00110001001111: color_data = 12'b010100000000;
		14'b00110001010000: color_data = 12'b010100000000;
		14'b00110001010001: color_data = 12'b010100000000;
		14'b00110001010010: color_data = 12'b101000000000;
		14'b00110001010011: color_data = 12'b101000000000;
		14'b00110001010100: color_data = 12'b101000000000;
		14'b00110001010101: color_data = 12'b101000000000;
		14'b00110001010110: color_data = 12'b010100000000;
		14'b00110001010111: color_data = 12'b010100000000;
		14'b00110001011000: color_data = 12'b010100000000;
		14'b00110001100111: color_data = 12'b010100000000;
		14'b00110001101000: color_data = 12'b010100000000;
		14'b00110001101001: color_data = 12'b010100000000;
		14'b00110010001000: color_data = 12'b010100000000;
		14'b00110010001001: color_data = 12'b010100000000;
		14'b00110010001010: color_data = 12'b010100000000;
		14'b00110010001011: color_data = 12'b010100000000;
		14'b00110010001101: color_data = 12'b010100000000;
		14'b00110010001110: color_data = 12'b010100000000;
		14'b00110010100101: color_data = 12'b010100000000;
		14'b00110010100110: color_data = 12'b010100000000;
		14'b00110010100111: color_data = 12'b101000000000;
		14'b00110010101000: color_data = 12'b101000000000;
		14'b00110010101001: color_data = 12'b101000000000;
		14'b00110010101010: color_data = 12'b101000000000;
		14'b00110010101011: color_data = 12'b010100000000;
		14'b00110010101100: color_data = 12'b010100000000;
		14'b00110011001000: color_data = 12'b010100000000;
		14'b00110011001001: color_data = 12'b010100000000;
		14'b00110011001010: color_data = 12'b101000000000;
		14'b00110011001011: color_data = 12'b101000000000;
		14'b00110011001100: color_data = 12'b101000000000;
		14'b00110011001101: color_data = 12'b101000000000;
		14'b00110011001110: color_data = 12'b101000000000;
		14'b00110011001111: color_data = 12'b010100000000;
		14'b00110011010000: color_data = 12'b010100000000;
		14'b00110011010001: color_data = 12'b101000000000;
		14'b00110011010010: color_data = 12'b101000000000;
		14'b00110011010011: color_data = 12'b101000000000;
		14'b00110011010100: color_data = 12'b101000000000;
		14'b00110011010101: color_data = 12'b101000000000;
		14'b00110011010110: color_data = 12'b010100000000;
		14'b00110011010111: color_data = 12'b010100000000;
		14'b00110011011000: color_data = 12'b010100000000;
		14'b00110011100111: color_data = 12'b010100000000;
		14'b00110011101000: color_data = 12'b010100000000;
		14'b00110011101001: color_data = 12'b010100000000;
		14'b00110100001000: color_data = 12'b010100000000;
		14'b00110100001001: color_data = 12'b010100000000;
		14'b00110100001010: color_data = 12'b010100000000;
		14'b00110100001011: color_data = 12'b010100000000;
		14'b00110100001110: color_data = 12'b010100000000;
		14'b00110100100100: color_data = 12'b010100000000;
		14'b00110100100101: color_data = 12'b010100000000;
		14'b00110100100110: color_data = 12'b101000000000;
		14'b00110100100111: color_data = 12'b101000000000;
		14'b00110100101000: color_data = 12'b101000000000;
		14'b00110100101001: color_data = 12'b101000000000;
		14'b00110100101010: color_data = 12'b101000000000;
		14'b00110100101011: color_data = 12'b010100000000;
		14'b00110101001000: color_data = 12'b010100000000;
		14'b00110101001001: color_data = 12'b101000000000;
		14'b00110101001010: color_data = 12'b101000000000;
		14'b00110101001011: color_data = 12'b010100000000;
		14'b00110101001100: color_data = 12'b010100000000;
		14'b00110101001101: color_data = 12'b101000000000;
		14'b00110101001110: color_data = 12'b101000000000;
		14'b00110101001111: color_data = 12'b010100000000;
		14'b00110101010000: color_data = 12'b010100000000;
		14'b00110101010001: color_data = 12'b101000000000;
		14'b00110101010010: color_data = 12'b101000000000;
		14'b00110101010011: color_data = 12'b101000000000;
		14'b00110101010100: color_data = 12'b101000000000;
		14'b00110101010101: color_data = 12'b101000000000;
		14'b00110101010110: color_data = 12'b010100000000;
		14'b00110101010111: color_data = 12'b010100000000;
		14'b00110101011000: color_data = 12'b010100000000;
		14'b00110101100111: color_data = 12'b010100000000;
		14'b00110101101000: color_data = 12'b010100000000;
		14'b00110101101001: color_data = 12'b010100000000;
		14'b00110110001000: color_data = 12'b010100000000;
		14'b00110110001001: color_data = 12'b010100000000;
		14'b00110110001010: color_data = 12'b010100000000;
		14'b00110110001011: color_data = 12'b010100000000;
		14'b00110110001111: color_data = 12'b010100000000;
		14'b00110110010000: color_data = 12'b010100000000;
		14'b00110110100001: color_data = 12'b010100000000;
		14'b00110110100010: color_data = 12'b010100000000;
		14'b00110110100011: color_data = 12'b010100000000;
		14'b00110110100100: color_data = 12'b010100000000;
		14'b00110110100101: color_data = 12'b101000000000;
		14'b00110110100110: color_data = 12'b101000000000;
		14'b00110110100111: color_data = 12'b101000000000;
		14'b00110110101000: color_data = 12'b101000000000;
		14'b00110110101001: color_data = 12'b101000000000;
		14'b00110110101010: color_data = 12'b010100000000;
		14'b00110111000111: color_data = 12'b010100000000;
		14'b00110111001000: color_data = 12'b010100000000;
		14'b00110111001001: color_data = 12'b010100000000;
		14'b00110111001010: color_data = 12'b010100000000;
		14'b00110111001011: color_data = 12'b010100000000;
		14'b00110111001100: color_data = 12'b101000000000;
		14'b00110111001101: color_data = 12'b101000000000;
		14'b00110111001110: color_data = 12'b101000000000;
		14'b00110111001111: color_data = 12'b010100000000;
		14'b00110111010000: color_data = 12'b010100000000;
		14'b00110111010001: color_data = 12'b101000000000;
		14'b00110111010010: color_data = 12'b101000000000;
		14'b00110111010011: color_data = 12'b101000000000;
		14'b00110111010100: color_data = 12'b101000000000;
		14'b00110111010101: color_data = 12'b101000000000;
		14'b00110111010110: color_data = 12'b010100000000;
		14'b00110111010111: color_data = 12'b010100000000;
		14'b00110111011000: color_data = 12'b010100000000;
		14'b00110111100111: color_data = 12'b010100000000;
		14'b00110111101000: color_data = 12'b010100000000;
		14'b00110111101001: color_data = 12'b010100000000;
		14'b00110111101010: color_data = 12'b010100000000;
		14'b00111000001001: color_data = 12'b010100000000;
		14'b00111000001010: color_data = 12'b010100000000;
		14'b00111000100001: color_data = 12'b010100000000;
		14'b00111000100010: color_data = 12'b010100000000;
		14'b00111000100011: color_data = 12'b101000000000;
		14'b00111000100100: color_data = 12'b101000000000;
		14'b00111000100101: color_data = 12'b101000000000;
		14'b00111000100110: color_data = 12'b101000000000;
		14'b00111000100111: color_data = 12'b101000000000;
		14'b00111000101000: color_data = 12'b101000000000;
		14'b00111000101001: color_data = 12'b010100000000;
		14'b00111000101010: color_data = 12'b010100000000;
		14'b00111001000110: color_data = 12'b010100000000;
		14'b00111001000111: color_data = 12'b010100000000;
		14'b00111001001000: color_data = 12'b010100000000;
		14'b00111001001001: color_data = 12'b010100000000;
		14'b00111001001010: color_data = 12'b101000000000;
		14'b00111001001011: color_data = 12'b101000000000;
		14'b00111001001100: color_data = 12'b101000000000;
		14'b00111001001101: color_data = 12'b101000000000;
		14'b00111001001110: color_data = 12'b101000000000;
		14'b00111001001111: color_data = 12'b010100000000;
		14'b00111001010000: color_data = 12'b010100000000;
		14'b00111001010001: color_data = 12'b010100000000;
		14'b00111001010010: color_data = 12'b101000000000;
		14'b00111001010011: color_data = 12'b101000000000;
		14'b00111001010100: color_data = 12'b101000000000;
		14'b00111001010101: color_data = 12'b101000000000;
		14'b00111001010110: color_data = 12'b010100000000;
		14'b00111001010111: color_data = 12'b010100000000;
		14'b00111001011000: color_data = 12'b010100000000;
		14'b00111001011001: color_data = 12'b010100000000;
		14'b00111001100111: color_data = 12'b010100000000;
		14'b00111001101000: color_data = 12'b010100000000;
		14'b00111001101001: color_data = 12'b010100000000;
		14'b00111001101010: color_data = 12'b010100000000;
		14'b00111010001001: color_data = 12'b010100000000;
		14'b00111010001010: color_data = 12'b010100000000;
		14'b00111010100000: color_data = 12'b010100000000;
		14'b00111010100001: color_data = 12'b010100000000;
		14'b00111010100010: color_data = 12'b101000000000;
		14'b00111010100011: color_data = 12'b101000000000;
		14'b00111010100100: color_data = 12'b101000000000;
		14'b00111010100101: color_data = 12'b101000000000;
		14'b00111010100110: color_data = 12'b101000000000;
		14'b00111010100111: color_data = 12'b010100000000;
		14'b00111010101000: color_data = 12'b010100000000;
		14'b00111011000101: color_data = 12'b010100000000;
		14'b00111011000110: color_data = 12'b010100000000;
		14'b00111011000111: color_data = 12'b101000000000;
		14'b00111011001000: color_data = 12'b101000000000;
		14'b00111011001001: color_data = 12'b101000000000;
		14'b00111011001010: color_data = 12'b101000000000;
		14'b00111011001011: color_data = 12'b101000000000;
		14'b00111011001100: color_data = 12'b101000000000;
		14'b00111011001101: color_data = 12'b101000000000;
		14'b00111011001110: color_data = 12'b101000000000;
		14'b00111011001111: color_data = 12'b101000000000;
		14'b00111011010000: color_data = 12'b010100000000;
		14'b00111011010001: color_data = 12'b010100000000;
		14'b00111011010010: color_data = 12'b010100000000;
		14'b00111011010011: color_data = 12'b101000000000;
		14'b00111011010100: color_data = 12'b101000000000;
		14'b00111011010101: color_data = 12'b101000000000;
		14'b00111011010110: color_data = 12'b101000000000;
		14'b00111011010111: color_data = 12'b010100000000;
		14'b00111011011000: color_data = 12'b010100000000;
		14'b00111011011001: color_data = 12'b010100000000;
		14'b00111011101001: color_data = 12'b010100000000;
		14'b00111011101010: color_data = 12'b010100000000;
		14'b00111100001010: color_data = 12'b010100000000;
		14'b00111100011111: color_data = 12'b010100000000;
		14'b00111100100000: color_data = 12'b010100000000;
		14'b00111100100001: color_data = 12'b101000000000;
		14'b00111100100010: color_data = 12'b101000000000;
		14'b00111100100011: color_data = 12'b101000000000;
		14'b00111100100100: color_data = 12'b101000000000;
		14'b00111100100101: color_data = 12'b101000000000;
		14'b00111100100110: color_data = 12'b010100000000;
		14'b00111100100111: color_data = 12'b010100000000;
		14'b00111101000011: color_data = 12'b010100000000;
		14'b00111101000100: color_data = 12'b010100000000;
		14'b00111101000101: color_data = 12'b101000000000;
		14'b00111101000110: color_data = 12'b101000000000;
		14'b00111101000111: color_data = 12'b101000000000;
		14'b00111101001000: color_data = 12'b101000000000;
		14'b00111101001001: color_data = 12'b101000000000;
		14'b00111101001010: color_data = 12'b101000000000;
		14'b00111101001011: color_data = 12'b101000000000;
		14'b00111101001100: color_data = 12'b101000000000;
		14'b00111101001101: color_data = 12'b101000000000;
		14'b00111101001110: color_data = 12'b101000000000;
		14'b00111101001111: color_data = 12'b101000000000;
		14'b00111101010000: color_data = 12'b010100000000;
		14'b00111101010001: color_data = 12'b010100000000;
		14'b00111101010010: color_data = 12'b010100000000;
		14'b00111101010011: color_data = 12'b010100000000;
		14'b00111101010100: color_data = 12'b101000000000;
		14'b00111101010101: color_data = 12'b101000000000;
		14'b00111101010110: color_data = 12'b101000000000;
		14'b00111101010111: color_data = 12'b010100000000;
		14'b00111101011000: color_data = 12'b010100000000;
		14'b00111101011001: color_data = 12'b010100000000;
		14'b00111101101001: color_data = 12'b010100000000;
		14'b00111101101010: color_data = 12'b010100000000;
		14'b00111110001011: color_data = 12'b010100000000;
		14'b00111110011110: color_data = 12'b010100000000;
		14'b00111110011111: color_data = 12'b010100000000;
		14'b00111110100000: color_data = 12'b010100000000;
		14'b00111110100001: color_data = 12'b010100000000;
		14'b00111110100010: color_data = 12'b010100000000;
		14'b00111110100011: color_data = 12'b010100000000;
		14'b00111110100100: color_data = 12'b010100000000;
		14'b00111110100101: color_data = 12'b010100000000;
		14'b00111110100110: color_data = 12'b010100000000;
		14'b00111111000010: color_data = 12'b010100000000;
		14'b00111111000011: color_data = 12'b101000000000;
		14'b00111111000100: color_data = 12'b101000000000;
		14'b00111111000101: color_data = 12'b101000000000;
		14'b00111111000110: color_data = 12'b101000000000;
		14'b00111111000111: color_data = 12'b101000000000;
		14'b00111111001000: color_data = 12'b101000000000;
		14'b00111111001001: color_data = 12'b101000000000;
		14'b00111111001010: color_data = 12'b101000000000;
		14'b00111111001011: color_data = 12'b101000000000;
		14'b00111111001100: color_data = 12'b101000000000;
		14'b00111111001101: color_data = 12'b101000000000;
		14'b00111111001110: color_data = 12'b101000000000;
		14'b00111111001111: color_data = 12'b101000000000;
		14'b00111111010000: color_data = 12'b101000000000;
		14'b00111111010001: color_data = 12'b010100000000;
		14'b00111111010010: color_data = 12'b010100000000;
		14'b00111111010011: color_data = 12'b010100000000;
		14'b00111111010100: color_data = 12'b010100000000;
		14'b00111111010101: color_data = 12'b101000000000;
		14'b00111111010110: color_data = 12'b101000000000;
		14'b00111111010111: color_data = 12'b101000000000;
		14'b00111111011000: color_data = 12'b010100000000;
		14'b00111111011001: color_data = 12'b010100000000;
		14'b00111111101010: color_data = 12'b010100000000;
		14'b01000000011101: color_data = 12'b010100000000;
		14'b01000000011110: color_data = 12'b010100000000;
		14'b01000000011111: color_data = 12'b010100000000;
		14'b01000000100000: color_data = 12'b010100000000;
		14'b01000000100001: color_data = 12'b010100000000;
		14'b01000000100010: color_data = 12'b010100000000;
		14'b01000000100011: color_data = 12'b010100000000;
		14'b01000000100100: color_data = 12'b010100000000;
		14'b01000001000001: color_data = 12'b010100000000;
		14'b01000001000010: color_data = 12'b101000000000;
		14'b01000001000011: color_data = 12'b101000000000;
		14'b01000001000100: color_data = 12'b101000000000;
		14'b01000001000101: color_data = 12'b101000000000;
		14'b01000001000110: color_data = 12'b101000000000;
		14'b01000001000111: color_data = 12'b101000000000;
		14'b01000001001000: color_data = 12'b101000000000;
		14'b01000001001001: color_data = 12'b101000000000;
		14'b01000001001010: color_data = 12'b101000000000;
		14'b01000001001011: color_data = 12'b101000000000;
		14'b01000001001100: color_data = 12'b101000000000;
		14'b01000001001101: color_data = 12'b101000000000;
		14'b01000001001110: color_data = 12'b101000000000;
		14'b01000001001111: color_data = 12'b101000000000;
		14'b01000001010000: color_data = 12'b101000000000;
		14'b01000001010001: color_data = 12'b101000000000;
		14'b01000001010010: color_data = 12'b010100000000;
		14'b01000001010011: color_data = 12'b010100000000;
		14'b01000001010100: color_data = 12'b010100000000;
		14'b01000001010101: color_data = 12'b010100000000;
		14'b01000001010110: color_data = 12'b010100000000;
		14'b01000001010111: color_data = 12'b010100000000;
		14'b01000001011000: color_data = 12'b010100000000;
		14'b01000001011001: color_data = 12'b010100000000;
		14'b01000010011101: color_data = 12'b010100000000;
		14'b01000010011110: color_data = 12'b010100000000;
		14'b01000010011111: color_data = 12'b010100000000;
		14'b01000010100000: color_data = 12'b010100000000;
		14'b01000010100001: color_data = 12'b010100000000;
		14'b01000010111111: color_data = 12'b010100000000;
		14'b01000011000000: color_data = 12'b010100000000;
		14'b01000011000001: color_data = 12'b101000000000;
		14'b01000011000010: color_data = 12'b101000000000;
		14'b01000011000011: color_data = 12'b101000000000;
		14'b01000011000100: color_data = 12'b101000000000;
		14'b01000011000101: color_data = 12'b101000000000;
		14'b01000011000110: color_data = 12'b101000000000;
		14'b01000011000111: color_data = 12'b101000000000;
		14'b01000011001000: color_data = 12'b101000000000;
		14'b01000011001001: color_data = 12'b101000000000;
		14'b01000011001010: color_data = 12'b101000000000;
		14'b01000011001011: color_data = 12'b101000000000;
		14'b01000011001100: color_data = 12'b101000000000;
		14'b01000011001101: color_data = 12'b101000000000;
		14'b01000011001110: color_data = 12'b101000000000;
		14'b01000011001111: color_data = 12'b101000000000;
		14'b01000011010000: color_data = 12'b101000000000;
		14'b01000011010001: color_data = 12'b101000000000;
		14'b01000011010010: color_data = 12'b010100000000;
		14'b01000011010011: color_data = 12'b010100000000;
		14'b01000011010110: color_data = 12'b010100000000;
		14'b01000011010111: color_data = 12'b010100000000;
		14'b01000011011000: color_data = 12'b010100000000;
		14'b01000011011001: color_data = 12'b010100000000;
		14'b01000011011010: color_data = 12'b010100000000;
		14'b01000100011101: color_data = 12'b010100000000;
		14'b01000100011110: color_data = 12'b010100000000;
		14'b01000100011111: color_data = 12'b010100000000;
		14'b01000100111101: color_data = 12'b010100000000;
		14'b01000100111110: color_data = 12'b010100000000;
		14'b01000100111111: color_data = 12'b101000000000;
		14'b01000101000000: color_data = 12'b101000000000;
		14'b01000101000001: color_data = 12'b101000000000;
		14'b01000101000010: color_data = 12'b101000000000;
		14'b01000101000011: color_data = 12'b101000000000;
		14'b01000101000100: color_data = 12'b101000000000;
		14'b01000101000101: color_data = 12'b101000000000;
		14'b01000101000110: color_data = 12'b101000000000;
		14'b01000101000111: color_data = 12'b101000000000;
		14'b01000101001000: color_data = 12'b101000000000;
		14'b01000101001001: color_data = 12'b101000000000;
		14'b01000101001010: color_data = 12'b101000000000;
		14'b01000101001011: color_data = 12'b101000000000;
		14'b01000101001100: color_data = 12'b101000000000;
		14'b01000101001101: color_data = 12'b101000000000;
		14'b01000101001110: color_data = 12'b101000000000;
		14'b01000101001111: color_data = 12'b101000000000;
		14'b01000101010000: color_data = 12'b101000000000;
		14'b01000101010001: color_data = 12'b101000000000;
		14'b01000101010010: color_data = 12'b101000000000;
		14'b01000101010011: color_data = 12'b010100000000;
		14'b01000101011000: color_data = 12'b010100000000;
		14'b01000101011001: color_data = 12'b010100000000;
		14'b01000101011010: color_data = 12'b010100000000;
		14'b01000110011101: color_data = 12'b010100000000;
		14'b01000110111011: color_data = 12'b010100000000;
		14'b01000110111100: color_data = 12'b010100000000;
		14'b01000110111101: color_data = 12'b101000000000;
		14'b01000110111110: color_data = 12'b101000000000;
		14'b01000110111111: color_data = 12'b101000000000;
		14'b01000111000000: color_data = 12'b101000000000;
		14'b01000111000001: color_data = 12'b101000000000;
		14'b01000111000010: color_data = 12'b101000000000;
		14'b01000111000011: color_data = 12'b101000000000;
		14'b01000111000100: color_data = 12'b101000000000;
		14'b01000111000101: color_data = 12'b101000000000;
		14'b01000111000110: color_data = 12'b101000000000;
		14'b01000111000111: color_data = 12'b101000000000;
		14'b01000111001000: color_data = 12'b101000000000;
		14'b01000111001001: color_data = 12'b101000000000;
		14'b01000111001010: color_data = 12'b101000000000;
		14'b01000111001011: color_data = 12'b101000000000;
		14'b01000111001100: color_data = 12'b101000000000;
		14'b01000111001101: color_data = 12'b101000000000;
		14'b01000111001110: color_data = 12'b101000000000;
		14'b01000111001111: color_data = 12'b101000000000;
		14'b01000111010000: color_data = 12'b101000000000;
		14'b01000111010001: color_data = 12'b101000000000;
		14'b01000111010010: color_data = 12'b101000000000;
		14'b01000111010011: color_data = 12'b101000000000;
		14'b01000111010100: color_data = 12'b010100000000;
		14'b01000111011001: color_data = 12'b010100000000;
		14'b01000111011010: color_data = 12'b010100000000;
		14'b01000111011011: color_data = 12'b010100000000;
		14'b01001000011110: color_data = 12'b010100000000;
		14'b01001000111001: color_data = 12'b010100000000;
		14'b01001000111010: color_data = 12'b010100000000;
		14'b01001000111011: color_data = 12'b101000000000;
		14'b01001000111100: color_data = 12'b101000000000;
		14'b01001000111101: color_data = 12'b101000000000;
		14'b01001000111110: color_data = 12'b101000000000;
		14'b01001000111111: color_data = 12'b101000000000;
		14'b01001001000000: color_data = 12'b101000000000;
		14'b01001001000001: color_data = 12'b101000000000;
		14'b01001001000010: color_data = 12'b101000000000;
		14'b01001001000011: color_data = 12'b101000000000;
		14'b01001001000100: color_data = 12'b101000000000;
		14'b01001001000101: color_data = 12'b101000000000;
		14'b01001001000110: color_data = 12'b101000000000;
		14'b01001001000111: color_data = 12'b101000000000;
		14'b01001001001000: color_data = 12'b101000000000;
		14'b01001001001001: color_data = 12'b101000000000;
		14'b01001001001010: color_data = 12'b101000000000;
		14'b01001001001011: color_data = 12'b101000000000;
		14'b01001001001100: color_data = 12'b101000000000;
		14'b01001001001101: color_data = 12'b101000000000;
		14'b01001001001110: color_data = 12'b101000000000;
		14'b01001001001111: color_data = 12'b101000000000;
		14'b01001001010000: color_data = 12'b101000000000;
		14'b01001001010001: color_data = 12'b101000000000;
		14'b01001001010010: color_data = 12'b101000000000;
		14'b01001001010011: color_data = 12'b101000000000;
		14'b01001001010100: color_data = 12'b010100000000;
		14'b01001001010101: color_data = 12'b010100000000;
		14'b01001001011011: color_data = 12'b010100000000;
		14'b01001010110111: color_data = 12'b010100000000;
		14'b01001010111000: color_data = 12'b010100000000;
		14'b01001010111001: color_data = 12'b101000000000;
		14'b01001010111010: color_data = 12'b101000000000;
		14'b01001010111011: color_data = 12'b101000000000;
		14'b01001010111100: color_data = 12'b101000000000;
		14'b01001010111101: color_data = 12'b101000000000;
		14'b01001010111110: color_data = 12'b101000000000;
		14'b01001010111111: color_data = 12'b101000000000;
		14'b01001011000000: color_data = 12'b101000000000;
		14'b01001011000001: color_data = 12'b101000000000;
		14'b01001011000010: color_data = 12'b101000000000;
		14'b01001011000011: color_data = 12'b101000000000;
		14'b01001011000100: color_data = 12'b101000000000;
		14'b01001011000101: color_data = 12'b101000000000;
		14'b01001011000110: color_data = 12'b101000000000;
		14'b01001011000111: color_data = 12'b101000000000;
		14'b01001011001000: color_data = 12'b101000000000;
		14'b01001011001001: color_data = 12'b101000000000;
		14'b01001011001010: color_data = 12'b101000000000;
		14'b01001011001011: color_data = 12'b101000000000;
		14'b01001011001100: color_data = 12'b101000000000;
		14'b01001011001101: color_data = 12'b101000000000;
		14'b01001011001110: color_data = 12'b010100000000;
		14'b01001011001111: color_data = 12'b010100000000;
		14'b01001011010000: color_data = 12'b010100000000;
		14'b01001011010001: color_data = 12'b101000000000;
		14'b01001011010010: color_data = 12'b101000000000;
		14'b01001011010011: color_data = 12'b101000000000;
		14'b01001011010100: color_data = 12'b101000000000;
		14'b01001011010101: color_data = 12'b101000000000;
		14'b01001011010110: color_data = 12'b010100000000;
		14'b01001100101100: color_data = 12'b010100000000;
		14'b01001100110100: color_data = 12'b010100000000;
		14'b01001100110101: color_data = 12'b010100000000;
		14'b01001100110110: color_data = 12'b010100000000;
		14'b01001100110111: color_data = 12'b010100000000;
		14'b01001100111000: color_data = 12'b101000000000;
		14'b01001100111001: color_data = 12'b101000000000;
		14'b01001100111010: color_data = 12'b101000000000;
		14'b01001100111011: color_data = 12'b101000000000;
		14'b01001100111100: color_data = 12'b101000000000;
		14'b01001100111101: color_data = 12'b101000000000;
		14'b01001100111110: color_data = 12'b101000000000;
		14'b01001100111111: color_data = 12'b101000000000;
		14'b01001101000000: color_data = 12'b101000000000;
		14'b01001101000001: color_data = 12'b101000000000;
		14'b01001101000010: color_data = 12'b101000000000;
		14'b01001101000011: color_data = 12'b101000000000;
		14'b01001101000100: color_data = 12'b101000000000;
		14'b01001101000101: color_data = 12'b101000000000;
		14'b01001101000110: color_data = 12'b101000000000;
		14'b01001101000111: color_data = 12'b101000000000;
		14'b01001101001000: color_data = 12'b101000000000;
		14'b01001101001001: color_data = 12'b101000000000;
		14'b01001101001010: color_data = 12'b101000000000;
		14'b01001101001011: color_data = 12'b101000000000;
		14'b01001101001100: color_data = 12'b101000000000;
		14'b01001101001101: color_data = 12'b101000000000;
		14'b01001101001110: color_data = 12'b101000000000;
		14'b01001101001111: color_data = 12'b101000000000;
		14'b01001101010000: color_data = 12'b010100000000;
		14'b01001101010001: color_data = 12'b010100000000;
		14'b01001101010010: color_data = 12'b010100000000;
		14'b01001101010011: color_data = 12'b101000000000;
		14'b01001101010100: color_data = 12'b101000000000;
		14'b01001101010101: color_data = 12'b101000000000;
		14'b01001101010110: color_data = 12'b101000000000;
		14'b01001101010111: color_data = 12'b010100000000;
		14'b01001110000000: color_data = 12'b010100000000;
		14'b01001110000001: color_data = 12'b010100000000;
		14'b01001110000010: color_data = 12'b010100000000;
		14'b01001110000011: color_data = 12'b010100000000;
		14'b01001110000100: color_data = 12'b010100000000;
		14'b01001110010010: color_data = 12'b010100000000;
		14'b01001110010011: color_data = 12'b101000000000;
		14'b01001110010100: color_data = 12'b010100000000;
		14'b01001110010101: color_data = 12'b010100000000;
		14'b01001110101010: color_data = 12'b010100000000;
		14'b01001110101011: color_data = 12'b010100000000;
		14'b01001110101100: color_data = 12'b010100000000;
		14'b01001110101101: color_data = 12'b010100000000;
		14'b01001110101110: color_data = 12'b010100000000;
		14'b01001110101111: color_data = 12'b010100000000;
		14'b01001110110000: color_data = 12'b010100000000;
		14'b01001110110001: color_data = 12'b010100000000;
		14'b01001110110010: color_data = 12'b010100000000;
		14'b01001110110011: color_data = 12'b010100000000;
		14'b01001110110100: color_data = 12'b010100000000;
		14'b01001110110101: color_data = 12'b010100000000;
		14'b01001110110110: color_data = 12'b101000000000;
		14'b01001110110111: color_data = 12'b101000000000;
		14'b01001110111000: color_data = 12'b101000000000;
		14'b01001110111001: color_data = 12'b101000000000;
		14'b01001110111010: color_data = 12'b101000000000;
		14'b01001110111011: color_data = 12'b101000000000;
		14'b01001110111100: color_data = 12'b101000000000;
		14'b01001110111101: color_data = 12'b101000000000;
		14'b01001110111110: color_data = 12'b101000000000;
		14'b01001110111111: color_data = 12'b101000000000;
		14'b01001111000000: color_data = 12'b101000000000;
		14'b01001111000001: color_data = 12'b101000000000;
		14'b01001111000010: color_data = 12'b101000000000;
		14'b01001111000011: color_data = 12'b101000000000;
		14'b01001111000100: color_data = 12'b101000000000;
		14'b01001111000101: color_data = 12'b101000000000;
		14'b01001111000110: color_data = 12'b101000000000;
		14'b01001111000111: color_data = 12'b101000000000;
		14'b01001111001000: color_data = 12'b101000000000;
		14'b01001111001001: color_data = 12'b101000000000;
		14'b01001111001010: color_data = 12'b101000000000;
		14'b01001111001011: color_data = 12'b101000000000;
		14'b01001111001100: color_data = 12'b101000000000;
		14'b01001111001101: color_data = 12'b101000000000;
		14'b01001111001110: color_data = 12'b101000000000;
		14'b01001111001111: color_data = 12'b101000000000;
		14'b01001111010000: color_data = 12'b101000000000;
		14'b01001111010001: color_data = 12'b101000000000;
		14'b01001111010010: color_data = 12'b101000000000;
		14'b01001111010011: color_data = 12'b010100000000;
		14'b01001111010100: color_data = 12'b101000000000;
		14'b01001111010101: color_data = 12'b101000000000;
		14'b01001111010110: color_data = 12'b101000000000;
		14'b01001111010111: color_data = 12'b101000000000;
		14'b01001111011000: color_data = 12'b010100000000;
		14'b01010000000010: color_data = 12'b010100000000;
		14'b01010000000011: color_data = 12'b010100000000;
		14'b01010000000100: color_data = 12'b101000000000;
		14'b01010000000101: color_data = 12'b010100000000;
		14'b01010000000110: color_data = 12'b010100000000;
		14'b01010000000111: color_data = 12'b010100000000;
		14'b01010000001101: color_data = 12'b010100000000;
		14'b01010000010011: color_data = 12'b010100000000;
		14'b01010000010100: color_data = 12'b101000000000;
		14'b01010000010101: color_data = 12'b101000000000;
		14'b01010000010110: color_data = 12'b101000000000;
		14'b01010000010111: color_data = 12'b101000000000;
		14'b01010000011000: color_data = 12'b010100000000;
		14'b01010000011001: color_data = 12'b010100000000;
		14'b01010000011010: color_data = 12'b010100000000;
		14'b01010000011011: color_data = 12'b010100000000;
		14'b01010000011100: color_data = 12'b010100000000;
		14'b01010000011101: color_data = 12'b010100000000;
		14'b01010000011110: color_data = 12'b010100000000;
		14'b01010000011111: color_data = 12'b010100000000;
		14'b01010000100000: color_data = 12'b010100000000;
		14'b01010000100001: color_data = 12'b010100000000;
		14'b01010000100101: color_data = 12'b010100000000;
		14'b01010000100110: color_data = 12'b010100000000;
		14'b01010000100111: color_data = 12'b010100000000;
		14'b01010000101000: color_data = 12'b010100000000;
		14'b01010000101001: color_data = 12'b010100000000;
		14'b01010000101010: color_data = 12'b010100000000;
		14'b01010000101011: color_data = 12'b010100000000;
		14'b01010000101100: color_data = 12'b010100000000;
		14'b01010000101101: color_data = 12'b010100000000;
		14'b01010000101110: color_data = 12'b010100000000;
		14'b01010000101111: color_data = 12'b010100000000;
		14'b01010000110000: color_data = 12'b010100000000;
		14'b01010000110001: color_data = 12'b101000000000;
		14'b01010000110010: color_data = 12'b101000000000;
		14'b01010000110011: color_data = 12'b101000000000;
		14'b01010000110100: color_data = 12'b101000000000;
		14'b01010000110101: color_data = 12'b101000000000;
		14'b01010000110110: color_data = 12'b101000000000;
		14'b01010000110111: color_data = 12'b101000000000;
		14'b01010000111000: color_data = 12'b101000000000;
		14'b01010000111001: color_data = 12'b101000000000;
		14'b01010000111010: color_data = 12'b101000000000;
		14'b01010000111011: color_data = 12'b101000000000;
		14'b01010000111100: color_data = 12'b101000000000;
		14'b01010000111101: color_data = 12'b101000000000;
		14'b01010000111110: color_data = 12'b010100000000;
		14'b01010000111111: color_data = 12'b010100000000;
		14'b01010001000000: color_data = 12'b010100000000;
		14'b01010001000001: color_data = 12'b010100000000;
		14'b01010001000010: color_data = 12'b010100000000;
		14'b01010001000011: color_data = 12'b010100000000;
		14'b01010001000100: color_data = 12'b010100000000;
		14'b01010001000101: color_data = 12'b010100000000;
		14'b01010001000110: color_data = 12'b010100000000;
		14'b01010001000111: color_data = 12'b010100000000;
		14'b01010001001000: color_data = 12'b101000000000;
		14'b01010001001001: color_data = 12'b101000000000;
		14'b01010001001010: color_data = 12'b101000000000;
		14'b01010001001011: color_data = 12'b101000000000;
		14'b01010001001100: color_data = 12'b010100000000;
		14'b01010001001101: color_data = 12'b010100000000;
		14'b01010001001110: color_data = 12'b010100000000;
		14'b01010001001111: color_data = 12'b101000000000;
		14'b01010001010000: color_data = 12'b101000000000;
		14'b01010001010001: color_data = 12'b101000000000;
		14'b01010001010010: color_data = 12'b101000000000;
		14'b01010001010011: color_data = 12'b101000000000;
		14'b01010001010100: color_data = 12'b010100000000;
		14'b01010001010101: color_data = 12'b101000000000;
		14'b01010001010110: color_data = 12'b101000000000;
		14'b01010001010111: color_data = 12'b101000000000;
		14'b01010001011000: color_data = 12'b101000000000;
		14'b01010001011001: color_data = 12'b101000000000;
		14'b01010001011010: color_data = 12'b010100000000;
		14'b01010010000100: color_data = 12'b010100000000;
		14'b01010010000101: color_data = 12'b010100000000;
		14'b01010010000110: color_data = 12'b101000000000;
		14'b01010010000111: color_data = 12'b101000000000;
		14'b01010010001000: color_data = 12'b101000000000;
		14'b01010010001001: color_data = 12'b010100000000;
		14'b01010010001010: color_data = 12'b010100000000;
		14'b01010010001011: color_data = 12'b010100000000;
		14'b01010010001110: color_data = 12'b010100000000;
		14'b01010010001111: color_data = 12'b010100000000;
		14'b01010010010000: color_data = 12'b010100000000;
		14'b01010010010100: color_data = 12'b010100000000;
		14'b01010010010101: color_data = 12'b101000000000;
		14'b01010010010110: color_data = 12'b101000000000;
		14'b01010010010111: color_data = 12'b101000000000;
		14'b01010010011000: color_data = 12'b101000000000;
		14'b01010010011001: color_data = 12'b101000000000;
		14'b01010010011010: color_data = 12'b101000000000;
		14'b01010010011011: color_data = 12'b101000000000;
		14'b01010010011100: color_data = 12'b101000000000;
		14'b01010010011101: color_data = 12'b101000000000;
		14'b01010010011110: color_data = 12'b101000000000;
		14'b01010010011111: color_data = 12'b101000000000;
		14'b01010010100000: color_data = 12'b101000000000;
		14'b01010010100001: color_data = 12'b101000000000;
		14'b01010010100010: color_data = 12'b010100000000;
		14'b01010010100011: color_data = 12'b010100000000;
		14'b01010010100100: color_data = 12'b010100000000;
		14'b01010010100101: color_data = 12'b010100000000;
		14'b01010010100110: color_data = 12'b010100000000;
		14'b01010010100111: color_data = 12'b010100000000;
		14'b01010010101000: color_data = 12'b010100000000;
		14'b01010010101001: color_data = 12'b010100000000;
		14'b01010010101010: color_data = 12'b010100000000;
		14'b01010010101011: color_data = 12'b010100000000;
		14'b01010010101100: color_data = 12'b010100000000;
		14'b01010010101101: color_data = 12'b010100000000;
		14'b01010010101110: color_data = 12'b101000000000;
		14'b01010010101111: color_data = 12'b101000000000;
		14'b01010010110000: color_data = 12'b101000000000;
		14'b01010010110001: color_data = 12'b101000000000;
		14'b01010010110010: color_data = 12'b101000000000;
		14'b01010010110011: color_data = 12'b101000000000;
		14'b01010010110100: color_data = 12'b101000000000;
		14'b01010010110101: color_data = 12'b101000000000;
		14'b01010010110110: color_data = 12'b101000000000;
		14'b01010010110111: color_data = 12'b101000000000;
		14'b01010010111000: color_data = 12'b101000000000;
		14'b01010010111001: color_data = 12'b101000000000;
		14'b01010010111010: color_data = 12'b101000000000;
		14'b01010010111011: color_data = 12'b101000000000;
		14'b01010010111100: color_data = 12'b101000000000;
		14'b01010010111101: color_data = 12'b010100000000;
		14'b01010010111110: color_data = 12'b010100000000;
		14'b01010010111111: color_data = 12'b010100000000;
		14'b01010011000000: color_data = 12'b010100000000;
		14'b01010011000001: color_data = 12'b010100000000;
		14'b01010011000010: color_data = 12'b010100000000;
		14'b01010011000011: color_data = 12'b010100000000;
		14'b01010011000100: color_data = 12'b010100000000;
		14'b01010011000101: color_data = 12'b010100000000;
		14'b01010011000110: color_data = 12'b010100000000;
		14'b01010011000111: color_data = 12'b010100000000;
		14'b01010011001000: color_data = 12'b010100000000;
		14'b01010011001001: color_data = 12'b010100000000;
		14'b01010011001010: color_data = 12'b010100000000;
		14'b01010011001011: color_data = 12'b010100000000;
		14'b01010011001100: color_data = 12'b010100000000;
		14'b01010011001101: color_data = 12'b010100000000;
		14'b01010011001110: color_data = 12'b010100000000;
		14'b01010011001111: color_data = 12'b010100000000;
		14'b01010011010000: color_data = 12'b010100000000;
		14'b01010011010001: color_data = 12'b010100000000;
		14'b01010011010010: color_data = 12'b101000000000;
		14'b01010011010011: color_data = 12'b101000000000;
		14'b01010011010100: color_data = 12'b101000000000;
		14'b01010011010101: color_data = 12'b101000000000;
		14'b01010011010110: color_data = 12'b101000000000;
		14'b01010011010111: color_data = 12'b101000000000;
		14'b01010011011000: color_data = 12'b101000000000;
		14'b01010011011001: color_data = 12'b101000000000;
		14'b01010011011010: color_data = 12'b101000000000;
		14'b01010011011011: color_data = 12'b010100000000;
		14'b01010100000110: color_data = 12'b010100000000;
		14'b01010100000111: color_data = 12'b010100000000;
		14'b01010100001000: color_data = 12'b010100000000;
		14'b01010100001001: color_data = 12'b010100000000;
		14'b01010100001010: color_data = 12'b101000000000;
		14'b01010100001011: color_data = 12'b101000000000;
		14'b01010100001100: color_data = 12'b101000000000;
		14'b01010100001101: color_data = 12'b010100000000;
		14'b01010100001110: color_data = 12'b010100000000;
		14'b01010100001111: color_data = 12'b101000000000;
		14'b01010100010000: color_data = 12'b101000000000;
		14'b01010100010001: color_data = 12'b010100000000;
		14'b01010100010101: color_data = 12'b010100000000;
		14'b01010100010110: color_data = 12'b010100000000;
		14'b01010100010111: color_data = 12'b101000000000;
		14'b01010100011000: color_data = 12'b101000000000;
		14'b01010100011001: color_data = 12'b101000000000;
		14'b01010100011010: color_data = 12'b101000000000;
		14'b01010100011011: color_data = 12'b010100000000;
		14'b01010100011100: color_data = 12'b010100000000;
		14'b01010100011101: color_data = 12'b010100000000;
		14'b01010100011110: color_data = 12'b010100000000;
		14'b01010100011111: color_data = 12'b010100000000;
		14'b01010100100000: color_data = 12'b101000000000;
		14'b01010100100001: color_data = 12'b101000000000;
		14'b01010100100010: color_data = 12'b101000000000;
		14'b01010100100011: color_data = 12'b101000000000;
		14'b01010100100100: color_data = 12'b101000000000;
		14'b01010100100101: color_data = 12'b101000000000;
		14'b01010100100110: color_data = 12'b101000000000;
		14'b01010100100111: color_data = 12'b101000000000;
		14'b01010100101000: color_data = 12'b010100000000;
		14'b01010100101001: color_data = 12'b010100000000;
		14'b01010100101010: color_data = 12'b010100000000;
		14'b01010100101011: color_data = 12'b010100000000;
		14'b01010100101100: color_data = 12'b010100000000;
		14'b01010100101101: color_data = 12'b010100000000;
		14'b01010100101110: color_data = 12'b101000000000;
		14'b01010100101111: color_data = 12'b101000000000;
		14'b01010100110000: color_data = 12'b101000000000;
		14'b01010100110001: color_data = 12'b101000000000;
		14'b01010100110010: color_data = 12'b101000000000;
		14'b01010100110011: color_data = 12'b101000000000;
		14'b01010100110100: color_data = 12'b101000000000;
		14'b01010100110101: color_data = 12'b101000000000;
		14'b01010100110110: color_data = 12'b101000000000;
		14'b01010100110111: color_data = 12'b101000000000;
		14'b01010100111000: color_data = 12'b101000000000;
		14'b01010100111001: color_data = 12'b010100000000;
		14'b01010100111010: color_data = 12'b010100000000;
		14'b01010100111011: color_data = 12'b101000000000;
		14'b01010100111100: color_data = 12'b010100000000;
		14'b01010100111101: color_data = 12'b010100000000;
		14'b01010100111110: color_data = 12'b010100000000;
		14'b01010100111111: color_data = 12'b010100000000;
		14'b01010101000000: color_data = 12'b010100000000;
		14'b01010101001101: color_data = 12'b010100000000;
		14'b01010101001110: color_data = 12'b010100000000;
		14'b01010101001111: color_data = 12'b010100000000;
		14'b01010101010000: color_data = 12'b010100000000;
		14'b01010101010001: color_data = 12'b010100000000;
		14'b01010101010010: color_data = 12'b010100000000;
		14'b01010101010011: color_data = 12'b010100000000;
		14'b01010101010100: color_data = 12'b101000000000;
		14'b01010101010101: color_data = 12'b101000000000;
		14'b01010101010110: color_data = 12'b010100000000;
		14'b01010101010111: color_data = 12'b010100000000;
		14'b01010101011000: color_data = 12'b101000000000;
		14'b01010101011001: color_data = 12'b101000000000;
		14'b01010101011010: color_data = 12'b101000000000;
		14'b01010101011011: color_data = 12'b101000000000;
		14'b01010101011100: color_data = 12'b010100000000;
		14'b01010110001100: color_data = 12'b010100000000;
		14'b01010110001101: color_data = 12'b010100000000;
		14'b01010110001110: color_data = 12'b010100000000;
		14'b01010110001111: color_data = 12'b010100000000;
		14'b01010110010000: color_data = 12'b101000000000;
		14'b01010110010001: color_data = 12'b101000000000;
		14'b01010110010010: color_data = 12'b010100000000;
		14'b01010110010111: color_data = 12'b010100000000;
		14'b01010110011000: color_data = 12'b010100000000;
		14'b01010110011001: color_data = 12'b101000000000;
		14'b01010110011010: color_data = 12'b101000000000;
		14'b01010110011011: color_data = 12'b101000000000;
		14'b01010110011100: color_data = 12'b101000000000;
		14'b01010110011101: color_data = 12'b010100000000;
		14'b01010110011110: color_data = 12'b010100000000;
		14'b01010110100001: color_data = 12'b010100000000;
		14'b01010110100010: color_data = 12'b010100000000;
		14'b01010110100011: color_data = 12'b101000000000;
		14'b01010110100100: color_data = 12'b101000000000;
		14'b01010110100101: color_data = 12'b101000000000;
		14'b01010110100110: color_data = 12'b101000000000;
		14'b01010110100111: color_data = 12'b101000000000;
		14'b01010110101000: color_data = 12'b101000000000;
		14'b01010110101001: color_data = 12'b101000000000;
		14'b01010110101010: color_data = 12'b010100000000;
		14'b01010110101011: color_data = 12'b010100000000;
		14'b01010110101100: color_data = 12'b010100000000;
		14'b01010110101101: color_data = 12'b010100000000;
		14'b01010110101110: color_data = 12'b101000000000;
		14'b01010110101111: color_data = 12'b101000000000;
		14'b01010110110000: color_data = 12'b101000000000;
		14'b01010110110001: color_data = 12'b101000000000;
		14'b01010110110010: color_data = 12'b101000000000;
		14'b01010110110011: color_data = 12'b101000000000;
		14'b01010110110100: color_data = 12'b101000000000;
		14'b01010110110101: color_data = 12'b101000000000;
		14'b01010110110110: color_data = 12'b101000000000;
		14'b01010110110111: color_data = 12'b010100000000;
		14'b01010110111000: color_data = 12'b010100000000;
		14'b01010110111001: color_data = 12'b010100000000;
		14'b01010110111010: color_data = 12'b010100000000;
		14'b01010110111011: color_data = 12'b010100000000;
		14'b01010110111100: color_data = 12'b010100000000;
		14'b01010110111101: color_data = 12'b010100000000;
		14'b01010111010010: color_data = 12'b010100000000;
		14'b01010111010011: color_data = 12'b010100000000;
		14'b01010111010100: color_data = 12'b010100000000;
		14'b01010111010101: color_data = 12'b101000000000;
		14'b01010111010110: color_data = 12'b101000000000;
		14'b01010111010111: color_data = 12'b010100000000;
		14'b01010111011000: color_data = 12'b010100000000;
		14'b01010111011001: color_data = 12'b101000000000;
		14'b01010111011010: color_data = 12'b101000000000;
		14'b01010111011011: color_data = 12'b101000000000;
		14'b01010111011100: color_data = 12'b101000000000;
		14'b01010111011101: color_data = 12'b010100000000;
		14'b01011000010000: color_data = 12'b010100000000;
		14'b01011000010001: color_data = 12'b010100000000;
		14'b01011000010010: color_data = 12'b101000000000;
		14'b01011000010011: color_data = 12'b101000000000;
		14'b01011000010100: color_data = 12'b010100000000;
		14'b01011000011001: color_data = 12'b010100000000;
		14'b01011000011010: color_data = 12'b010100000000;
		14'b01011000011011: color_data = 12'b101000000000;
		14'b01011000011100: color_data = 12'b101000000000;
		14'b01011000011101: color_data = 12'b101000000000;
		14'b01011000011110: color_data = 12'b101000000000;
		14'b01011000011111: color_data = 12'b010100000000;
		14'b01011000100100: color_data = 12'b010100000000;
		14'b01011000100101: color_data = 12'b101000000000;
		14'b01011000100110: color_data = 12'b101000000000;
		14'b01011000100111: color_data = 12'b101000000000;
		14'b01011000101000: color_data = 12'b101000000000;
		14'b01011000101001: color_data = 12'b101000000000;
		14'b01011000101010: color_data = 12'b101000000000;
		14'b01011000101011: color_data = 12'b101000000000;
		14'b01011000101100: color_data = 12'b010100000000;
		14'b01011000101101: color_data = 12'b010100000000;
		14'b01011000101110: color_data = 12'b101000000000;
		14'b01011000101111: color_data = 12'b101000000000;
		14'b01011000110000: color_data = 12'b101000000000;
		14'b01011000110001: color_data = 12'b101000000000;
		14'b01011000110010: color_data = 12'b101000000000;
		14'b01011000110011: color_data = 12'b101000000000;
		14'b01011000110100: color_data = 12'b101000000000;
		14'b01011000110101: color_data = 12'b101000000000;
		14'b01011000110110: color_data = 12'b010100000000;
		14'b01011000110111: color_data = 12'b010100000000;
		14'b01011000111000: color_data = 12'b010100000000;
		14'b01011000111001: color_data = 12'b010100000000;
		14'b01011000111010: color_data = 12'b010100000000;
		14'b01011001010101: color_data = 12'b010100000000;
		14'b01011001010110: color_data = 12'b010100000000;
		14'b01011001010111: color_data = 12'b010100000000;
		14'b01011001011000: color_data = 12'b010100000000;
		14'b01011001011001: color_data = 12'b101000000000;
		14'b01011001011010: color_data = 12'b101000000000;
		14'b01011001011011: color_data = 12'b101000000000;
		14'b01011001011100: color_data = 12'b101000000000;
		14'b01011001011101: color_data = 12'b101000000000;
		14'b01011001011110: color_data = 12'b010100000000;
		14'b01011010010010: color_data = 12'b010100000000;
		14'b01011010010011: color_data = 12'b101000000000;
		14'b01011010010100: color_data = 12'b101000000000;
		14'b01011010010101: color_data = 12'b010100000000;
		14'b01011010011011: color_data = 12'b010100000000;
		14'b01011010011100: color_data = 12'b101000000000;
		14'b01011010011101: color_data = 12'b101000000000;
		14'b01011010011110: color_data = 12'b101000000000;
		14'b01011010011111: color_data = 12'b101000000000;
		14'b01011010100000: color_data = 12'b101000000000;
		14'b01011010100001: color_data = 12'b010100000000;
		14'b01011010100101: color_data = 12'b010100000000;
		14'b01011010100110: color_data = 12'b101000000000;
		14'b01011010100111: color_data = 12'b101000000000;
		14'b01011010101000: color_data = 12'b101000000000;
		14'b01011010101001: color_data = 12'b101000000000;
		14'b01011010101010: color_data = 12'b101000000000;
		14'b01011010101011: color_data = 12'b101000000000;
		14'b01011010101100: color_data = 12'b101000000000;
		14'b01011010101101: color_data = 12'b101000000000;
		14'b01011010101110: color_data = 12'b101000000000;
		14'b01011010101111: color_data = 12'b101000000000;
		14'b01011010110000: color_data = 12'b101000000000;
		14'b01011010110001: color_data = 12'b101000000000;
		14'b01011010110010: color_data = 12'b101000000000;
		14'b01011010110011: color_data = 12'b101000000000;
		14'b01011010110100: color_data = 12'b010100000000;
		14'b01011010110101: color_data = 12'b010100000000;
		14'b01011010110110: color_data = 12'b010100000000;
		14'b01011010110111: color_data = 12'b010100000000;
		14'b01011010111000: color_data = 12'b010100000000;
		14'b01011010111001: color_data = 12'b010100000000;
		14'b01011011010111: color_data = 12'b010100000000;
		14'b01011011011000: color_data = 12'b010100000000;
		14'b01011011011001: color_data = 12'b010100000000;
		14'b01011011011010: color_data = 12'b101000000000;
		14'b01011011011011: color_data = 12'b101000000000;
		14'b01011011011100: color_data = 12'b101000000000;
		14'b01011011011101: color_data = 12'b101000000000;
		14'b01011011011110: color_data = 12'b101000000000;
		14'b01011011011111: color_data = 12'b010100000000;
		14'b01011100010011: color_data = 12'b010100000000;
		14'b01011100010100: color_data = 12'b101000000000;
		14'b01011100010101: color_data = 12'b101000000000;
		14'b01011100010110: color_data = 12'b101000000000;
		14'b01011100010111: color_data = 12'b010100000000;
		14'b01011100011100: color_data = 12'b010100000000;
		14'b01011100011101: color_data = 12'b101000000000;
		14'b01011100011110: color_data = 12'b101000000000;
		14'b01011100011111: color_data = 12'b101000000000;
		14'b01011100100000: color_data = 12'b101000000000;
		14'b01011100100001: color_data = 12'b101000000000;
		14'b01011100100010: color_data = 12'b010100000000;
		14'b01011100100111: color_data = 12'b010100000000;
		14'b01011100101000: color_data = 12'b101000000000;
		14'b01011100101001: color_data = 12'b101000000000;
		14'b01011100101010: color_data = 12'b101000000000;
		14'b01011100101011: color_data = 12'b101000000000;
		14'b01011100101100: color_data = 12'b101000000000;
		14'b01011100101101: color_data = 12'b101000000000;
		14'b01011100101110: color_data = 12'b101000000000;
		14'b01011100101111: color_data = 12'b101000000000;
		14'b01011100110000: color_data = 12'b101000000000;
		14'b01011100110001: color_data = 12'b101000000000;
		14'b01011100110010: color_data = 12'b010100000000;
		14'b01011100110011: color_data = 12'b010100000000;
		14'b01011100110100: color_data = 12'b010100000000;
		14'b01011100110101: color_data = 12'b010100000000;
		14'b01011100110110: color_data = 12'b010100000000;
		14'b01011100110111: color_data = 12'b010100000000;
		14'b01011100111000: color_data = 12'b010100000000;
		14'b01011101011001: color_data = 12'b010100000000;
		14'b01011101011010: color_data = 12'b010100000000;
		14'b01011101011011: color_data = 12'b101000000000;
		14'b01011101011100: color_data = 12'b101000000000;
		14'b01011101011101: color_data = 12'b101000000000;
		14'b01011101011110: color_data = 12'b101000000000;
		14'b01011101011111: color_data = 12'b101000000000;
		14'b01011110010100: color_data = 12'b010100000000;
		14'b01011110010101: color_data = 12'b101000000000;
		14'b01011110010110: color_data = 12'b101000000000;
		14'b01011110010111: color_data = 12'b101000000000;
		14'b01011110011000: color_data = 12'b010100000000;
		14'b01011110011101: color_data = 12'b010100000000;
		14'b01011110011110: color_data = 12'b101000000000;
		14'b01011110011111: color_data = 12'b101000000000;
		14'b01011110100000: color_data = 12'b101000000000;
		14'b01011110100001: color_data = 12'b101000000000;
		14'b01011110100010: color_data = 12'b101000000000;
		14'b01011110100011: color_data = 12'b010100000000;
		14'b01011110100101: color_data = 12'b010100000000;
		14'b01011110101000: color_data = 12'b010100000000;
		14'b01011110101001: color_data = 12'b101000000000;
		14'b01011110101010: color_data = 12'b101000000000;
		14'b01011110101011: color_data = 12'b101000000000;
		14'b01011110101100: color_data = 12'b101000000000;
		14'b01011110101101: color_data = 12'b101000000000;
		14'b01011110101110: color_data = 12'b010100000000;
		14'b01011110101111: color_data = 12'b010100000000;
		14'b01011110110000: color_data = 12'b010100000000;
		14'b01011110110011: color_data = 12'b010100000000;
		14'b01011110110100: color_data = 12'b010100000000;
		14'b01011110110101: color_data = 12'b010100000000;
		14'b01011110110110: color_data = 12'b010100000000;
		14'b01011110110111: color_data = 12'b010100000000;
		14'b01011110111000: color_data = 12'b010100000000;
		14'b01011111000001: color_data = 12'b010100000000;
		14'b01011111000010: color_data = 12'b010100000000;
		14'b01011111011010: color_data = 12'b010100000000;
		14'b01011111011011: color_data = 12'b010100000000;
		14'b01011111011100: color_data = 12'b101000000000;
		14'b01011111011101: color_data = 12'b101000000000;
		14'b01011111011110: color_data = 12'b101000000000;
		14'b01011111011111: color_data = 12'b101000000000;
		14'b01011111100000: color_data = 12'b101000000000;
		14'b01011111100110: color_data = 12'b010100000000;
		14'b01011111100111: color_data = 12'b010100000000;
		14'b01100000010101: color_data = 12'b010100000000;
		14'b01100000010110: color_data = 12'b101000000000;
		14'b01100000010111: color_data = 12'b101000000000;
		14'b01100000011000: color_data = 12'b101000000000;
		14'b01100000011001: color_data = 12'b010100000000;
		14'b01100000011110: color_data = 12'b101000000000;
		14'b01100000011111: color_data = 12'b101000000000;
		14'b01100000100000: color_data = 12'b101000000000;
		14'b01100000100001: color_data = 12'b101000000000;
		14'b01100000100010: color_data = 12'b101000000000;
		14'b01100000100011: color_data = 12'b101000000000;
		14'b01100000100100: color_data = 12'b010100000000;
		14'b01100000100101: color_data = 12'b010100000000;
		14'b01100000100110: color_data = 12'b010100000000;
		14'b01100000101010: color_data = 12'b101000000000;
		14'b01100000101011: color_data = 12'b101000000000;
		14'b01100000101100: color_data = 12'b101000000000;
		14'b01100000101101: color_data = 12'b010100000000;
		14'b01100000110010: color_data = 12'b010100000000;
		14'b01100000110011: color_data = 12'b010100000000;
		14'b01100000110100: color_data = 12'b010100000000;
		14'b01100000110101: color_data = 12'b010100000000;
		14'b01100001000101: color_data = 12'b010100000000;
		14'b01100001011011: color_data = 12'b010100000000;
		14'b01100001011100: color_data = 12'b010100000000;
		14'b01100001011101: color_data = 12'b101000000000;
		14'b01100001011110: color_data = 12'b101000000000;
		14'b01100001011111: color_data = 12'b101000000000;
		14'b01100001100000: color_data = 12'b101000000000;
		14'b01100001100001: color_data = 12'b010100000000;
		14'b01100001100111: color_data = 12'b010100000000;
		14'b01100010010110: color_data = 12'b010100000000;
		14'b01100010010111: color_data = 12'b010100000000;
		14'b01100010011000: color_data = 12'b101000000000;
		14'b01100010011001: color_data = 12'b101000000000;
		14'b01100010011010: color_data = 12'b010100000000;
		14'b01100010011110: color_data = 12'b010100000000;
		14'b01100010011111: color_data = 12'b101000000000;
		14'b01100010100000: color_data = 12'b101000000000;
		14'b01100010100001: color_data = 12'b101000000000;
		14'b01100010100010: color_data = 12'b101000000000;
		14'b01100010100011: color_data = 12'b101000000000;
		14'b01100010100100: color_data = 12'b101000000000;
		14'b01100010100101: color_data = 12'b101000000000;
		14'b01100010100110: color_data = 12'b010100000000;
		14'b01100010100111: color_data = 12'b010100000000;
		14'b01100010101011: color_data = 12'b010100000000;
		14'b01100010110000: color_data = 12'b010100000000;
		14'b01100010110001: color_data = 12'b010100000000;
		14'b01100010110010: color_data = 12'b010100000000;
		14'b01100010110011: color_data = 12'b010100000000;
		14'b01100010110100: color_data = 12'b010100000000;
		14'b01100011000111: color_data = 12'b010100000000;
		14'b01100011001000: color_data = 12'b010100000000;
		14'b01100011011100: color_data = 12'b010100000000;
		14'b01100011011101: color_data = 12'b010100000000;
		14'b01100011011110: color_data = 12'b101000000000;
		14'b01100011011111: color_data = 12'b101000000000;
		14'b01100011100000: color_data = 12'b101000000000;
		14'b01100011100001: color_data = 12'b101000000000;
		14'b01100011100010: color_data = 12'b010100000000;
		14'b01100011101000: color_data = 12'b010100000000;
		14'b01100100011000: color_data = 12'b010100000000;
		14'b01100100011001: color_data = 12'b101000000000;
		14'b01100100011010: color_data = 12'b101000000000;
		14'b01100100011011: color_data = 12'b010100000000;
		14'b01100100011111: color_data = 12'b010100000000;
		14'b01100100100000: color_data = 12'b101000000000;
		14'b01100100100001: color_data = 12'b101000000000;
		14'b01100100100010: color_data = 12'b101000000000;
		14'b01100100100011: color_data = 12'b101000000000;
		14'b01100100100100: color_data = 12'b101000000000;
		14'b01100100100101: color_data = 12'b101000000000;
		14'b01100100100110: color_data = 12'b101000000000;
		14'b01100100100111: color_data = 12'b010100000000;
		14'b01100100101000: color_data = 12'b010100000000;
		14'b01100100101111: color_data = 12'b010100000000;
		14'b01100100110000: color_data = 12'b010100000000;
		14'b01100100110001: color_data = 12'b101000000000;
		14'b01100100110010: color_data = 12'b010100000000;
		14'b01100101001000: color_data = 12'b010100000000;
		14'b01100101001001: color_data = 12'b010100000000;
		14'b01100101001010: color_data = 12'b010100000000;
		14'b01100101011101: color_data = 12'b010100000000;
		14'b01100101011110: color_data = 12'b010100000000;
		14'b01100101011111: color_data = 12'b101000000000;
		14'b01100101100000: color_data = 12'b101000000000;
		14'b01100101100001: color_data = 12'b101000000000;
		14'b01100101100010: color_data = 12'b101000000000;
		14'b01100101100011: color_data = 12'b010100000000;
		14'b01100101101001: color_data = 12'b010100000000;
		14'b01100110011001: color_data = 12'b010100000000;
		14'b01100110011010: color_data = 12'b101000000000;
		14'b01100110011011: color_data = 12'b101000000000;
		14'b01100110011100: color_data = 12'b010100000000;
		14'b01100110100000: color_data = 12'b010100000000;
		14'b01100110100001: color_data = 12'b101000000000;
		14'b01100110100010: color_data = 12'b101000000000;
		14'b01100110100011: color_data = 12'b101000000000;
		14'b01100110100100: color_data = 12'b101000000000;
		14'b01100110100101: color_data = 12'b101000000000;
		14'b01100110100110: color_data = 12'b101000000000;
		14'b01100110100111: color_data = 12'b010100000000;
		14'b01100110101000: color_data = 12'b010100000000;
		14'b01100110101001: color_data = 12'b010100000000;
		14'b01100110101010: color_data = 12'b010100000000;
		14'b01100110101011: color_data = 12'b010100000000;
		14'b01100110101100: color_data = 12'b010100000000;
		14'b01100110101101: color_data = 12'b010100000000;
		14'b01100110101110: color_data = 12'b010100000000;
		14'b01100110101111: color_data = 12'b101000000000;
		14'b01100110110000: color_data = 12'b101000000000;
		14'b01100110110001: color_data = 12'b010100000000;
		14'b01100111001001: color_data = 12'b010100000000;
		14'b01100111001010: color_data = 12'b010100000000;
		14'b01100111001011: color_data = 12'b010100000000;
		14'b01100111011110: color_data = 12'b010100000000;
		14'b01100111011111: color_data = 12'b010100000000;
		14'b01100111100000: color_data = 12'b101000000000;
		14'b01100111100001: color_data = 12'b101000000000;
		14'b01100111100010: color_data = 12'b101000000000;
		14'b01100111100011: color_data = 12'b101000000000;
		14'b01100111100100: color_data = 12'b101000000000;
		14'b01100111101001: color_data = 12'b010100000000;
		14'b01100111101010: color_data = 12'b010100000000;
		14'b01101000011010: color_data = 12'b010100000000;
		14'b01101000011011: color_data = 12'b101000000000;
		14'b01101000011100: color_data = 12'b101000000000;
		14'b01101000100001: color_data = 12'b010100000000;
		14'b01101000100010: color_data = 12'b101000000000;
		14'b01101000100011: color_data = 12'b101000000000;
		14'b01101000100100: color_data = 12'b101000000000;
		14'b01101000100101: color_data = 12'b101000000000;
		14'b01101000100110: color_data = 12'b101000000000;
		14'b01101000100111: color_data = 12'b010100000000;
		14'b01101000101000: color_data = 12'b010100000000;
		14'b01101000101001: color_data = 12'b010100000000;
		14'b01101000101010: color_data = 12'b010100000000;
		14'b01101000101011: color_data = 12'b010100000000;
		14'b01101000101100: color_data = 12'b010100000000;
		14'b01101000101101: color_data = 12'b010100000000;
		14'b01101000101110: color_data = 12'b101000000000;
		14'b01101000101111: color_data = 12'b101000000000;
		14'b01101000110000: color_data = 12'b101000000000;
		14'b01101001000100: color_data = 12'b010100000000;
		14'b01101001001001: color_data = 12'b010100000000;
		14'b01101001001010: color_data = 12'b010100000000;
		14'b01101001001011: color_data = 12'b010100000000;
		14'b01101001100000: color_data = 12'b010100000000;
		14'b01101001100001: color_data = 12'b101000000000;
		14'b01101001100010: color_data = 12'b101000000000;
		14'b01101001100011: color_data = 12'b101000000000;
		14'b01101001100100: color_data = 12'b101000000000;
		14'b01101001100101: color_data = 12'b101000000000;
		14'b01101001100110: color_data = 12'b010100000000;
		14'b01101001101010: color_data = 12'b010100000000;
		14'b01101010011011: color_data = 12'b010100000000;
		14'b01101010011100: color_data = 12'b101000000000;
		14'b01101010011101: color_data = 12'b010100000000;
		14'b01101010100010: color_data = 12'b101000000000;
		14'b01101010100011: color_data = 12'b101000000000;
		14'b01101010100100: color_data = 12'b101000000000;
		14'b01101010100101: color_data = 12'b101000000000;
		14'b01101010100110: color_data = 12'b101000000000;
		14'b01101010100111: color_data = 12'b101000000000;
		14'b01101010101000: color_data = 12'b010100000000;
		14'b01101010101001: color_data = 12'b010100000000;
		14'b01101010101010: color_data = 12'b010100000000;
		14'b01101010101011: color_data = 12'b010100000000;
		14'b01101010101100: color_data = 12'b010100000000;
		14'b01101010101101: color_data = 12'b010100000000;
		14'b01101010101110: color_data = 12'b101000000000;
		14'b01101010101111: color_data = 12'b101000000000;
		14'b01101010110000: color_data = 12'b010100000000;
		14'b01101010111000: color_data = 12'b010100000000;
		14'b01101010111001: color_data = 12'b010100000000;
		14'b01101010111010: color_data = 12'b010100000000;
		14'b01101010111011: color_data = 12'b010100000000;
		14'b01101010111100: color_data = 12'b010100000000;
		14'b01101010111101: color_data = 12'b010100000000;
		14'b01101010111110: color_data = 12'b010100000000;
		14'b01101010111111: color_data = 12'b010100000000;
		14'b01101011000000: color_data = 12'b010100000000;
		14'b01101011000010: color_data = 12'b010100000000;
		14'b01101011000011: color_data = 12'b010100000000;
		14'b01101011000100: color_data = 12'b010100000000;
		14'b01101011000101: color_data = 12'b010100000000;
		14'b01101011000110: color_data = 12'b010100000000;
		14'b01101011000111: color_data = 12'b010100000000;
		14'b01101011001000: color_data = 12'b010100000000;
		14'b01101011001001: color_data = 12'b010100000000;
		14'b01101011001010: color_data = 12'b010100000000;
		14'b01101011001011: color_data = 12'b010100000000;
		14'b01101011001100: color_data = 12'b010100000000;
		14'b01101011100001: color_data = 12'b010100000000;
		14'b01101011100010: color_data = 12'b101000000000;
		14'b01101011100011: color_data = 12'b101000000000;
		14'b01101011100100: color_data = 12'b101000000000;
		14'b01101011100101: color_data = 12'b101000000000;
		14'b01101011100110: color_data = 12'b101000000000;
		14'b01101011100111: color_data = 12'b010100000000;
		14'b01101100011100: color_data = 12'b010100000000;
		14'b01101100011101: color_data = 12'b010100000000;
		14'b01101100100010: color_data = 12'b101000000000;
		14'b01101100100011: color_data = 12'b101000000000;
		14'b01101100100100: color_data = 12'b101000000000;
		14'b01101100100101: color_data = 12'b101000000000;
		14'b01101100100110: color_data = 12'b101000000000;
		14'b01101100100111: color_data = 12'b101000000000;
		14'b01101100101000: color_data = 12'b101000000000;
		14'b01101100101001: color_data = 12'b010100000000;
		14'b01101100101010: color_data = 12'b010100000000;
		14'b01101100101011: color_data = 12'b010100000000;
		14'b01101100101100: color_data = 12'b010100000000;
		14'b01101100101101: color_data = 12'b101000000000;
		14'b01101100101110: color_data = 12'b101000000000;
		14'b01101100101111: color_data = 12'b010100000000;
		14'b01101100111011: color_data = 12'b010100000000;
		14'b01101100111100: color_data = 12'b010100000000;
		14'b01101100111101: color_data = 12'b010100000000;
		14'b01101100111110: color_data = 12'b010100000000;
		14'b01101100111111: color_data = 12'b010100000000;
		14'b01101101000000: color_data = 12'b010100000000;
		14'b01101101000001: color_data = 12'b010100000000;
		14'b01101101000010: color_data = 12'b010100000000;
		14'b01101101000011: color_data = 12'b101000000000;
		14'b01101101000100: color_data = 12'b101000000000;
		14'b01101101000101: color_data = 12'b010100000000;
		14'b01101101000110: color_data = 12'b101000000000;
		14'b01101101000111: color_data = 12'b101000000000;
		14'b01101101001000: color_data = 12'b010100000000;
		14'b01101101001001: color_data = 12'b010100000000;
		14'b01101101001010: color_data = 12'b010100000000;
		14'b01101101001011: color_data = 12'b010100000000;
		14'b01101101001100: color_data = 12'b010100000000;
		14'b01101101100001: color_data = 12'b010100000000;
		14'b01101101100010: color_data = 12'b010100000000;
		14'b01101101100011: color_data = 12'b101000000000;
		14'b01101101100100: color_data = 12'b101000000000;
		14'b01101101100101: color_data = 12'b101000000000;
		14'b01101101100110: color_data = 12'b101000000000;
		14'b01101101100111: color_data = 12'b101000000000;
		14'b01101101101000: color_data = 12'b010100000000;
		14'b01101110011100: color_data = 12'b010100000000;
		14'b01101110011101: color_data = 12'b010100000000;
		14'b01101110100010: color_data = 12'b010100000000;
		14'b01101110100011: color_data = 12'b101000000000;
		14'b01101110100100: color_data = 12'b101000000000;
		14'b01101110100101: color_data = 12'b101000000000;
		14'b01101110100110: color_data = 12'b101000000000;
		14'b01101110100111: color_data = 12'b101000000000;
		14'b01101110101000: color_data = 12'b010100000000;
		14'b01101110101001: color_data = 12'b010100000000;
		14'b01101110101010: color_data = 12'b010100000000;
		14'b01101110101011: color_data = 12'b010100000000;
		14'b01101110101100: color_data = 12'b101000000000;
		14'b01101110101101: color_data = 12'b101000000000;
		14'b01101110101110: color_data = 12'b101000000000;
		14'b01101110101111: color_data = 12'b010100000000;
		14'b01101110111100: color_data = 12'b010100000000;
		14'b01101110111101: color_data = 12'b010100000000;
		14'b01101110111110: color_data = 12'b101000000000;
		14'b01101110111111: color_data = 12'b010100000000;
		14'b01101111000000: color_data = 12'b010100000000;
		14'b01101111000001: color_data = 12'b010100000000;
		14'b01101111000010: color_data = 12'b101000000000;
		14'b01101111000011: color_data = 12'b101000000000;
		14'b01101111000100: color_data = 12'b101000000000;
		14'b01101111000101: color_data = 12'b010100000000;
		14'b01101111000110: color_data = 12'b101000000000;
		14'b01101111000111: color_data = 12'b101000000000;
		14'b01101111001000: color_data = 12'b101000000000;
		14'b01101111001001: color_data = 12'b101000000000;
		14'b01101111001010: color_data = 12'b010100000000;
		14'b01101111001011: color_data = 12'b010100000000;
		14'b01101111001100: color_data = 12'b010100000000;
		14'b01101111100010: color_data = 12'b010100000000;
		14'b01101111100011: color_data = 12'b010100000000;
		14'b01101111100100: color_data = 12'b101000000000;
		14'b01101111100101: color_data = 12'b101000000000;
		14'b01101111100110: color_data = 12'b101000000000;
		14'b01101111100111: color_data = 12'b101000000000;
		14'b01101111101000: color_data = 12'b101000000000;
		14'b01101111101001: color_data = 12'b010100000000;
		14'b01110000011100: color_data = 12'b010100000000;
		14'b01110000011101: color_data = 12'b010100000000;
		14'b01110000100010: color_data = 12'b010100000000;
		14'b01110000100011: color_data = 12'b101000000000;
		14'b01110000100100: color_data = 12'b101000000000;
		14'b01110000100101: color_data = 12'b101000000000;
		14'b01110000100110: color_data = 12'b101000000000;
		14'b01110000100111: color_data = 12'b101000000000;
		14'b01110000101000: color_data = 12'b010100000000;
		14'b01110000101001: color_data = 12'b010100000000;
		14'b01110000101010: color_data = 12'b010100000000;
		14'b01110000101011: color_data = 12'b101000000000;
		14'b01110000101100: color_data = 12'b101000000000;
		14'b01110000101101: color_data = 12'b101000000000;
		14'b01110000101110: color_data = 12'b010100000000;
		14'b01110000111011: color_data = 12'b010100000000;
		14'b01110000111100: color_data = 12'b010100000000;
		14'b01110000111101: color_data = 12'b101000000000;
		14'b01110000111110: color_data = 12'b101000000000;
		14'b01110000111111: color_data = 12'b101000000000;
		14'b01110001000000: color_data = 12'b101000000000;
		14'b01110001000001: color_data = 12'b101000000000;
		14'b01110001000010: color_data = 12'b101000000000;
		14'b01110001000011: color_data = 12'b101000000000;
		14'b01110001000100: color_data = 12'b101000000000;
		14'b01110001000101: color_data = 12'b101000000000;
		14'b01110001000110: color_data = 12'b101000000000;
		14'b01110001000111: color_data = 12'b101000000000;
		14'b01110001001000: color_data = 12'b101000000000;
		14'b01110001001001: color_data = 12'b101000000000;
		14'b01110001001010: color_data = 12'b101000000000;
		14'b01110001001011: color_data = 12'b101000000000;
		14'b01110001001100: color_data = 12'b010100000000;
		14'b01110001001101: color_data = 12'b010100000000;
		14'b01110001100011: color_data = 12'b010100000000;
		14'b01110001100100: color_data = 12'b101000000000;
		14'b01110001100101: color_data = 12'b101000000000;
		14'b01110001100110: color_data = 12'b101000000000;
		14'b01110001100111: color_data = 12'b101000000000;
		14'b01110001101000: color_data = 12'b101000000000;
		14'b01110001101001: color_data = 12'b101000000000;
		14'b01110001101010: color_data = 12'b010100000000;
		14'b01110010011100: color_data = 12'b010100000000;
		14'b01110010011101: color_data = 12'b010100000000;
		14'b01110010100010: color_data = 12'b010100000000;
		14'b01110010100011: color_data = 12'b101000000000;
		14'b01110010100100: color_data = 12'b101000000000;
		14'b01110010100101: color_data = 12'b101000000000;
		14'b01110010100110: color_data = 12'b101000000000;
		14'b01110010100111: color_data = 12'b010100000000;
		14'b01110010101000: color_data = 12'b010100000000;
		14'b01110010101001: color_data = 12'b010100000000;
		14'b01110010101010: color_data = 12'b010100000000;
		14'b01110010101011: color_data = 12'b101000000000;
		14'b01110010101100: color_data = 12'b101000000000;
		14'b01110010101101: color_data = 12'b101000000000;
		14'b01110010101110: color_data = 12'b010100000000;
		14'b01110010111010: color_data = 12'b010100000000;
		14'b01110010111011: color_data = 12'b010100000000;
		14'b01110010111100: color_data = 12'b101000000000;
		14'b01110010111101: color_data = 12'b101000000000;
		14'b01110010111110: color_data = 12'b101000000000;
		14'b01110010111111: color_data = 12'b101000000000;
		14'b01110011000000: color_data = 12'b101000000000;
		14'b01110011000001: color_data = 12'b101000000000;
		14'b01110011000010: color_data = 12'b101000000000;
		14'b01110011000011: color_data = 12'b101000000000;
		14'b01110011000100: color_data = 12'b101000000000;
		14'b01110011000101: color_data = 12'b101000000000;
		14'b01110011000110: color_data = 12'b101000000000;
		14'b01110011000111: color_data = 12'b101000000000;
		14'b01110011001000: color_data = 12'b101000000000;
		14'b01110011001001: color_data = 12'b101000000000;
		14'b01110011001010: color_data = 12'b101000000000;
		14'b01110011001011: color_data = 12'b101000000000;
		14'b01110011001100: color_data = 12'b101000000000;
		14'b01110011001101: color_data = 12'b101000000000;
		14'b01110011001110: color_data = 12'b010100000000;
		14'b01110011100100: color_data = 12'b010100000000;
		14'b01110011100101: color_data = 12'b101000000000;
		14'b01110011100110: color_data = 12'b101000000000;
		14'b01110011100111: color_data = 12'b101000000000;
		14'b01110011101000: color_data = 12'b101000000000;
		14'b01110011101001: color_data = 12'b101000000000;
		14'b01110011101010: color_data = 12'b101000000000;
		14'b01110100011100: color_data = 12'b010100000000;
		14'b01110100011101: color_data = 12'b010100000000;
		14'b01110100100010: color_data = 12'b010100000000;
		14'b01110100100011: color_data = 12'b101000000000;
		14'b01110100100100: color_data = 12'b101000000000;
		14'b01110100100101: color_data = 12'b101000000000;
		14'b01110100100110: color_data = 12'b101000000000;
		14'b01110100100111: color_data = 12'b010100000000;
		14'b01110100101000: color_data = 12'b010100000000;
		14'b01110100101001: color_data = 12'b010100000000;
		14'b01110100101010: color_data = 12'b101000000000;
		14'b01110100101011: color_data = 12'b101000000000;
		14'b01110100101100: color_data = 12'b101000000000;
		14'b01110100101101: color_data = 12'b010100000000;
		14'b01110100111001: color_data = 12'b010100000000;
		14'b01110100111010: color_data = 12'b101000000000;
		14'b01110100111011: color_data = 12'b101000000000;
		14'b01110100111100: color_data = 12'b101000000000;
		14'b01110100111101: color_data = 12'b101000000000;
		14'b01110100111110: color_data = 12'b101000000000;
		14'b01110100111111: color_data = 12'b101000000000;
		14'b01110101000000: color_data = 12'b101000000000;
		14'b01110101000001: color_data = 12'b101000000000;
		14'b01110101000010: color_data = 12'b101000000000;
		14'b01110101000011: color_data = 12'b101000000000;
		14'b01110101000100: color_data = 12'b101000000000;
		14'b01110101000101: color_data = 12'b101000000000;
		14'b01110101000110: color_data = 12'b101000000000;
		14'b01110101000111: color_data = 12'b101000000000;
		14'b01110101001000: color_data = 12'b010100000000;
		14'b01110101001001: color_data = 12'b101000000000;
		14'b01110101001010: color_data = 12'b101000000000;
		14'b01110101001011: color_data = 12'b101000000000;
		14'b01110101001100: color_data = 12'b101000000000;
		14'b01110101001101: color_data = 12'b101000000000;
		14'b01110101001110: color_data = 12'b010100000000;
		14'b01110101001111: color_data = 12'b010100000000;
		14'b01110101100100: color_data = 12'b010100000000;
		14'b01110101100101: color_data = 12'b010100000000;
		14'b01110101100110: color_data = 12'b101000000000;
		14'b01110101100111: color_data = 12'b101000000000;
		14'b01110101101000: color_data = 12'b101000000000;
		14'b01110101101001: color_data = 12'b101000000000;
		14'b01110101101010: color_data = 12'b101000000000;
		14'b01110110011100: color_data = 12'b010100000000;
		14'b01110110011101: color_data = 12'b010100000000;
		14'b01110110011110: color_data = 12'b010100000000;
		14'b01110110100010: color_data = 12'b010100000000;
		14'b01110110100011: color_data = 12'b101000000000;
		14'b01110110100100: color_data = 12'b101000000000;
		14'b01110110100101: color_data = 12'b101000000000;
		14'b01110110100110: color_data = 12'b101000000000;
		14'b01110110100111: color_data = 12'b010100000000;
		14'b01110110101000: color_data = 12'b010100000000;
		14'b01110110101001: color_data = 12'b101000000000;
		14'b01110110101010: color_data = 12'b101000000000;
		14'b01110110101011: color_data = 12'b101000000000;
		14'b01110110101100: color_data = 12'b101000000000;
		14'b01110110101101: color_data = 12'b010100000000;
		14'b01110110111000: color_data = 12'b010100000000;
		14'b01110110111001: color_data = 12'b101000000000;
		14'b01110110111010: color_data = 12'b101000000000;
		14'b01110110111011: color_data = 12'b010100000000;
		14'b01110110111100: color_data = 12'b101000000000;
		14'b01110110111101: color_data = 12'b101000000000;
		14'b01110110111110: color_data = 12'b101000000000;
		14'b01110110111111: color_data = 12'b101000000000;
		14'b01110111000000: color_data = 12'b101000000000;
		14'b01110111000001: color_data = 12'b010100000000;
		14'b01110111000010: color_data = 12'b010100000000;
		14'b01110111000011: color_data = 12'b010100000000;
		14'b01110111000100: color_data = 12'b010100000000;
		14'b01110111000101: color_data = 12'b101000000000;
		14'b01110111000110: color_data = 12'b101000000000;
		14'b01110111000111: color_data = 12'b101000000000;
		14'b01110111001000: color_data = 12'b010100000000;
		14'b01110111001001: color_data = 12'b010100000000;
		14'b01110111001010: color_data = 12'b010100000000;
		14'b01110111001011: color_data = 12'b101000000000;
		14'b01110111001100: color_data = 12'b101000000000;
		14'b01110111001101: color_data = 12'b101000000000;
		14'b01110111001110: color_data = 12'b101000000000;
		14'b01110111001111: color_data = 12'b010100000000;
		14'b01110111100101: color_data = 12'b010100000000;
		14'b01110111100110: color_data = 12'b101000000000;
		14'b01110111100111: color_data = 12'b101000000000;
		14'b01110111101000: color_data = 12'b101000000000;
		14'b01110111101001: color_data = 12'b101000000000;
		14'b01110111101010: color_data = 12'b101000000000;
		14'b01111000011100: color_data = 12'b010100000000;
		14'b01111000011101: color_data = 12'b010100000000;
		14'b01111000011110: color_data = 12'b010100000000;
		14'b01111000100010: color_data = 12'b010100000000;
		14'b01111000100011: color_data = 12'b101000000000;
		14'b01111000100100: color_data = 12'b101000000000;
		14'b01111000100101: color_data = 12'b101000000000;
		14'b01111000100110: color_data = 12'b101000000000;
		14'b01111000100111: color_data = 12'b010100000000;
		14'b01111000101000: color_data = 12'b010100000000;
		14'b01111000101001: color_data = 12'b101000000000;
		14'b01111000101010: color_data = 12'b101000000000;
		14'b01111000101011: color_data = 12'b101000000000;
		14'b01111000101100: color_data = 12'b010100000000;
		14'b01111000110111: color_data = 12'b010100000000;
		14'b01111000111000: color_data = 12'b010100000000;
		14'b01111000111001: color_data = 12'b010100000000;
		14'b01111000111010: color_data = 12'b010100000000;
		14'b01111000111011: color_data = 12'b010100000000;
		14'b01111000111100: color_data = 12'b010100000000;
		14'b01111000111101: color_data = 12'b101000000000;
		14'b01111000111110: color_data = 12'b101000000000;
		14'b01111000111111: color_data = 12'b101000000000;
		14'b01111001000000: color_data = 12'b010100000000;
		14'b01111001000101: color_data = 12'b010100000000;
		14'b01111001000110: color_data = 12'b101000000000;
		14'b01111001000111: color_data = 12'b101000000000;
		14'b01111001001000: color_data = 12'b010100000000;
		14'b01111001001011: color_data = 12'b010100000000;
		14'b01111001001100: color_data = 12'b010100000000;
		14'b01111001001101: color_data = 12'b101000000000;
		14'b01111001001110: color_data = 12'b101000000000;
		14'b01111001001111: color_data = 12'b101000000000;
		14'b01111001010000: color_data = 12'b010100000000;
		14'b01111001100101: color_data = 12'b010100000000;
		14'b01111001100110: color_data = 12'b010100000000;
		14'b01111001100111: color_data = 12'b101000000000;
		14'b01111001101000: color_data = 12'b101000000000;
		14'b01111001101001: color_data = 12'b101000000000;
		14'b01111001101010: color_data = 12'b101000000000;
		14'b01111010011100: color_data = 12'b010100000000;
		14'b01111010011101: color_data = 12'b010100000000;
		14'b01111010100010: color_data = 12'b010100000000;
		14'b01111010100011: color_data = 12'b101000000000;
		14'b01111010100100: color_data = 12'b101000000000;
		14'b01111010100101: color_data = 12'b010100000000;
		14'b01111010100110: color_data = 12'b010100000000;
		14'b01111010100111: color_data = 12'b010100000000;
		14'b01111010101000: color_data = 12'b010100000000;
		14'b01111010101001: color_data = 12'b101000000000;
		14'b01111010101010: color_data = 12'b101000000000;
		14'b01111010101011: color_data = 12'b101000000000;
		14'b01111010101100: color_data = 12'b010100000000;
		14'b01111010110111: color_data = 12'b010100000000;
		14'b01111010111000: color_data = 12'b010100000000;
		14'b01111010111010: color_data = 12'b010100000000;
		14'b01111010111011: color_data = 12'b010100000000;
		14'b01111010111100: color_data = 12'b010100000000;
		14'b01111010111101: color_data = 12'b101000000000;
		14'b01111010111110: color_data = 12'b101000000000;
		14'b01111010111111: color_data = 12'b010100000000;
		14'b01111011000101: color_data = 12'b010100000000;
		14'b01111011000110: color_data = 12'b101000000000;
		14'b01111011000111: color_data = 12'b101000000000;
		14'b01111011001000: color_data = 12'b101000000000;
		14'b01111011001001: color_data = 12'b010100000000;
		14'b01111011001101: color_data = 12'b010100000000;
		14'b01111011001110: color_data = 12'b101000000000;
		14'b01111011001111: color_data = 12'b101000000000;
		14'b01111011010000: color_data = 12'b101000000000;
		14'b01111011010001: color_data = 12'b010100000000;
		14'b01111011100110: color_data = 12'b010100000000;
		14'b01111011100111: color_data = 12'b101000000000;
		14'b01111011101000: color_data = 12'b101000000000;
		14'b01111011101001: color_data = 12'b101000000000;
		14'b01111011101010: color_data = 12'b101000000000;
		14'b01111100011011: color_data = 12'b010100000000;
		14'b01111100011100: color_data = 12'b010100000000;
		14'b01111100100010: color_data = 12'b101000000000;
		14'b01111100100011: color_data = 12'b101000000000;
		14'b01111100100100: color_data = 12'b010100000000;
		14'b01111100100101: color_data = 12'b010100000000;
		14'b01111100100110: color_data = 12'b010100000000;
		14'b01111100100111: color_data = 12'b010100000000;
		14'b01111100101000: color_data = 12'b010100000000;
		14'b01111100101001: color_data = 12'b101000000000;
		14'b01111100101010: color_data = 12'b101000000000;
		14'b01111100101011: color_data = 12'b010100000000;
		14'b01111100110110: color_data = 12'b010100000000;
		14'b01111100110111: color_data = 12'b010100000000;
		14'b01111100111010: color_data = 12'b010100000000;
		14'b01111100111011: color_data = 12'b010100000000;
		14'b01111100111100: color_data = 12'b101000000000;
		14'b01111100111101: color_data = 12'b101000000000;
		14'b01111100111110: color_data = 12'b010100000000;
		14'b01111101000100: color_data = 12'b010100000000;
		14'b01111101000101: color_data = 12'b010100000000;
		14'b01111101000110: color_data = 12'b101000000000;
		14'b01111101000111: color_data = 12'b101000000000;
		14'b01111101001000: color_data = 12'b101000000000;
		14'b01111101001001: color_data = 12'b101000000000;
		14'b01111101001010: color_data = 12'b010100000000;
		14'b01111101001110: color_data = 12'b010100000000;
		14'b01111101001111: color_data = 12'b101000000000;
		14'b01111101010000: color_data = 12'b101000000000;
		14'b01111101010001: color_data = 12'b010100000000;
		14'b01111101010010: color_data = 12'b010100000000;
		14'b01111101100111: color_data = 12'b010100000000;
		14'b01111101101000: color_data = 12'b101000000000;
		14'b01111101101001: color_data = 12'b101000000000;
		14'b01111101101010: color_data = 12'b101000000000;
		14'b01111101101011: color_data = 12'b010100000000;
		14'b01111110100001: color_data = 12'b010100000000;
		14'b01111110100010: color_data = 12'b010100000000;
		14'b01111110100011: color_data = 12'b010100000000;
		14'b01111110100100: color_data = 12'b010100000000;
		14'b01111110100101: color_data = 12'b010100000000;
		14'b01111110100110: color_data = 12'b010100000000;
		14'b01111110100111: color_data = 12'b010100000000;
		14'b01111110101000: color_data = 12'b101000000000;
		14'b01111110101001: color_data = 12'b101000000000;
		14'b01111110101010: color_data = 12'b101000000000;
		14'b01111110101011: color_data = 12'b010100000000;
		14'b01111110110110: color_data = 12'b010100000000;
		14'b01111110111010: color_data = 12'b010100000000;
		14'b01111110111011: color_data = 12'b101000000000;
		14'b01111110111100: color_data = 12'b101000000000;
		14'b01111110111101: color_data = 12'b010100000000;
		14'b01111111000001: color_data = 12'b010100000000;
		14'b01111111000010: color_data = 12'b010100000000;
		14'b01111111000011: color_data = 12'b010100000000;
		14'b01111111000100: color_data = 12'b101000000000;
		14'b01111111000101: color_data = 12'b101000000000;
		14'b01111111000110: color_data = 12'b101000000000;
		14'b01111111000111: color_data = 12'b101000000000;
		14'b01111111001000: color_data = 12'b101000000000;
		14'b01111111001001: color_data = 12'b101000000000;
		14'b01111111001010: color_data = 12'b101000000000;
		14'b01111111001011: color_data = 12'b010100000000;
		14'b01111111001111: color_data = 12'b010100000000;
		14'b01111111010000: color_data = 12'b010100000000;
		14'b01111111010001: color_data = 12'b010100000000;
		14'b01111111010010: color_data = 12'b010100000000;
		14'b01111111100111: color_data = 12'b010100000000;
		14'b01111111101000: color_data = 12'b101000000000;
		14'b01111111101001: color_data = 12'b101000000000;
		14'b01111111101010: color_data = 12'b101000000000;
		14'b01111111101011: color_data = 12'b101000000000;
		14'b10000000100000: color_data = 12'b010100000000;
		14'b10000000100001: color_data = 12'b010100000000;
		14'b10000000100010: color_data = 12'b010100000000;
		14'b10000000100011: color_data = 12'b010100000000;
		14'b10000000100100: color_data = 12'b101000000000;
		14'b10000000100101: color_data = 12'b010100000000;
		14'b10000000100110: color_data = 12'b010100000000;
		14'b10000000100111: color_data = 12'b010100000000;
		14'b10000000101000: color_data = 12'b101000000000;
		14'b10000000101001: color_data = 12'b101000000000;
		14'b10000000101010: color_data = 12'b010100000000;
		14'b10000000101011: color_data = 12'b010100000000;
		14'b10000000111001: color_data = 12'b010100000000;
		14'b10000000111010: color_data = 12'b010100000000;
		14'b10000000111011: color_data = 12'b010100000000;
		14'b10000000111100: color_data = 12'b010100000000;
		14'b10000000111101: color_data = 12'b010100000000;
		14'b10000000111110: color_data = 12'b010100000000;
		14'b10000000111111: color_data = 12'b010100000000;
		14'b10000001000000: color_data = 12'b101000000000;
		14'b10000001000001: color_data = 12'b101000000000;
		14'b10000001000010: color_data = 12'b101000000000;
		14'b10000001000011: color_data = 12'b101000000000;
		14'b10000001000100: color_data = 12'b101000000000;
		14'b10000001000101: color_data = 12'b101000000000;
		14'b10000001000110: color_data = 12'b101000000000;
		14'b10000001000111: color_data = 12'b101000000000;
		14'b10000001001000: color_data = 12'b101000000000;
		14'b10000001001001: color_data = 12'b101000000000;
		14'b10000001001010: color_data = 12'b101000000000;
		14'b10000001001011: color_data = 12'b101000000000;
		14'b10000001001100: color_data = 12'b010100000000;
		14'b10000001010000: color_data = 12'b010100000000;
		14'b10000001010001: color_data = 12'b010100000000;
		14'b10000001010010: color_data = 12'b010100000000;
		14'b10000001010011: color_data = 12'b010100000000;
		14'b10000001101000: color_data = 12'b010100000000;
		14'b10000001101001: color_data = 12'b101000000000;
		14'b10000001101010: color_data = 12'b101000000000;
		14'b10000001101011: color_data = 12'b101000000000;
		14'b10000001101100: color_data = 12'b010100000000;
		14'b10000010011101: color_data = 12'b010100000000;
		14'b10000010100000: color_data = 12'b010100000000;
		14'b10000010100001: color_data = 12'b101000000000;
		14'b10000010100010: color_data = 12'b101000000000;
		14'b10000010100011: color_data = 12'b101000000000;
		14'b10000010100100: color_data = 12'b101000000000;
		14'b10000010100101: color_data = 12'b010100000000;
		14'b10000010100110: color_data = 12'b010100000000;
		14'b10000010100111: color_data = 12'b010100000000;
		14'b10000010101000: color_data = 12'b101000000000;
		14'b10000010101001: color_data = 12'b101000000000;
		14'b10000010101010: color_data = 12'b010100000000;
		14'b10000010101011: color_data = 12'b010100000000;
		14'b10000010111000: color_data = 12'b010100000000;
		14'b10000010111001: color_data = 12'b010100000000;
		14'b10000010111011: color_data = 12'b010100000000;
		14'b10000010111100: color_data = 12'b010100000000;
		14'b10000010111101: color_data = 12'b010100000000;
		14'b10000010111110: color_data = 12'b101000000000;
		14'b10000010111111: color_data = 12'b101000000000;
		14'b10000011000000: color_data = 12'b101000000000;
		14'b10000011000001: color_data = 12'b101000000000;
		14'b10000011000010: color_data = 12'b101000000000;
		14'b10000011000011: color_data = 12'b101000000000;
		14'b10000011000100: color_data = 12'b101000000000;
		14'b10000011000101: color_data = 12'b101000000000;
		14'b10000011000110: color_data = 12'b101000000000;
		14'b10000011000111: color_data = 12'b101000000000;
		14'b10000011001000: color_data = 12'b101000000000;
		14'b10000011001001: color_data = 12'b101000000000;
		14'b10000011001010: color_data = 12'b101000000000;
		14'b10000011001011: color_data = 12'b101000000000;
		14'b10000011001100: color_data = 12'b101000000000;
		14'b10000011001101: color_data = 12'b010100000000;
		14'b10000011010000: color_data = 12'b010100000000;
		14'b10000011010001: color_data = 12'b010100000000;
		14'b10000011101000: color_data = 12'b010100000000;
		14'b10000011101001: color_data = 12'b101000000000;
		14'b10000011101010: color_data = 12'b101000000000;
		14'b10000011101011: color_data = 12'b101000000000;
		14'b10000011101100: color_data = 12'b010100000000;
		14'b10000100011111: color_data = 12'b010100000000;
		14'b10000100100000: color_data = 12'b101000000000;
		14'b10000100100001: color_data = 12'b101000000000;
		14'b10000100100010: color_data = 12'b101000000000;
		14'b10000100100011: color_data = 12'b101000000000;
		14'b10000100100100: color_data = 12'b101000000000;
		14'b10000100100101: color_data = 12'b010100000000;
		14'b10000100100110: color_data = 12'b010100000000;
		14'b10000100100111: color_data = 12'b010100000000;
		14'b10000100101000: color_data = 12'b101000000000;
		14'b10000100101001: color_data = 12'b010100000000;
		14'b10000100101010: color_data = 12'b010100000000;
		14'b10000100101011: color_data = 12'b010100000000;
		14'b10000100111100: color_data = 12'b010100000000;
		14'b10000100111101: color_data = 12'b101000000000;
		14'b10000100111110: color_data = 12'b101000000000;
		14'b10000100111111: color_data = 12'b101000000000;
		14'b10000101000000: color_data = 12'b101000000000;
		14'b10000101000001: color_data = 12'b010100000000;
		14'b10000101000010: color_data = 12'b010100000000;
		14'b10000101000011: color_data = 12'b101000000000;
		14'b10000101000100: color_data = 12'b101000000000;
		14'b10000101000101: color_data = 12'b101000000000;
		14'b10000101000110: color_data = 12'b101000000000;
		14'b10000101000111: color_data = 12'b101000000000;
		14'b10000101001000: color_data = 12'b101000000000;
		14'b10000101001001: color_data = 12'b101000000000;
		14'b10000101001010: color_data = 12'b101000000000;
		14'b10000101001011: color_data = 12'b101000000000;
		14'b10000101001100: color_data = 12'b101000000000;
		14'b10000101001101: color_data = 12'b101000000000;
		14'b10000101001110: color_data = 12'b010100000000;
		14'b10000101001111: color_data = 12'b010100000000;
		14'b10000101010001: color_data = 12'b010100000000;
		14'b10000101010010: color_data = 12'b010100000000;
		14'b10000101101001: color_data = 12'b010100000000;
		14'b10000101101010: color_data = 12'b101000000000;
		14'b10000101101011: color_data = 12'b101000000000;
		14'b10000101101100: color_data = 12'b101000000000;
		14'b10000101101101: color_data = 12'b010100000000;
		14'b10000110000000: color_data = 12'b010100000000;
		14'b10000110011110: color_data = 12'b010100000000;
		14'b10000110011111: color_data = 12'b101000000000;
		14'b10000110100000: color_data = 12'b101000000000;
		14'b10000110100001: color_data = 12'b101000000000;
		14'b10000110100010: color_data = 12'b101000000000;
		14'b10000110100011: color_data = 12'b101000000000;
		14'b10000110100100: color_data = 12'b101000000000;
		14'b10000110100101: color_data = 12'b010100000000;
		14'b10000110100110: color_data = 12'b010100000000;
		14'b10000110100111: color_data = 12'b010100000000;
		14'b10000110101000: color_data = 12'b101000000000;
		14'b10000110101001: color_data = 12'b010100000000;
		14'b10000110101010: color_data = 12'b010100000000;
		14'b10000110101011: color_data = 12'b010100000000;
		14'b10000110111011: color_data = 12'b010100000000;
		14'b10000110111100: color_data = 12'b010100000000;
		14'b10000110111101: color_data = 12'b101000000000;
		14'b10000110111110: color_data = 12'b101000000000;
		14'b10000110111111: color_data = 12'b010100000000;
		14'b10000111000000: color_data = 12'b010100000000;
		14'b10000111000001: color_data = 12'b010100000000;
		14'b10000111000010: color_data = 12'b010100000000;
		14'b10000111000011: color_data = 12'b101000000000;
		14'b10000111000100: color_data = 12'b101000000000;
		14'b10000111000101: color_data = 12'b101000000000;
		14'b10000111000110: color_data = 12'b101000000000;
		14'b10000111000111: color_data = 12'b101000000000;
		14'b10000111001000: color_data = 12'b010100000000;
		14'b10000111001001: color_data = 12'b010100000000;
		14'b10000111001010: color_data = 12'b101000000000;
		14'b10000111001011: color_data = 12'b101000000000;
		14'b10000111001100: color_data = 12'b101000000000;
		14'b10000111001101: color_data = 12'b101000000000;
		14'b10000111001110: color_data = 12'b101000000000;
		14'b10000111001111: color_data = 12'b010100000000;
		14'b10000111010000: color_data = 12'b010100000000;
		14'b10000111010001: color_data = 12'b010100000000;
		14'b10000111010010: color_data = 12'b010100000000;
		14'b10000111010011: color_data = 12'b010100000000;
		14'b10000111101001: color_data = 12'b010100000000;
		14'b10000111101010: color_data = 12'b010100000000;
		14'b10000111101011: color_data = 12'b101000000000;
		14'b10000111101100: color_data = 12'b101000000000;
		14'b10000111101101: color_data = 12'b010100000000;
		14'b10001000000000: color_data = 12'b010100000000;
		14'b10001000011110: color_data = 12'b010100000000;
		14'b10001000011111: color_data = 12'b101000000000;
		14'b10001000100000: color_data = 12'b101000000000;
		14'b10001000100001: color_data = 12'b101000000000;
		14'b10001000100010: color_data = 12'b101000000000;
		14'b10001000100011: color_data = 12'b101000000000;
		14'b10001000100100: color_data = 12'b101000000000;
		14'b10001000100101: color_data = 12'b101000000000;
		14'b10001000100110: color_data = 12'b010100000000;
		14'b10001000100111: color_data = 12'b010100000000;
		14'b10001000101000: color_data = 12'b010100000000;
		14'b10001000101001: color_data = 12'b010100000000;
		14'b10001000101010: color_data = 12'b101000000000;
		14'b10001000101011: color_data = 12'b010100000000;
		14'b10001000111011: color_data = 12'b010100000000;
		14'b10001000111100: color_data = 12'b010100000000;
		14'b10001000111101: color_data = 12'b010100000000;
		14'b10001000111110: color_data = 12'b010100000000;
		14'b10001001000000: color_data = 12'b010100000000;
		14'b10001001000001: color_data = 12'b010100000000;
		14'b10001001000010: color_data = 12'b101000000000;
		14'b10001001000011: color_data = 12'b101000000000;
		14'b10001001000100: color_data = 12'b101000000000;
		14'b10001001000101: color_data = 12'b101000000000;
		14'b10001001000110: color_data = 12'b010100000000;
		14'b10001001001010: color_data = 12'b101000000000;
		14'b10001001001011: color_data = 12'b010100000000;
		14'b10001001001100: color_data = 12'b010100000000;
		14'b10001001001101: color_data = 12'b101000000000;
		14'b10001001001110: color_data = 12'b101000000000;
		14'b10001001001111: color_data = 12'b101000000000;
		14'b10001001010000: color_data = 12'b010100000000;
		14'b10001001010001: color_data = 12'b010100000000;
		14'b10001001010010: color_data = 12'b101000000000;
		14'b10001001010011: color_data = 12'b010100000000;
		14'b10001001101010: color_data = 12'b010100000000;
		14'b10001001101011: color_data = 12'b101000000000;
		14'b10001001101100: color_data = 12'b101000000000;
		14'b10001001101101: color_data = 12'b010100000000;
		14'b10001010000000: color_data = 12'b010100000000;
		14'b10001010011110: color_data = 12'b101000000000;
		14'b10001010011111: color_data = 12'b101000000000;
		14'b10001010100000: color_data = 12'b101000000000;
		14'b10001010100001: color_data = 12'b101000000000;
		14'b10001010100010: color_data = 12'b101000000000;
		14'b10001010100011: color_data = 12'b101000000000;
		14'b10001010100100: color_data = 12'b101000000000;
		14'b10001010100101: color_data = 12'b101000000000;
		14'b10001010100110: color_data = 12'b010100000000;
		14'b10001010100111: color_data = 12'b010100000000;
		14'b10001010101000: color_data = 12'b010100000000;
		14'b10001010101001: color_data = 12'b010100000000;
		14'b10001010101010: color_data = 12'b101000000000;
		14'b10001010101011: color_data = 12'b010100000000;
		14'b10001011000000: color_data = 12'b010100000000;
		14'b10001011000001: color_data = 12'b101000000000;
		14'b10001011000010: color_data = 12'b101000000000;
		14'b10001011000011: color_data = 12'b101000000000;
		14'b10001011000100: color_data = 12'b010100000000;
		14'b10001011000101: color_data = 12'b010100000000;
		14'b10001011001001: color_data = 12'b010100000000;
		14'b10001011001010: color_data = 12'b101000000000;
		14'b10001011001011: color_data = 12'b010100000000;
		14'b10001011001100: color_data = 12'b010100000000;
		14'b10001011001101: color_data = 12'b010100000000;
		14'b10001011001110: color_data = 12'b101000000000;
		14'b10001011001111: color_data = 12'b101000000000;
		14'b10001011010000: color_data = 12'b101000000000;
		14'b10001011010001: color_data = 12'b010100000000;
		14'b10001011010010: color_data = 12'b010100000000;
		14'b10001011010011: color_data = 12'b101000000000;
		14'b10001011010100: color_data = 12'b010100000000;
		14'b10001011101010: color_data = 12'b010100000000;
		14'b10001011101011: color_data = 12'b101000000000;
		14'b10001011101100: color_data = 12'b101000000000;
		14'b10001011101101: color_data = 12'b101000000000;
		14'b10001100000000: color_data = 12'b010100000000;
		14'b10001100011010: color_data = 12'b010100000000;
		14'b10001100011101: color_data = 12'b010100000000;
		14'b10001100011110: color_data = 12'b101000000000;
		14'b10001100011111: color_data = 12'b101000000000;
		14'b10001100100000: color_data = 12'b101000000000;
		14'b10001100100001: color_data = 12'b101000000000;
		14'b10001100100010: color_data = 12'b101000000000;
		14'b10001100100011: color_data = 12'b101000000000;
		14'b10001100100100: color_data = 12'b101000000000;
		14'b10001100100101: color_data = 12'b010100000000;
		14'b10001100100110: color_data = 12'b010100000000;
		14'b10001100100111: color_data = 12'b010100000000;
		14'b10001100101000: color_data = 12'b010100000000;
		14'b10001100101001: color_data = 12'b101000000000;
		14'b10001100101010: color_data = 12'b101000000000;
		14'b10001100101011: color_data = 12'b010100000000;
		14'b10001100111110: color_data = 12'b010100000000;
		14'b10001100111111: color_data = 12'b010100000000;
		14'b10001101000000: color_data = 12'b101000000000;
		14'b10001101000001: color_data = 12'b101000000000;
		14'b10001101000010: color_data = 12'b101000000000;
		14'b10001101000011: color_data = 12'b101000000000;
		14'b10001101000100: color_data = 12'b010100000000;
		14'b10001101001000: color_data = 12'b010100000000;
		14'b10001101001001: color_data = 12'b101000000000;
		14'b10001101001010: color_data = 12'b101000000000;
		14'b10001101001011: color_data = 12'b010100000000;
		14'b10001101001101: color_data = 12'b010100000000;
		14'b10001101001110: color_data = 12'b101000000000;
		14'b10001101001111: color_data = 12'b101000000000;
		14'b10001101010000: color_data = 12'b101000000000;
		14'b10001101010001: color_data = 12'b101000000000;
		14'b10001101010010: color_data = 12'b010100000000;
		14'b10001101010011: color_data = 12'b010100000000;
		14'b10001101010100: color_data = 12'b010100000000;
		14'b10001101101010: color_data = 12'b010100000000;
		14'b10001101101011: color_data = 12'b101000000000;
		14'b10001101101100: color_data = 12'b101000000000;
		14'b10001101101101: color_data = 12'b101000000000;
		14'b10001110000000: color_data = 12'b010100000000;
		14'b10001110010101: color_data = 12'b010100000000;
		14'b10001110011010: color_data = 12'b010100000000;
		14'b10001110011101: color_data = 12'b010100000000;
		14'b10001110011110: color_data = 12'b101000000000;
		14'b10001110011111: color_data = 12'b101000000000;
		14'b10001110100000: color_data = 12'b101000000000;
		14'b10001110100001: color_data = 12'b101000000000;
		14'b10001110100010: color_data = 12'b101000000000;
		14'b10001110100011: color_data = 12'b010100000000;
		14'b10001110100100: color_data = 12'b010100000000;
		14'b10001110100101: color_data = 12'b010100000000;
		14'b10001110100110: color_data = 12'b010100000000;
		14'b10001110100111: color_data = 12'b101000000000;
		14'b10001110101000: color_data = 12'b101000000000;
		14'b10001110101001: color_data = 12'b101000000000;
		14'b10001110101010: color_data = 12'b101000000000;
		14'b10001110101011: color_data = 12'b010100000000;
		14'b10001110111101: color_data = 12'b010100000000;
		14'b10001110111110: color_data = 12'b010100000000;
		14'b10001110111111: color_data = 12'b101000000000;
		14'b10001111000000: color_data = 12'b101000000000;
		14'b10001111000001: color_data = 12'b101000000000;
		14'b10001111000010: color_data = 12'b101000000000;
		14'b10001111000011: color_data = 12'b010100000000;
		14'b10001111000100: color_data = 12'b010100000000;
		14'b10001111000101: color_data = 12'b010100000000;
		14'b10001111000110: color_data = 12'b010100000000;
		14'b10001111000111: color_data = 12'b101000000000;
		14'b10001111001000: color_data = 12'b101000000000;
		14'b10001111001001: color_data = 12'b101000000000;
		14'b10001111001010: color_data = 12'b101000000000;
		14'b10001111001011: color_data = 12'b101000000000;
		14'b10001111001100: color_data = 12'b010100000000;
		14'b10001111001101: color_data = 12'b010100000000;
		14'b10001111001110: color_data = 12'b101000000000;
		14'b10001111001111: color_data = 12'b101000000000;
		14'b10001111010000: color_data = 12'b101000000000;
		14'b10001111010001: color_data = 12'b101000000000;
		14'b10001111010010: color_data = 12'b010100000000;
		14'b10001111010011: color_data = 12'b010100000000;
		14'b10001111010100: color_data = 12'b010100000000;
		14'b10001111101010: color_data = 12'b010100000000;
		14'b10001111101011: color_data = 12'b101000000000;
		14'b10001111101100: color_data = 12'b101000000000;
		14'b10001111101101: color_data = 12'b101000000000;
		14'b10010000000000: color_data = 12'b010100000000;
		14'b10010000010101: color_data = 12'b010100000000;
		14'b10010000010110: color_data = 12'b010100000000;
		14'b10010000011101: color_data = 12'b010100000000;
		14'b10010000011110: color_data = 12'b101000000000;
		14'b10010000011111: color_data = 12'b101000000000;
		14'b10010000100000: color_data = 12'b101000000000;
		14'b10010000100001: color_data = 12'b101000000000;
		14'b10010000100010: color_data = 12'b010100000000;
		14'b10010000100011: color_data = 12'b010100000000;
		14'b10010000100100: color_data = 12'b010100000000;
		14'b10010000100101: color_data = 12'b010100000000;
		14'b10010000100110: color_data = 12'b101000000000;
		14'b10010000100111: color_data = 12'b101000000000;
		14'b10010000101000: color_data = 12'b101000000000;
		14'b10010000101001: color_data = 12'b101000000000;
		14'b10010000101010: color_data = 12'b101000000000;
		14'b10010000101011: color_data = 12'b010100000000;
		14'b10010000111100: color_data = 12'b010100000000;
		14'b10010000111101: color_data = 12'b101000000000;
		14'b10010000111110: color_data = 12'b101000000000;
		14'b10010000111111: color_data = 12'b101000000000;
		14'b10010001000000: color_data = 12'b101000000000;
		14'b10010001000001: color_data = 12'b101000000000;
		14'b10010001000010: color_data = 12'b101000000000;
		14'b10010001000011: color_data = 12'b101000000000;
		14'b10010001000100: color_data = 12'b101000000000;
		14'b10010001000101: color_data = 12'b101000000000;
		14'b10010001000110: color_data = 12'b010100000000;
		14'b10010001000111: color_data = 12'b010100000000;
		14'b10010001001000: color_data = 12'b010100000000;
		14'b10010001001001: color_data = 12'b101000000000;
		14'b10010001001010: color_data = 12'b101000000000;
		14'b10010001001011: color_data = 12'b101000000000;
		14'b10010001001100: color_data = 12'b101000000000;
		14'b10010001001101: color_data = 12'b101000000000;
		14'b10010001001110: color_data = 12'b101000000000;
		14'b10010001001111: color_data = 12'b101000000000;
		14'b10010001010000: color_data = 12'b101000000000;
		14'b10010001010001: color_data = 12'b101000000000;
		14'b10010001010010: color_data = 12'b101000000000;
		14'b10010001010011: color_data = 12'b010100000000;
		14'b10010001101010: color_data = 12'b010100000000;
		14'b10010001101011: color_data = 12'b101000000000;
		14'b10010001101100: color_data = 12'b101000000000;
		14'b10010001101101: color_data = 12'b101000000000;
		14'b10010010000000: color_data = 12'b010100000000;
		14'b10010010001100: color_data = 12'b010100000000;
		14'b10010010001101: color_data = 12'b010100000000;
		14'b10010010001110: color_data = 12'b010100000000;
		14'b10010010001111: color_data = 12'b010100000000;
		14'b10010010010001: color_data = 12'b010100000000;
		14'b10010010010010: color_data = 12'b010100000000;
		14'b10010010010011: color_data = 12'b010100000000;
		14'b10010010010100: color_data = 12'b010100000000;
		14'b10010010010101: color_data = 12'b010100000000;
		14'b10010010010110: color_data = 12'b010100000000;
		14'b10010010011101: color_data = 12'b010100000000;
		14'b10010010011110: color_data = 12'b101000000000;
		14'b10010010011111: color_data = 12'b101000000000;
		14'b10010010100000: color_data = 12'b101000000000;
		14'b10010010100001: color_data = 12'b010100000000;
		14'b10010010100010: color_data = 12'b010100000000;
		14'b10010010100011: color_data = 12'b010100000000;
		14'b10010010100100: color_data = 12'b010100000000;
		14'b10010010100101: color_data = 12'b101000000000;
		14'b10010010100110: color_data = 12'b101000000000;
		14'b10010010100111: color_data = 12'b101000000000;
		14'b10010010101000: color_data = 12'b101000000000;
		14'b10010010101001: color_data = 12'b101000000000;
		14'b10010010101010: color_data = 12'b101000000000;
		14'b10010010101011: color_data = 12'b010100000000;
		14'b10010010111010: color_data = 12'b010100000000;
		14'b10010010111011: color_data = 12'b010100000000;
		14'b10010010111100: color_data = 12'b101000000000;
		14'b10010010111101: color_data = 12'b101000000000;
		14'b10010010111110: color_data = 12'b101000000000;
		14'b10010010111111: color_data = 12'b101000000000;
		14'b10010011000000: color_data = 12'b101000000000;
		14'b10010011000001: color_data = 12'b101000000000;
		14'b10010011000010: color_data = 12'b101000000000;
		14'b10010011000011: color_data = 12'b101000000000;
		14'b10010011000100: color_data = 12'b101000000000;
		14'b10010011000101: color_data = 12'b010100000000;
		14'b10010011001000: color_data = 12'b010100000000;
		14'b10010011001001: color_data = 12'b101000000000;
		14'b10010011001010: color_data = 12'b101000000000;
		14'b10010011001011: color_data = 12'b101000000000;
		14'b10010011001100: color_data = 12'b101000000000;
		14'b10010011001101: color_data = 12'b101000000000;
		14'b10010011001110: color_data = 12'b101000000000;
		14'b10010011001111: color_data = 12'b101000000000;
		14'b10010011010000: color_data = 12'b101000000000;
		14'b10010011010001: color_data = 12'b101000000000;
		14'b10010011010010: color_data = 12'b101000000000;
		14'b10010011010011: color_data = 12'b010100000000;
		14'b10010011101010: color_data = 12'b010100000000;
		14'b10010011101011: color_data = 12'b101000000000;
		14'b10010011101100: color_data = 12'b101000000000;
		14'b10010011101101: color_data = 12'b101000000000;
		14'b10010100000000: color_data = 12'b010100000000;
		14'b10010100000001: color_data = 12'b010100000000;
		14'b10010100001101: color_data = 12'b010100000000;
		14'b10010100001110: color_data = 12'b010100000000;
		14'b10010100001111: color_data = 12'b010100000000;
		14'b10010100010000: color_data = 12'b010100000000;
		14'b10010100010001: color_data = 12'b101000000000;
		14'b10010100010010: color_data = 12'b101000000000;
		14'b10010100010011: color_data = 12'b101000000000;
		14'b10010100010100: color_data = 12'b101000000000;
		14'b10010100010101: color_data = 12'b010100000000;
		14'b10010100010110: color_data = 12'b010100000000;
		14'b10010100011101: color_data = 12'b010100000000;
		14'b10010100011110: color_data = 12'b101000000000;
		14'b10010100011111: color_data = 12'b101000000000;
		14'b10010100100000: color_data = 12'b010100000000;
		14'b10010100100001: color_data = 12'b010100000000;
		14'b10010100100010: color_data = 12'b010100000000;
		14'b10010100100011: color_data = 12'b101000000000;
		14'b10010100100100: color_data = 12'b101000000000;
		14'b10010100100101: color_data = 12'b101000000000;
		14'b10010100100110: color_data = 12'b101000000000;
		14'b10010100100111: color_data = 12'b101000000000;
		14'b10010100101000: color_data = 12'b101000000000;
		14'b10010100101001: color_data = 12'b101000000000;
		14'b10010100101010: color_data = 12'b010100000000;
		14'b10010100101011: color_data = 12'b010100000000;
		14'b10010100111010: color_data = 12'b010100000000;
		14'b10010100111011: color_data = 12'b101000000000;
		14'b10010100111100: color_data = 12'b101000000000;
		14'b10010100111101: color_data = 12'b101000000000;
		14'b10010100111110: color_data = 12'b101000000000;
		14'b10010100111111: color_data = 12'b101000000000;
		14'b10010101000000: color_data = 12'b101000000000;
		14'b10010101000001: color_data = 12'b010100000000;
		14'b10010101000010: color_data = 12'b010100000000;
		14'b10010101000011: color_data = 12'b010100000000;
		14'b10010101000100: color_data = 12'b010100000000;
		14'b10010101001000: color_data = 12'b010100000000;
		14'b10010101001001: color_data = 12'b101000000000;
		14'b10010101001010: color_data = 12'b101000000000;
		14'b10010101001011: color_data = 12'b101000000000;
		14'b10010101001100: color_data = 12'b101000000000;
		14'b10010101001101: color_data = 12'b101000000000;
		14'b10010101001110: color_data = 12'b101000000000;
		14'b10010101001111: color_data = 12'b101000000000;
		14'b10010101010000: color_data = 12'b010100000000;
		14'b10010101010001: color_data = 12'b010100000000;
		14'b10010101010010: color_data = 12'b101000000000;
		14'b10010101010011: color_data = 12'b010100000000;
		14'b10010101101010: color_data = 12'b010100000000;
		14'b10010101101011: color_data = 12'b101000000000;
		14'b10010101101100: color_data = 12'b101000000000;
		14'b10010101101101: color_data = 12'b101000000000;
		14'b10010110000000: color_data = 12'b010100000000;
		14'b10010110000001: color_data = 12'b010100000000;
		14'b10010110001101: color_data = 12'b010100000000;
		14'b10010110001110: color_data = 12'b101000000000;
		14'b10010110001111: color_data = 12'b101000000000;
		14'b10010110010000: color_data = 12'b101000000000;
		14'b10010110010001: color_data = 12'b101000000000;
		14'b10010110010010: color_data = 12'b101000000000;
		14'b10010110010011: color_data = 12'b101000000000;
		14'b10010110010100: color_data = 12'b101000000000;
		14'b10010110010101: color_data = 12'b101000000000;
		14'b10010110010110: color_data = 12'b010100000000;
		14'b10010110010111: color_data = 12'b010100000000;
		14'b10010110011101: color_data = 12'b010100000000;
		14'b10010110011110: color_data = 12'b101000000000;
		14'b10010110011111: color_data = 12'b101000000000;
		14'b10010110100000: color_data = 12'b010100000000;
		14'b10010110100001: color_data = 12'b010100000000;
		14'b10010110100010: color_data = 12'b101000000000;
		14'b10010110100011: color_data = 12'b101000000000;
		14'b10010110100100: color_data = 12'b101000000000;
		14'b10010110100101: color_data = 12'b101000000000;
		14'b10010110100110: color_data = 12'b101000000000;
		14'b10010110100111: color_data = 12'b101000000000;
		14'b10010110101000: color_data = 12'b010100000000;
		14'b10010110101001: color_data = 12'b010100000000;
		14'b10010110101010: color_data = 12'b010100000000;
		14'b10010110111001: color_data = 12'b010100000000;
		14'b10010110111010: color_data = 12'b101000000000;
		14'b10010110111011: color_data = 12'b101000000000;
		14'b10010110111100: color_data = 12'b101000000000;
		14'b10010110111101: color_data = 12'b101000000000;
		14'b10010110111110: color_data = 12'b101000000000;
		14'b10010110111111: color_data = 12'b010100000000;
		14'b10010111000000: color_data = 12'b010100000000;
		14'b10010111001000: color_data = 12'b010100000000;
		14'b10010111001001: color_data = 12'b010100000000;
		14'b10010111001010: color_data = 12'b101000000000;
		14'b10010111001011: color_data = 12'b101000000000;
		14'b10010111001100: color_data = 12'b101000000000;
		14'b10010111001101: color_data = 12'b101000000000;
		14'b10010111001110: color_data = 12'b101000000000;
		14'b10010111001111: color_data = 12'b101000000000;
		14'b10010111010000: color_data = 12'b101000000000;
		14'b10010111010001: color_data = 12'b010100000000;
		14'b10010111010010: color_data = 12'b010100000000;
		14'b10010111010011: color_data = 12'b010100000000;
		14'b10010111101011: color_data = 12'b101000000000;
		14'b10010111101100: color_data = 12'b101000000000;
		14'b10010111101101: color_data = 12'b101000000000;
		14'b10011000000000: color_data = 12'b010100000000;
		14'b10011000000001: color_data = 12'b010100000000;
		14'b10011000001100: color_data = 12'b010100000000;
		14'b10011000001101: color_data = 12'b101000000000;
		14'b10011000001110: color_data = 12'b101000000000;
		14'b10011000001111: color_data = 12'b101000000000;
		14'b10011000010000: color_data = 12'b101000000000;
		14'b10011000010001: color_data = 12'b101000000000;
		14'b10011000010010: color_data = 12'b101000000000;
		14'b10011000010011: color_data = 12'b101000000000;
		14'b10011000010100: color_data = 12'b101000000000;
		14'b10011000010101: color_data = 12'b101000000000;
		14'b10011000010110: color_data = 12'b101000000000;
		14'b10011000010111: color_data = 12'b010100000000;
		14'b10011000011101: color_data = 12'b010100000000;
		14'b10011000011110: color_data = 12'b101000000000;
		14'b10011000011111: color_data = 12'b101000000000;
		14'b10011000100000: color_data = 12'b101000000000;
		14'b10011000100001: color_data = 12'b101000000000;
		14'b10011000100010: color_data = 12'b101000000000;
		14'b10011000100011: color_data = 12'b101000000000;
		14'b10011000100100: color_data = 12'b101000000000;
		14'b10011000100101: color_data = 12'b101000000000;
		14'b10011000100110: color_data = 12'b010100000000;
		14'b10011000100111: color_data = 12'b010100000000;
		14'b10011000101000: color_data = 12'b010100000000;
		14'b10011000111000: color_data = 12'b010100000000;
		14'b10011000111001: color_data = 12'b101000000000;
		14'b10011000111010: color_data = 12'b101000000000;
		14'b10011000111011: color_data = 12'b101000000000;
		14'b10011000111100: color_data = 12'b010100000000;
		14'b10011000111101: color_data = 12'b010100000000;
		14'b10011001001000: color_data = 12'b010100000000;
		14'b10011001001001: color_data = 12'b010100000000;
		14'b10011001001010: color_data = 12'b101000000000;
		14'b10011001001011: color_data = 12'b101000000000;
		14'b10011001001100: color_data = 12'b101000000000;
		14'b10011001001101: color_data = 12'b101000000000;
		14'b10011001001110: color_data = 12'b101000000000;
		14'b10011001001111: color_data = 12'b101000000000;
		14'b10011001010000: color_data = 12'b010100000000;
		14'b10011001010010: color_data = 12'b010100000000;
		14'b10011001010011: color_data = 12'b010100000000;
		14'b10011001101011: color_data = 12'b101000000000;
		14'b10011001101100: color_data = 12'b101000000000;
		14'b10011001101101: color_data = 12'b101000000000;
		14'b10011010000000: color_data = 12'b010100000000;
		14'b10011010000001: color_data = 12'b010100000000;
		14'b10011010001011: color_data = 12'b010100000000;
		14'b10011010001100: color_data = 12'b101000000000;
		14'b10011010001101: color_data = 12'b101000000000;
		14'b10011010001110: color_data = 12'b101000000000;
		14'b10011010001111: color_data = 12'b101000000000;
		14'b10011010010000: color_data = 12'b010100000000;
		14'b10011010010001: color_data = 12'b010100000000;
		14'b10011010010010: color_data = 12'b101000000000;
		14'b10011010010011: color_data = 12'b101000000000;
		14'b10011010010100: color_data = 12'b010100000000;
		14'b10011010010101: color_data = 12'b010100000000;
		14'b10011010010110: color_data = 12'b101000000000;
		14'b10011010010111: color_data = 12'b101000000000;
		14'b10011010011000: color_data = 12'b010100000000;
		14'b10011010011011: color_data = 12'b010100000000;
		14'b10011010011101: color_data = 12'b010100000000;
		14'b10011010011110: color_data = 12'b101000000000;
		14'b10011010011111: color_data = 12'b101000000000;
		14'b10011010100000: color_data = 12'b101000000000;
		14'b10011010100001: color_data = 12'b101000000000;
		14'b10011010100010: color_data = 12'b101000000000;
		14'b10011010100011: color_data = 12'b101000000000;
		14'b10011010100100: color_data = 12'b101000000000;
		14'b10011010100101: color_data = 12'b010100000000;
		14'b10011010110111: color_data = 12'b010100000000;
		14'b10011010111000: color_data = 12'b010100000000;
		14'b10011010111001: color_data = 12'b101000000000;
		14'b10011010111010: color_data = 12'b010100000000;
		14'b10011010111011: color_data = 12'b010100000000;
		14'b10011011000011: color_data = 12'b010100000000;
		14'b10011011000100: color_data = 12'b010100000000;
		14'b10011011001000: color_data = 12'b010100000000;
		14'b10011011001001: color_data = 12'b010100000000;
		14'b10011011001010: color_data = 12'b010100000000;
		14'b10011011001011: color_data = 12'b010100000000;
		14'b10011011001100: color_data = 12'b010100000000;
		14'b10011011001101: color_data = 12'b010100000000;
		14'b10011011001110: color_data = 12'b010100000000;
		14'b10011011001111: color_data = 12'b010100000000;
		14'b10011011010000: color_data = 12'b010100000000;
		14'b10011011010011: color_data = 12'b010100000000;
		14'b10011011101011: color_data = 12'b101000000000;
		14'b10011011101100: color_data = 12'b101000000000;
		14'b10011011101101: color_data = 12'b101000000000;
		14'b10011100000000: color_data = 12'b010100000000;
		14'b10011100000001: color_data = 12'b010100000000;
		14'b10011100001011: color_data = 12'b010100000000;
		14'b10011100001100: color_data = 12'b010100000000;
		14'b10011100001101: color_data = 12'b010100000000;
		14'b10011100001110: color_data = 12'b101000000000;
		14'b10011100001111: color_data = 12'b010100000000;
		14'b10011100010010: color_data = 12'b010100000000;
		14'b10011100010011: color_data = 12'b101000000000;
		14'b10011100010100: color_data = 12'b010100000000;
		14'b10011100010110: color_data = 12'b010100000000;
		14'b10011100010111: color_data = 12'b101000000000;
		14'b10011100011000: color_data = 12'b010100000000;
		14'b10011100011011: color_data = 12'b010100000000;
		14'b10011100011101: color_data = 12'b010100000000;
		14'b10011100011110: color_data = 12'b101000000000;
		14'b10011100011111: color_data = 12'b101000000000;
		14'b10011100100000: color_data = 12'b101000000000;
		14'b10011100100001: color_data = 12'b101000000000;
		14'b10011100100010: color_data = 12'b101000000000;
		14'b10011100100011: color_data = 12'b101000000000;
		14'b10011100100100: color_data = 12'b010100000000;
		14'b10011100110101: color_data = 12'b010100000000;
		14'b10011100110110: color_data = 12'b010100000000;
		14'b10011100110111: color_data = 12'b010100000000;
		14'b10011100111000: color_data = 12'b101000000000;
		14'b10011100111001: color_data = 12'b101000000000;
		14'b10011100111010: color_data = 12'b010100000000;
		14'b10011101000101: color_data = 12'b010100000000;
		14'b10011101000110: color_data = 12'b010100000000;
		14'b10011101001001: color_data = 12'b010100000000;
		14'b10011101001010: color_data = 12'b010100000000;
		14'b10011101001011: color_data = 12'b010100000000;
		14'b10011101001100: color_data = 12'b010100000000;
		14'b10011101001101: color_data = 12'b010100000000;
		14'b10011101001110: color_data = 12'b010100000000;
		14'b10011101001111: color_data = 12'b101000000000;
		14'b10011101010000: color_data = 12'b010100000000;
		14'b10011101010011: color_data = 12'b010100000000;
		14'b10011101101011: color_data = 12'b101000000000;
		14'b10011101101100: color_data = 12'b101000000000;
		14'b10011101101101: color_data = 12'b101000000000;
		14'b10011110000000: color_data = 12'b010100000000;
		14'b10011110000001: color_data = 12'b010100000000;
		14'b10011110001100: color_data = 12'b010100000000;
		14'b10011110001101: color_data = 12'b101000000000;
		14'b10011110001110: color_data = 12'b010100000000;
		14'b10011110010010: color_data = 12'b010100000000;
		14'b10011110010011: color_data = 12'b101000000000;
		14'b10011110010100: color_data = 12'b010100000000;
		14'b10011110010111: color_data = 12'b010100000000;
		14'b10011110011000: color_data = 12'b101000000000;
		14'b10011110011100: color_data = 12'b010100000000;
		14'b10011110011101: color_data = 12'b010100000000;
		14'b10011110011110: color_data = 12'b101000000000;
		14'b10011110011111: color_data = 12'b101000000000;
		14'b10011110100000: color_data = 12'b101000000000;
		14'b10011110100001: color_data = 12'b101000000000;
		14'b10011110100010: color_data = 12'b101000000000;
		14'b10011110100011: color_data = 12'b101000000000;
		14'b10011110100100: color_data = 12'b010100000000;
		14'b10011110110101: color_data = 12'b010100000000;
		14'b10011110110110: color_data = 12'b010100000000;
		14'b10011110110111: color_data = 12'b101000000000;
		14'b10011110111000: color_data = 12'b101000000000;
		14'b10011110111001: color_data = 12'b010100000000;
		14'b10011111000101: color_data = 12'b010100000000;
		14'b10011111000110: color_data = 12'b010100000000;
		14'b10011111001001: color_data = 12'b010100000000;
		14'b10011111001010: color_data = 12'b010100000000;
		14'b10011111001110: color_data = 12'b010100000000;
		14'b10011111001111: color_data = 12'b101000000000;
		14'b10011111010000: color_data = 12'b010100000000;
		14'b10011111010011: color_data = 12'b010100000000;
		14'b10011111101011: color_data = 12'b101000000000;
		14'b10011111101100: color_data = 12'b101000000000;
		14'b10011111101101: color_data = 12'b101000000000;
		14'b10100000000000: color_data = 12'b010100000000;
		14'b10100000000001: color_data = 12'b010100000000;
		14'b10100000001100: color_data = 12'b010100000000;
		14'b10100000001101: color_data = 12'b010100000000;
		14'b10100000010000: color_data = 12'b010100000000;
		14'b10100000010001: color_data = 12'b010100000000;
		14'b10100000010010: color_data = 12'b101000000000;
		14'b10100000010011: color_data = 12'b101000000000;
		14'b10100000010100: color_data = 12'b101000000000;
		14'b10100000010101: color_data = 12'b010100000000;
		14'b10100000010111: color_data = 12'b010100000000;
		14'b10100000011000: color_data = 12'b010100000000;
		14'b10100000011001: color_data = 12'b010100000000;
		14'b10100000011100: color_data = 12'b010100000000;
		14'b10100000011101: color_data = 12'b010100000000;
		14'b10100000011110: color_data = 12'b101000000000;
		14'b10100000011111: color_data = 12'b101000000000;
		14'b10100000100000: color_data = 12'b101000000000;
		14'b10100000100001: color_data = 12'b101000000000;
		14'b10100000100010: color_data = 12'b101000000000;
		14'b10100000100011: color_data = 12'b101000000000;
		14'b10100000100100: color_data = 12'b010100000000;
		14'b10100000110101: color_data = 12'b010100000000;
		14'b10100000110110: color_data = 12'b101000000000;
		14'b10100000110111: color_data = 12'b101000000000;
		14'b10100000111000: color_data = 12'b010100000000;
		14'b10100001000111: color_data = 12'b010100000000;
		14'b10100001001101: color_data = 12'b010100000000;
		14'b10100001001110: color_data = 12'b101000000000;
		14'b10100001001111: color_data = 12'b101000000000;
		14'b10100001010000: color_data = 12'b010100000000;
		14'b10100001010011: color_data = 12'b010100000000;
		14'b10100001101011: color_data = 12'b101000000000;
		14'b10100001101100: color_data = 12'b101000000000;
		14'b10100001101101: color_data = 12'b101000000000;
		14'b10100010000000: color_data = 12'b010100000000;
		14'b10100010000001: color_data = 12'b010100000000;
		14'b10100010001011: color_data = 12'b010100000000;
		14'b10100010001100: color_data = 12'b010100000000;
		14'b10100010001101: color_data = 12'b010100000000;
		14'b10100010001110: color_data = 12'b010100000000;
		14'b10100010001111: color_data = 12'b101000000000;
		14'b10100010010000: color_data = 12'b101000000000;
		14'b10100010010001: color_data = 12'b101000000000;
		14'b10100010010010: color_data = 12'b101000000000;
		14'b10100010010011: color_data = 12'b101000000000;
		14'b10100010010100: color_data = 12'b101000000000;
		14'b10100010010101: color_data = 12'b101000000000;
		14'b10100010010110: color_data = 12'b010100000000;
		14'b10100010011000: color_data = 12'b010100000000;
		14'b10100010011001: color_data = 12'b010100000000;
		14'b10100010011100: color_data = 12'b010100000000;
		14'b10100010011101: color_data = 12'b010100000000;
		14'b10100010011110: color_data = 12'b101000000000;
		14'b10100010011111: color_data = 12'b101000000000;
		14'b10100010100000: color_data = 12'b101000000000;
		14'b10100010100001: color_data = 12'b101000000000;
		14'b10100010100010: color_data = 12'b101000000000;
		14'b10100010100011: color_data = 12'b101000000000;
		14'b10100010100100: color_data = 12'b010100000000;
		14'b10100010110100: color_data = 12'b010100000000;
		14'b10100010110101: color_data = 12'b010100000000;
		14'b10100010110110: color_data = 12'b101000000000;
		14'b10100010110111: color_data = 12'b010100000000;
		14'b10100010111000: color_data = 12'b010100000000;
		14'b10100011000110: color_data = 12'b010100000000;
		14'b10100011000111: color_data = 12'b101000000000;
		14'b10100011001100: color_data = 12'b010100000000;
		14'b10100011001101: color_data = 12'b101000000000;
		14'b10100011001110: color_data = 12'b101000000000;
		14'b10100011001111: color_data = 12'b101000000000;
		14'b10100011010000: color_data = 12'b010100000000;
		14'b10100011101010: color_data = 12'b010100000000;
		14'b10100011101011: color_data = 12'b101000000000;
		14'b10100011101100: color_data = 12'b101000000000;
		14'b10100011101101: color_data = 12'b101000000000;
		14'b10100100000000: color_data = 12'b010100000000;
		14'b10100100000001: color_data = 12'b010100000000;
		14'b10100100001100: color_data = 12'b010100000000;
		14'b10100100001101: color_data = 12'b101000000000;
		14'b10100100001110: color_data = 12'b101000000000;
		14'b10100100001111: color_data = 12'b010100000000;
		14'b10100100010000: color_data = 12'b101000000000;
		14'b10100100010001: color_data = 12'b101000000000;
		14'b10100100010010: color_data = 12'b101000000000;
		14'b10100100010011: color_data = 12'b101000000000;
		14'b10100100010100: color_data = 12'b101000000000;
		14'b10100100010101: color_data = 12'b101000000000;
		14'b10100100010110: color_data = 12'b101000000000;
		14'b10100100010111: color_data = 12'b010100000000;
		14'b10100100011000: color_data = 12'b010100000000;
		14'b10100100011001: color_data = 12'b010100000000;
		14'b10100100011101: color_data = 12'b010100000000;
		14'b10100100011110: color_data = 12'b101000000000;
		14'b10100100011111: color_data = 12'b101000000000;
		14'b10100100100000: color_data = 12'b101000000000;
		14'b10100100100001: color_data = 12'b101000000000;
		14'b10100100100010: color_data = 12'b101000000000;
		14'b10100100100011: color_data = 12'b101000000000;
		14'b10100100100100: color_data = 12'b101000000000;
		14'b10100100110100: color_data = 12'b010100000000;
		14'b10100100110101: color_data = 12'b101000000000;
		14'b10100100110110: color_data = 12'b010100000000;
		14'b10100100110111: color_data = 12'b010100000000;
		14'b10100100111000: color_data = 12'b010100000000;
		14'b10100101000111: color_data = 12'b010100000000;
		14'b10100101001100: color_data = 12'b010100000000;
		14'b10100101001101: color_data = 12'b101000000000;
		14'b10100101001110: color_data = 12'b101000000000;
		14'b10100101001111: color_data = 12'b101000000000;
		14'b10100101101010: color_data = 12'b010100000000;
		14'b10100101101011: color_data = 12'b101000000000;
		14'b10100101101100: color_data = 12'b101000000000;
		14'b10100101101101: color_data = 12'b101000000000;
		14'b10100110000000: color_data = 12'b010100000000;
		14'b10100110001100: color_data = 12'b010100000000;
		14'b10100110001101: color_data = 12'b010100000000;
		14'b10100110001110: color_data = 12'b010100000000;
		14'b10100110001111: color_data = 12'b010100000000;
		14'b10100110010000: color_data = 12'b101000000000;
		14'b10100110010001: color_data = 12'b101000000000;
		14'b10100110010010: color_data = 12'b101000000000;
		14'b10100110010011: color_data = 12'b010100000000;
		14'b10100110010100: color_data = 12'b010100000000;
		14'b10100110010101: color_data = 12'b101000000000;
		14'b10100110010110: color_data = 12'b101000000000;
		14'b10100110010111: color_data = 12'b010100000000;
		14'b10100110011000: color_data = 12'b010100000000;
		14'b10100110011001: color_data = 12'b010100000000;
		14'b10100110011101: color_data = 12'b010100000000;
		14'b10100110011110: color_data = 12'b101000000000;
		14'b10100110011111: color_data = 12'b101000000000;
		14'b10100110100000: color_data = 12'b101000000000;
		14'b10100110100001: color_data = 12'b101000000000;
		14'b10100110100010: color_data = 12'b101000000000;
		14'b10100110100011: color_data = 12'b101000000000;
		14'b10100110100100: color_data = 12'b101000000000;
		14'b10100110100101: color_data = 12'b010100000000;
		14'b10100110110011: color_data = 12'b010100000000;
		14'b10100110110100: color_data = 12'b010100000000;
		14'b10100110110101: color_data = 12'b010100000000;
		14'b10100110110110: color_data = 12'b010100000000;
		14'b10100110110111: color_data = 12'b010100000000;
		14'b10100111001011: color_data = 12'b010100000000;
		14'b10100111001100: color_data = 12'b101000000000;
		14'b10100111001101: color_data = 12'b101000000000;
		14'b10100111001110: color_data = 12'b101000000000;
		14'b10100111001111: color_data = 12'b010100000000;
		14'b10100111101010: color_data = 12'b010100000000;
		14'b10100111101011: color_data = 12'b101000000000;
		14'b10100111101100: color_data = 12'b101000000000;
		14'b10100111101101: color_data = 12'b101000000000;
		14'b10101000000000: color_data = 12'b010100000000;
		14'b10101000001110: color_data = 12'b010100000000;
		14'b10101000001111: color_data = 12'b101000000000;
		14'b10101000010000: color_data = 12'b101000000000;
		14'b10101000010001: color_data = 12'b010100000000;
		14'b10101000010100: color_data = 12'b010100000000;
		14'b10101000010101: color_data = 12'b010100000000;
		14'b10101000010110: color_data = 12'b101000000000;
		14'b10101000010111: color_data = 12'b101000000000;
		14'b10101000011000: color_data = 12'b010100000000;
		14'b10101000011001: color_data = 12'b010100000000;
		14'b10101000011110: color_data = 12'b010100000000;
		14'b10101000011111: color_data = 12'b101000000000;
		14'b10101000100000: color_data = 12'b101000000000;
		14'b10101000100001: color_data = 12'b101000000000;
		14'b10101000100010: color_data = 12'b101000000000;
		14'b10101000100011: color_data = 12'b101000000000;
		14'b10101000100100: color_data = 12'b010100000000;
		14'b10101000100101: color_data = 12'b010100000000;
		14'b10101000110011: color_data = 12'b010100000000;
		14'b10101000110100: color_data = 12'b010100000000;
		14'b10101000110101: color_data = 12'b010100000000;
		14'b10101000111000: color_data = 12'b010100000000;
		14'b10101001001010: color_data = 12'b010100000000;
		14'b10101001001011: color_data = 12'b101000000000;
		14'b10101001001100: color_data = 12'b101000000000;
		14'b10101001001101: color_data = 12'b101000000000;
		14'b10101001001110: color_data = 12'b101000000000;
		14'b10101001001111: color_data = 12'b010100000000;
		14'b10101001101010: color_data = 12'b010100000000;
		14'b10101001101011: color_data = 12'b101000000000;
		14'b10101001101100: color_data = 12'b101000000000;
		14'b10101001101101: color_data = 12'b101000000000;
		14'b10101010000000: color_data = 12'b010100000000;
		14'b10101010001101: color_data = 12'b010100000000;
		14'b10101010001110: color_data = 12'b101000000000;
		14'b10101010001111: color_data = 12'b101000000000;
		14'b10101010010000: color_data = 12'b010100000000;
		14'b10101010010001: color_data = 12'b010100000000;
		14'b10101010010010: color_data = 12'b010100000000;
		14'b10101010010011: color_data = 12'b010100000000;
		14'b10101010010100: color_data = 12'b101000000000;
		14'b10101010010101: color_data = 12'b010100000000;
		14'b10101010010110: color_data = 12'b010100000000;
		14'b10101010010111: color_data = 12'b101000000000;
		14'b10101010011000: color_data = 12'b010100000000;
		14'b10101010011001: color_data = 12'b010100000000;
		14'b10101010011110: color_data = 12'b010100000000;
		14'b10101010011111: color_data = 12'b101000000000;
		14'b10101010100000: color_data = 12'b101000000000;
		14'b10101010100001: color_data = 12'b101000000000;
		14'b10101010100010: color_data = 12'b101000000000;
		14'b10101010100011: color_data = 12'b101000000000;
		14'b10101010100100: color_data = 12'b010100000000;
		14'b10101010110011: color_data = 12'b010100000000;
		14'b10101010110100: color_data = 12'b010100000000;
		14'b10101010110101: color_data = 12'b010100000000;
		14'b10101010111000: color_data = 12'b010100000000;
		14'b10101011001001: color_data = 12'b010100000000;
		14'b10101011001010: color_data = 12'b101000000000;
		14'b10101011001011: color_data = 12'b101000000000;
		14'b10101011001100: color_data = 12'b101000000000;
		14'b10101011001101: color_data = 12'b101000000000;
		14'b10101011001110: color_data = 12'b010100000000;
		14'b10101011101010: color_data = 12'b010100000000;
		14'b10101011101011: color_data = 12'b101000000000;
		14'b10101011101100: color_data = 12'b101000000000;
		14'b10101011101101: color_data = 12'b101000000000;
		14'b10101100000000: color_data = 12'b010100000000;
		14'b10101100001100: color_data = 12'b010100000000;
		14'b10101100001101: color_data = 12'b101000000000;
		14'b10101100001110: color_data = 12'b101000000000;
		14'b10101100001111: color_data = 12'b101000000000;
		14'b10101100010000: color_data = 12'b101000000000;
		14'b10101100010001: color_data = 12'b010100000000;
		14'b10101100010010: color_data = 12'b010100000000;
		14'b10101100010011: color_data = 12'b101000000000;
		14'b10101100010100: color_data = 12'b101000000000;
		14'b10101100010101: color_data = 12'b101000000000;
		14'b10101100010110: color_data = 12'b101000000000;
		14'b10101100010111: color_data = 12'b101000000000;
		14'b10101100011000: color_data = 12'b101000000000;
		14'b10101100011001: color_data = 12'b010100000000;
		14'b10101100011110: color_data = 12'b010100000000;
		14'b10101100011111: color_data = 12'b101000000000;
		14'b10101100100000: color_data = 12'b101000000000;
		14'b10101100100001: color_data = 12'b101000000000;
		14'b10101100100010: color_data = 12'b101000000000;
		14'b10101100100011: color_data = 12'b010100000000;
		14'b10101100110011: color_data = 12'b010100000000;
		14'b10101100110100: color_data = 12'b010100000000;
		14'b10101100110101: color_data = 12'b010100000000;
		14'b10101100111000: color_data = 12'b010100000000;
		14'b10101100111001: color_data = 12'b010100000000;
		14'b10101101000111: color_data = 12'b010100000000;
		14'b10101101001000: color_data = 12'b010100000000;
		14'b10101101001001: color_data = 12'b101000000000;
		14'b10101101001010: color_data = 12'b101000000000;
		14'b10101101001011: color_data = 12'b101000000000;
		14'b10101101001100: color_data = 12'b101000000000;
		14'b10101101001101: color_data = 12'b010100000000;
		14'b10101101101001: color_data = 12'b010100000000;
		14'b10101101101010: color_data = 12'b101000000000;
		14'b10101101101011: color_data = 12'b101000000000;
		14'b10101101101100: color_data = 12'b101000000000;
		14'b10101101101101: color_data = 12'b010100000000;
		14'b10101110001011: color_data = 12'b010100000000;
		14'b10101110001100: color_data = 12'b101000000000;
		14'b10101110001101: color_data = 12'b101000000000;
		14'b10101110001110: color_data = 12'b101000000000;
		14'b10101110001111: color_data = 12'b101000000000;
		14'b10101110010000: color_data = 12'b010100000000;
		14'b10101110010001: color_data = 12'b010100000000;
		14'b10101110010011: color_data = 12'b010100000000;
		14'b10101110010100: color_data = 12'b101000000000;
		14'b10101110010101: color_data = 12'b101000000000;
		14'b10101110010110: color_data = 12'b101000000000;
		14'b10101110010111: color_data = 12'b101000000000;
		14'b10101110011000: color_data = 12'b101000000000;
		14'b10101110011001: color_data = 12'b010100000000;
		14'b10101110011111: color_data = 12'b010100000000;
		14'b10101110100000: color_data = 12'b101000000000;
		14'b10101110100001: color_data = 12'b101000000000;
		14'b10101110100010: color_data = 12'b101000000000;
		14'b10101110100011: color_data = 12'b010100000000;
		14'b10101110110011: color_data = 12'b010100000000;
		14'b10101110110100: color_data = 12'b010100000000;
		14'b10101110111010: color_data = 12'b010100000000;
		14'b10101111000110: color_data = 12'b010100000000;
		14'b10101111000111: color_data = 12'b010100000000;
		14'b10101111001000: color_data = 12'b101000000000;
		14'b10101111001001: color_data = 12'b101000000000;
		14'b10101111001010: color_data = 12'b101000000000;
		14'b10101111001011: color_data = 12'b101000000000;
		14'b10101111001100: color_data = 12'b010100000000;
		14'b10101111001101: color_data = 12'b010100000000;
		14'b10101111101001: color_data = 12'b010100000000;
		14'b10101111101010: color_data = 12'b101000000000;
		14'b10101111101011: color_data = 12'b101000000000;
		14'b10101111101100: color_data = 12'b101000000000;
		14'b10101111101101: color_data = 12'b010100000000;
		14'b10110000001010: color_data = 12'b010100000000;
		14'b10110000001011: color_data = 12'b101000000000;
		14'b10110000001100: color_data = 12'b101000000000;
		14'b10110000001101: color_data = 12'b101000000000;
		14'b10110000001110: color_data = 12'b010100000000;
		14'b10110000001111: color_data = 12'b010100000000;
		14'b10110000010011: color_data = 12'b010100000000;
		14'b10110000010100: color_data = 12'b101000000000;
		14'b10110000010101: color_data = 12'b101000000000;
		14'b10110000010110: color_data = 12'b101000000000;
		14'b10110000010111: color_data = 12'b010100000000;
		14'b10110000011000: color_data = 12'b010100000000;
		14'b10110000011111: color_data = 12'b010100000000;
		14'b10110000100000: color_data = 12'b101000000000;
		14'b10110000100001: color_data = 12'b101000000000;
		14'b10110000100010: color_data = 12'b101000000000;
		14'b10110000110011: color_data = 12'b010100000000;
		14'b10110001000101: color_data = 12'b010100000000;
		14'b10110001000110: color_data = 12'b010100000000;
		14'b10110001000111: color_data = 12'b101000000000;
		14'b10110001001000: color_data = 12'b101000000000;
		14'b10110001001001: color_data = 12'b101000000000;
		14'b10110001001010: color_data = 12'b101000000000;
		14'b10110001001011: color_data = 12'b010100000000;
		14'b10110001001100: color_data = 12'b010100000000;
		14'b10110001101000: color_data = 12'b010100000000;
		14'b10110001101001: color_data = 12'b101000000000;
		14'b10110001101010: color_data = 12'b101000000000;
		14'b10110001101011: color_data = 12'b101000000000;
		14'b10110001101100: color_data = 12'b101000000000;
		14'b10110001101101: color_data = 12'b010100000000;
		14'b10110010001001: color_data = 12'b010100000000;
		14'b10110010001010: color_data = 12'b101000000000;
		14'b10110010001011: color_data = 12'b101000000000;
		14'b10110010001100: color_data = 12'b010100000000;
		14'b10110010010011: color_data = 12'b010100000000;
		14'b10110010010100: color_data = 12'b101000000000;
		14'b10110010010101: color_data = 12'b101000000000;
		14'b10110010010110: color_data = 12'b101000000000;
		14'b10110010010111: color_data = 12'b010100000000;
		14'b10110010011000: color_data = 12'b010100000000;
		14'b10110010011111: color_data = 12'b010100000000;
		14'b10110010100000: color_data = 12'b101000000000;
		14'b10110010100001: color_data = 12'b101000000000;
		14'b10110010100010: color_data = 12'b101000000000;
		14'b10110010110011: color_data = 12'b010100000000;
		14'b10110011000100: color_data = 12'b010100000000;
		14'b10110011000101: color_data = 12'b010100000000;
		14'b10110011000110: color_data = 12'b101000000000;
		14'b10110011000111: color_data = 12'b101000000000;
		14'b10110011001000: color_data = 12'b101000000000;
		14'b10110011001001: color_data = 12'b101000000000;
		14'b10110011001010: color_data = 12'b010100000000;
		14'b10110011101000: color_data = 12'b010100000000;
		14'b10110011101001: color_data = 12'b101000000000;
		14'b10110011101010: color_data = 12'b101000000000;
		14'b10110011101011: color_data = 12'b101000000000;
		14'b10110011101100: color_data = 12'b010100000000;
		14'b10110011101101: color_data = 12'b010100000000;
		14'b10110100001000: color_data = 12'b010100000000;
		14'b10110100001001: color_data = 12'b010100000000;
		14'b10110100001010: color_data = 12'b010100000000;
		14'b10110100010011: color_data = 12'b010100000000;
		14'b10110100010100: color_data = 12'b010100000000;
		14'b10110100010101: color_data = 12'b010100000000;
		14'b10110100010110: color_data = 12'b010100000000;
		14'b10110100010111: color_data = 12'b010100000000;
		14'b10110100100000: color_data = 12'b101000000000;
		14'b10110100100001: color_data = 12'b101000000000;
		14'b10110100100010: color_data = 12'b010100000000;
		14'b10110100100011: color_data = 12'b010100000000;
		14'b10110100110011: color_data = 12'b010100000000;
		14'b10110101000011: color_data = 12'b010100000000;
		14'b10110101000100: color_data = 12'b010100000000;
		14'b10110101000101: color_data = 12'b101000000000;
		14'b10110101000110: color_data = 12'b101000000000;
		14'b10110101000111: color_data = 12'b101000000000;
		14'b10110101001000: color_data = 12'b101000000000;
		14'b10110101001001: color_data = 12'b010100000000;
		14'b10110101100111: color_data = 12'b010100000000;
		14'b10110101101000: color_data = 12'b101000000000;
		14'b10110101101001: color_data = 12'b101000000000;
		14'b10110101101010: color_data = 12'b101000000000;
		14'b10110101101011: color_data = 12'b010100000000;
		14'b10110101101100: color_data = 12'b010100000000;
		14'b10110110001000: color_data = 12'b010100000000;
		14'b10110110001001: color_data = 12'b101000000000;
		14'b10110110001010: color_data = 12'b010100000000;
		14'b10110110010011: color_data = 12'b010100000000;
		14'b10110110010101: color_data = 12'b010100000000;
		14'b10110110010110: color_data = 12'b010100000000;
		14'b10110110100000: color_data = 12'b101000000000;
		14'b10110110100001: color_data = 12'b101000000000;
		14'b10110110100010: color_data = 12'b010100000000;
		14'b10110110100011: color_data = 12'b010100000000;
		14'b10110110110011: color_data = 12'b010100000000;
		14'b10110111000011: color_data = 12'b010100000000;
		14'b10110111000100: color_data = 12'b010100000000;
		14'b10110111000101: color_data = 12'b101000000000;
		14'b10110111000110: color_data = 12'b010100000000;
		14'b10110111000111: color_data = 12'b010100000000;
		14'b10110111001000: color_data = 12'b010100000000;
		14'b10110111100110: color_data = 12'b010100000000;
		14'b10110111100111: color_data = 12'b010100000000;
		14'b10110111101000: color_data = 12'b101000000000;
		14'b10110111101001: color_data = 12'b010100000000;
		14'b10110111101010: color_data = 12'b010100000000;
		14'b10110111101011: color_data = 12'b010100000000;
		14'b10111000000111: color_data = 12'b010100000000;
		14'b10111000001000: color_data = 12'b101000000000;
		14'b10111000001001: color_data = 12'b010100000000;
		14'b10111000010001: color_data = 12'b010100000000;
		14'b10111000010101: color_data = 12'b010100000000;
		14'b10111000010110: color_data = 12'b010100000000;
		14'b10111000100000: color_data = 12'b010100000000;
		14'b10111000100001: color_data = 12'b101000000000;
		14'b10111000100010: color_data = 12'b010100000000;
		14'b10111000100011: color_data = 12'b010100000000;
		14'b10111000110011: color_data = 12'b010100000000;
		14'b10111001000010: color_data = 12'b010100000000;
		14'b10111001000011: color_data = 12'b010100000000;
		14'b10111001000100: color_data = 12'b010100000000;
		14'b10111001000101: color_data = 12'b010100000000;
		14'b10111001000110: color_data = 12'b010100000000;
		14'b10111001000111: color_data = 12'b010100000000;
		14'b10111001100110: color_data = 12'b010100000000;
		14'b10111001100111: color_data = 12'b101000000000;
		14'b10111001101000: color_data = 12'b101000000000;
		14'b10111001101001: color_data = 12'b010100000000;
		14'b10111001101010: color_data = 12'b010100000000;
		14'b10111001101011: color_data = 12'b010100000000;
		14'b10111010000111: color_data = 12'b010100000000;
		14'b10111010001000: color_data = 12'b010100000000;
		14'b10111010010001: color_data = 12'b010100000000;
		14'b10111010010100: color_data = 12'b010100000000;
		14'b10111010010101: color_data = 12'b101000000000;
		14'b10111010010110: color_data = 12'b010100000000;
		14'b10111010100000: color_data = 12'b010100000000;
		14'b10111010100001: color_data = 12'b101000000000;
		14'b10111010100010: color_data = 12'b101000000000;
		14'b10111010100011: color_data = 12'b010100000000;
		14'b10111011000001: color_data = 12'b010100000000;
		14'b10111011000010: color_data = 12'b010100000000;
		14'b10111011000011: color_data = 12'b010100000000;
		14'b10111011000100: color_data = 12'b010100000000;
		14'b10111011000101: color_data = 12'b010100000000;
		14'b10111011000110: color_data = 12'b010100000000;
		14'b10111011100110: color_data = 12'b010100000000;
		14'b10111011100111: color_data = 12'b101000000000;
		14'b10111011101000: color_data = 12'b010100000000;
		14'b10111011101001: color_data = 12'b010100000000;
		14'b10111011101010: color_data = 12'b101000000000;
		14'b10111011101011: color_data = 12'b010100000000;
		14'b10111100000110: color_data = 12'b010100000000;
		14'b10111100000111: color_data = 12'b010100000000;
		14'b10111100001000: color_data = 12'b010100000000;
		14'b10111100010011: color_data = 12'b010100000000;
		14'b10111100010100: color_data = 12'b101000000000;
		14'b10111100010101: color_data = 12'b101000000000;
		14'b10111100100000: color_data = 12'b010100000000;
		14'b10111100100001: color_data = 12'b101000000000;
		14'b10111100100010: color_data = 12'b101000000000;
		14'b10111100100011: color_data = 12'b010100000000;
		14'b10111101000001: color_data = 12'b010100000000;
		14'b10111101000010: color_data = 12'b010100000000;
		14'b10111101000011: color_data = 12'b010100000000;
		14'b10111101000100: color_data = 12'b010100000000;
		14'b10111101100110: color_data = 12'b010100000000;
		14'b10111101100111: color_data = 12'b010100000000;
		14'b10111101101000: color_data = 12'b010100000000;
		14'b10111101101001: color_data = 12'b010100000000;
		14'b10111101101010: color_data = 12'b010100000000;
		14'b10111101101011: color_data = 12'b010100000000;
		14'b10111110000110: color_data = 12'b010100000000;
		14'b10111110010010: color_data = 12'b010100000000;
		14'b10111110010011: color_data = 12'b101000000000;
		14'b10111110010100: color_data = 12'b101000000000;
		14'b10111110010101: color_data = 12'b010100000000;
		14'b10111110100000: color_data = 12'b010100000000;
		14'b10111110100001: color_data = 12'b101000000000;
		14'b10111110100010: color_data = 12'b101000000000;
		14'b10111110100011: color_data = 12'b010100000000;
		14'b10111111000000: color_data = 12'b010100000000;
		14'b10111111000001: color_data = 12'b010100000000;
		14'b10111111000010: color_data = 12'b010100000000;
		14'b10111111100101: color_data = 12'b010100000000;
		14'b10111111100110: color_data = 12'b010100000000;
		14'b10111111100111: color_data = 12'b010100000000;
		14'b10111111101000: color_data = 12'b010100000000;
		14'b10111111101001: color_data = 12'b010100000000;
		14'b11000000000110: color_data = 12'b010100000000;
		14'b11000000001001: color_data = 12'b010100000000;
		14'b11000000010001: color_data = 12'b010100000000;
		14'b11000000010010: color_data = 12'b101000000000;
		14'b11000000010011: color_data = 12'b101000000000;
		14'b11000000010100: color_data = 12'b010100000000;
		14'b11000000100000: color_data = 12'b010100000000;
		14'b11000000100001: color_data = 12'b101000000000;
		14'b11000000100010: color_data = 12'b101000000000;
		14'b11000000100011: color_data = 12'b010100000000;
		14'b11000000100100: color_data = 12'b010100000000;
		14'b11000001000000: color_data = 12'b010100000000;
		14'b11000001100100: color_data = 12'b010100000000;
		14'b11000001100101: color_data = 12'b010100000000;
		14'b11000001100110: color_data = 12'b010100000000;
		14'b11000001100111: color_data = 12'b010100000000;
		14'b11000010000110: color_data = 12'b010100000000;
		14'b11000010010000: color_data = 12'b010100000000;
		14'b11000010010001: color_data = 12'b101000000000;
		14'b11000010010010: color_data = 12'b101000000000;
		14'b11000010010011: color_data = 12'b010100000000;
		14'b11000010100000: color_data = 12'b010100000000;
		14'b11000010100001: color_data = 12'b101000000000;
		14'b11000010100010: color_data = 12'b101000000000;
		14'b11000010100011: color_data = 12'b101000000000;
		14'b11000010100100: color_data = 12'b010100000000;
		14'b11000010100101: color_data = 12'b010100000000;
		14'b11000010100110: color_data = 12'b010100000000;
		14'b11000011000000: color_data = 12'b010100000000;
		14'b11000011100011: color_data = 12'b010100000000;
		14'b11000011100100: color_data = 12'b010100000000;
		14'b11000011100101: color_data = 12'b010100000000;
		14'b11000011100110: color_data = 12'b010100000000;
		14'b11000100001111: color_data = 12'b010100000000;
		14'b11000100010000: color_data = 12'b101000000000;
		14'b11000100010001: color_data = 12'b101000000000;
		14'b11000100010010: color_data = 12'b010100000000;
		14'b11000100100000: color_data = 12'b101000000000;
		14'b11000100100001: color_data = 12'b101000000000;
		14'b11000100100010: color_data = 12'b101000000000;
		14'b11000100100011: color_data = 12'b101000000000;
		14'b11000100100100: color_data = 12'b101000000000;
		14'b11000100100101: color_data = 12'b010100000000;
		14'b11000100100110: color_data = 12'b010100000000;
		14'b11000100100111: color_data = 12'b010100000000;
		14'b11000101000000: color_data = 12'b010100000000;
		14'b11000101100010: color_data = 12'b010100000000;
		14'b11000101100011: color_data = 12'b101000000000;
		14'b11000101100100: color_data = 12'b010100000000;
		14'b11000110001111: color_data = 12'b010100000000;
		14'b11000110010000: color_data = 12'b101000000000;
		14'b11000110010001: color_data = 12'b010100000000;
		14'b11000110011111: color_data = 12'b010100000000;
		14'b11000110100000: color_data = 12'b101000000000;
		14'b11000110100001: color_data = 12'b101000000000;
		14'b11000110100010: color_data = 12'b010100000000;
		14'b11000110100011: color_data = 12'b101000000000;
		14'b11000110100100: color_data = 12'b101000000000;
		14'b11000110100101: color_data = 12'b010100000000;
		14'b11000110100110: color_data = 12'b010100000000;
		14'b11000110100111: color_data = 12'b010100000000;
		14'b11000110101000: color_data = 12'b010100000000;
		14'b11000111100001: color_data = 12'b010100000000;
		14'b11000111100010: color_data = 12'b010100000000;
		14'b11000111100011: color_data = 12'b101000000000;
		14'b11000111100100: color_data = 12'b010100000000;
		14'b11001000001110: color_data = 12'b010100000000;
		14'b11001000001111: color_data = 12'b010100000000;
		14'b11001000010000: color_data = 12'b010100000000;
		14'b11001000011110: color_data = 12'b010100000000;
		14'b11001000011111: color_data = 12'b101000000000;
		14'b11001000100000: color_data = 12'b101000000000;
		14'b11001000100001: color_data = 12'b101000000000;
		14'b11001000100010: color_data = 12'b010100000000;
		14'b11001000100011: color_data = 12'b101000000000;
		14'b11001000100100: color_data = 12'b101000000000;
		14'b11001000100101: color_data = 12'b101000000000;
		14'b11001000100110: color_data = 12'b010100000000;
		14'b11001000100111: color_data = 12'b010100000000;
		14'b11001000101000: color_data = 12'b010100000000;
		14'b11001000101001: color_data = 12'b010100000000;
		14'b11001001100000: color_data = 12'b010100000000;
		14'b11001001100001: color_data = 12'b010100000000;
		14'b11001001100010: color_data = 12'b101000000000;
		14'b11001001100011: color_data = 12'b010100000000;
		14'b11001010001101: color_data = 12'b010100000000;
		14'b11001010001110: color_data = 12'b010100000000;
		14'b11001010001111: color_data = 12'b010100000000;
		14'b11001010011100: color_data = 12'b010100000000;
		14'b11001010011101: color_data = 12'b010100000000;
		14'b11001010011110: color_data = 12'b101000000000;
		14'b11001010011111: color_data = 12'b101000000000;
		14'b11001010100000: color_data = 12'b101000000000;
		14'b11001010100001: color_data = 12'b101000000000;
		14'b11001010100010: color_data = 12'b010100000000;
		14'b11001010100011: color_data = 12'b101000000000;
		14'b11001010100100: color_data = 12'b101000000000;
		14'b11001010100101: color_data = 12'b101000000000;
		14'b11001010100110: color_data = 12'b101000000000;
		14'b11001010100111: color_data = 12'b101000000000;
		14'b11001010101000: color_data = 12'b010100000000;
		14'b11001010101001: color_data = 12'b010100000000;
		14'b11001011011110: color_data = 12'b010100000000;
		14'b11001011011111: color_data = 12'b010100000000;
		14'b11001011100000: color_data = 12'b010100000000;
		14'b11001011100001: color_data = 12'b101000000000;
		14'b11001011100010: color_data = 12'b101000000000;
		14'b11001011100011: color_data = 12'b010100000000;
		14'b11001100001101: color_data = 12'b010100000000;
		14'b11001100011001: color_data = 12'b010100000000;
		14'b11001100011010: color_data = 12'b010100000000;
		14'b11001100011011: color_data = 12'b010100000000;
		14'b11001100011100: color_data = 12'b101000000000;
		14'b11001100011101: color_data = 12'b101000000000;
		14'b11001100011110: color_data = 12'b101000000000;
		14'b11001100011111: color_data = 12'b101000000000;
		14'b11001100100000: color_data = 12'b101000000000;
		14'b11001100100001: color_data = 12'b010100000000;
		14'b11001100100010: color_data = 12'b101000000000;
		14'b11001100100011: color_data = 12'b101000000000;
		14'b11001100100100: color_data = 12'b101000000000;
		14'b11001100100101: color_data = 12'b101000000000;
		14'b11001100100110: color_data = 12'b101000000000;
		14'b11001100100111: color_data = 12'b101000000000;
		14'b11001100101000: color_data = 12'b010100000000;
		14'b11001100101001: color_data = 12'b010100000000;
		14'b11001101011100: color_data = 12'b010100000000;
		14'b11001101011101: color_data = 12'b010100000000;
		14'b11001101011110: color_data = 12'b010100000000;
		14'b11001101011111: color_data = 12'b010100000000;
		14'b11001101100000: color_data = 12'b101000000000;
		14'b11001101100001: color_data = 12'b101000000000;
		14'b11001101100010: color_data = 12'b010100000000;
		14'b11001110010110: color_data = 12'b010100000000;
		14'b11001110010111: color_data = 12'b010100000000;
		14'b11001110011000: color_data = 12'b010100000000;
		14'b11001110011001: color_data = 12'b101000000000;
		14'b11001110011010: color_data = 12'b101000000000;
		14'b11001110011011: color_data = 12'b101000000000;
		14'b11001110011100: color_data = 12'b101000000000;
		14'b11001110011101: color_data = 12'b101000000000;
		14'b11001110011110: color_data = 12'b101000000000;
		14'b11001110011111: color_data = 12'b101000000000;
		14'b11001110100000: color_data = 12'b010100000000;
		14'b11001110100001: color_data = 12'b010100000000;
		14'b11001110100010: color_data = 12'b101000000000;
		14'b11001110100011: color_data = 12'b101000000000;
		14'b11001110100100: color_data = 12'b101000000000;
		14'b11001110100101: color_data = 12'b101000000000;
		14'b11001110100110: color_data = 12'b101000000000;
		14'b11001110100111: color_data = 12'b101000000000;
		14'b11001110101000: color_data = 12'b010100000000;
		14'b11001110101001: color_data = 12'b010100000000;
		14'b11001111011010: color_data = 12'b010100000000;
		14'b11001111011011: color_data = 12'b010100000000;
		14'b11001111011100: color_data = 12'b010100000000;
		14'b11001111011101: color_data = 12'b010100000000;
		14'b11001111011110: color_data = 12'b010100000000;
		14'b11001111011111: color_data = 12'b101000000000;
		14'b11001111100000: color_data = 12'b101000000000;
		14'b11001111100001: color_data = 12'b101000000000;
		14'b11001111100010: color_data = 12'b010100000000;
		14'b11010000010011: color_data = 12'b010100000000;
		14'b11010000010100: color_data = 12'b010100000000;
		14'b11010000010101: color_data = 12'b101000000000;
		14'b11010000010110: color_data = 12'b101000000000;
		14'b11010000010111: color_data = 12'b101000000000;
		14'b11010000011000: color_data = 12'b101000000000;
		14'b11010000011001: color_data = 12'b101000000000;
		14'b11010000011010: color_data = 12'b101000000000;
		14'b11010000011011: color_data = 12'b101000000000;
		14'b11010000011100: color_data = 12'b101000000000;
		14'b11010000011101: color_data = 12'b101000000000;
		14'b11010000011110: color_data = 12'b101000000000;
		14'b11010000011111: color_data = 12'b101000000000;
		14'b11010000100000: color_data = 12'b101000000000;
		14'b11010000100001: color_data = 12'b101000000000;
		14'b11010000100010: color_data = 12'b101000000000;
		14'b11010000100011: color_data = 12'b101000000000;
		14'b11010000100100: color_data = 12'b101000000000;
		14'b11010000100101: color_data = 12'b101000000000;
		14'b11010000100110: color_data = 12'b010100000000;
		14'b11010000100111: color_data = 12'b010100000000;
		14'b11010000101000: color_data = 12'b010100000000;
		14'b11010000101001: color_data = 12'b010100000000;
		14'b11010001010111: color_data = 12'b010100000000;
		14'b11010001011000: color_data = 12'b010100000000;
		14'b11010001011001: color_data = 12'b010100000000;
		14'b11010001011010: color_data = 12'b010100000000;
		14'b11010001011011: color_data = 12'b010100000000;
		14'b11010001011100: color_data = 12'b010100000000;
		14'b11010001011101: color_data = 12'b010100000000;
		14'b11010001011110: color_data = 12'b101000000000;
		14'b11010001011111: color_data = 12'b101000000000;
		14'b11010001100000: color_data = 12'b101000000000;
		14'b11010001100001: color_data = 12'b101000000000;
		14'b11010001100010: color_data = 12'b010100000000;
		14'b11010010001111: color_data = 12'b010100000000;
		14'b11010010010000: color_data = 12'b010100000000;
		14'b11010010010001: color_data = 12'b010100000000;
		14'b11010010010010: color_data = 12'b010100000000;
		14'b11010010010011: color_data = 12'b010100000000;
		14'b11010010010100: color_data = 12'b010100000000;
		14'b11010010010101: color_data = 12'b010100000000;
		14'b11010010010110: color_data = 12'b010100000000;
		14'b11010010010111: color_data = 12'b101000000000;
		14'b11010010011000: color_data = 12'b101000000000;
		14'b11010010011001: color_data = 12'b101000000000;
		14'b11010010011010: color_data = 12'b101000000000;
		14'b11010010011011: color_data = 12'b101000000000;
		14'b11010010011100: color_data = 12'b101000000000;
		14'b11010010011101: color_data = 12'b101000000000;
		14'b11010010011110: color_data = 12'b101000000000;
		14'b11010010011111: color_data = 12'b101000000000;
		14'b11010010100000: color_data = 12'b101000000000;
		14'b11010010100001: color_data = 12'b101000000000;
		14'b11010010100010: color_data = 12'b101000000000;
		14'b11010010100011: color_data = 12'b010100000000;
		14'b11010010100100: color_data = 12'b010100000000;
		14'b11010010100101: color_data = 12'b010100000000;
		14'b11010010100110: color_data = 12'b010100000000;
		14'b11010010100111: color_data = 12'b010100000000;
		14'b11010010101000: color_data = 12'b010100000000;
		14'b11010011010011: color_data = 12'b010100000000;
		14'b11010011010100: color_data = 12'b010100000000;
		14'b11010011010101: color_data = 12'b010100000000;
		14'b11010011010110: color_data = 12'b010100000000;
		14'b11010011010111: color_data = 12'b010100000000;
		14'b11010011011000: color_data = 12'b010100000000;
		14'b11010011011001: color_data = 12'b010100000000;
		14'b11010011011010: color_data = 12'b010100000000;
		14'b11010011011011: color_data = 12'b010100000000;
		14'b11010011011100: color_data = 12'b010100000000;
		14'b11010011011101: color_data = 12'b101000000000;
		14'b11010011011110: color_data = 12'b101000000000;
		14'b11010011011111: color_data = 12'b101000000000;
		14'b11010011100000: color_data = 12'b101000000000;
		14'b11010011100001: color_data = 12'b010100000000;
		14'b11010011100010: color_data = 12'b010100000000;
		14'b11010100001000: color_data = 12'b010100000000;
		14'b11010100001111: color_data = 12'b010100000000;
		14'b11010100010000: color_data = 12'b010100000000;
		14'b11010100010001: color_data = 12'b010100000000;
		14'b11010100010010: color_data = 12'b010100000000;
		14'b11010100010011: color_data = 12'b010100000000;
		14'b11010100010100: color_data = 12'b010100000000;
		14'b11010100010101: color_data = 12'b010100000000;
		14'b11010100010110: color_data = 12'b101000000000;
		14'b11010100010111: color_data = 12'b101000000000;
		14'b11010100011000: color_data = 12'b101000000000;
		14'b11010100011001: color_data = 12'b101000000000;
		14'b11010100011010: color_data = 12'b101000000000;
		14'b11010100011011: color_data = 12'b101000000000;
		14'b11010100011100: color_data = 12'b010100000000;
		14'b11010100011101: color_data = 12'b010100000000;
		14'b11010100011110: color_data = 12'b010100000000;
		14'b11010100011111: color_data = 12'b010100000000;
		14'b11010100100000: color_data = 12'b010100000000;
		14'b11010100100001: color_data = 12'b010100000000;
		14'b11010100100010: color_data = 12'b010100000000;
		14'b11010100100011: color_data = 12'b010100000000;
		14'b11010100100100: color_data = 12'b010100000000;
		14'b11010100100101: color_data = 12'b010100000000;
		14'b11010101000100: color_data = 12'b010100000000;
		14'b11010101010000: color_data = 12'b010100000000;
		14'b11010101010001: color_data = 12'b010100000000;
		14'b11010101010010: color_data = 12'b010100000000;
		14'b11010101010011: color_data = 12'b010100000000;
		14'b11010101010100: color_data = 12'b010100000000;
		14'b11010101010101: color_data = 12'b010100000000;
		14'b11010101010110: color_data = 12'b010100000000;
		14'b11010101010111: color_data = 12'b010100000000;
		14'b11010101011000: color_data = 12'b010100000000;
		14'b11010101011001: color_data = 12'b010100000000;
		14'b11010101011010: color_data = 12'b010100000000;
		14'b11010101011011: color_data = 12'b010100000000;
		14'b11010101011100: color_data = 12'b101000000000;
		14'b11010101011101: color_data = 12'b101000000000;
		14'b11010101011110: color_data = 12'b101000000000;
		14'b11010101011111: color_data = 12'b010100000000;
		14'b11010101100000: color_data = 12'b010100000000;
		14'b11010110001011: color_data = 12'b010100000000;
		14'b11010110001100: color_data = 12'b010100000000;
		14'b11010110001101: color_data = 12'b010100000000;
		14'b11010110001110: color_data = 12'b010100000000;
		14'b11010110001111: color_data = 12'b010100000000;
		14'b11010110010000: color_data = 12'b010100000000;
		14'b11010110010001: color_data = 12'b010100000000;
		14'b11010110010010: color_data = 12'b010100000000;
		14'b11010110010011: color_data = 12'b010100000000;
		14'b11010110010100: color_data = 12'b010100000000;
		14'b11010110010101: color_data = 12'b010100000000;
		14'b11010110010110: color_data = 12'b010100000000;
		14'b11010110010111: color_data = 12'b010100000000;
		14'b11010110011000: color_data = 12'b010100000000;
		14'b11010110011001: color_data = 12'b010100000000;
		14'b11010110011010: color_data = 12'b010100000000;
		14'b11010110011011: color_data = 12'b010100000000;
		14'b11010110011100: color_data = 12'b010100000000;
		14'b11010110011101: color_data = 12'b010100000000;
		14'b11010110011110: color_data = 12'b010100000000;
		14'b11010110011111: color_data = 12'b010100000000;
		14'b11010110100000: color_data = 12'b010100000000;
		14'b11010111000101: color_data = 12'b010100000000;
		14'b11010111000110: color_data = 12'b010100000000;
		14'b11010111000111: color_data = 12'b010100000000;
		14'b11010111001111: color_data = 12'b010100000000;
		14'b11010111010000: color_data = 12'b101000000000;
		14'b11010111010001: color_data = 12'b101000000000;
		14'b11010111010010: color_data = 12'b101000000000;
		14'b11010111010011: color_data = 12'b101000000000;
		14'b11010111010100: color_data = 12'b101000000000;
		14'b11010111010101: color_data = 12'b101000000000;
		14'b11010111010110: color_data = 12'b010100000000;
		14'b11010111010111: color_data = 12'b010100000000;
		14'b11010111011000: color_data = 12'b010100000000;
		14'b11010111011001: color_data = 12'b010100000000;
		14'b11010111011010: color_data = 12'b010100000000;
		14'b11010111011011: color_data = 12'b101000000000;
		14'b11010111011100: color_data = 12'b010100000000;
		14'b11010111011101: color_data = 12'b010100000000;
		14'b11010111011110: color_data = 12'b010100000000;
		14'b11010111011111: color_data = 12'b010100000000;
		14'b11011000001111: color_data = 12'b010100000000;
		14'b11011000010000: color_data = 12'b010100000000;
		14'b11011000010001: color_data = 12'b010100000000;
		14'b11011000010010: color_data = 12'b010100000000;
		14'b11011000010011: color_data = 12'b010100000000;
		14'b11011000010100: color_data = 12'b010100000000;
		14'b11011000010101: color_data = 12'b010100000000;
		14'b11011000010110: color_data = 12'b010100000000;
		14'b11011000110100: color_data = 12'b010100000000;
		14'b11011000110101: color_data = 12'b010100000000;
		14'b11011001000110: color_data = 12'b010100000000;
		14'b11011001000111: color_data = 12'b101000000000;
		14'b11011001001000: color_data = 12'b101000000000;
		14'b11011001001001: color_data = 12'b101000000000;
		14'b11011001001010: color_data = 12'b101000000000;
		14'b11011001001011: color_data = 12'b101000000000;
		14'b11011001001100: color_data = 12'b101000000000;
		14'b11011001001101: color_data = 12'b101000000000;
		14'b11011001001110: color_data = 12'b101000000000;
		14'b11011001001111: color_data = 12'b101000000000;
		14'b11011001010000: color_data = 12'b101000000000;
		14'b11011001010001: color_data = 12'b101000000000;
		14'b11011001010010: color_data = 12'b101000000000;
		14'b11011001010011: color_data = 12'b101000000000;
		14'b11011001010100: color_data = 12'b101000000000;
		14'b11011001010101: color_data = 12'b101000000000;
		14'b11011001010110: color_data = 12'b010100000000;
		14'b11011001010111: color_data = 12'b010100000000;
		14'b11011001011000: color_data = 12'b010100000000;
		14'b11011001011001: color_data = 12'b010100000000;
		14'b11011001011010: color_data = 12'b010100000000;
		14'b11011001011011: color_data = 12'b010100000000;
		14'b11011010110110: color_data = 12'b010100000000;
		14'b11011011001000: color_data = 12'b010100000000;
		14'b11011011001001: color_data = 12'b010100000000;
		14'b11011011001010: color_data = 12'b010100000000;
		14'b11011011001011: color_data = 12'b010100000000;
		14'b11011011001100: color_data = 12'b101000000000;
		14'b11011011001101: color_data = 12'b101000000000;
		14'b11011011001110: color_data = 12'b101000000000;
		14'b11011011001111: color_data = 12'b101000000000;
		14'b11011011010000: color_data = 12'b101000000000;
		14'b11011011010001: color_data = 12'b101000000000;
		14'b11011011010010: color_data = 12'b101000000000;
		14'b11011011010011: color_data = 12'b101000000000;
		14'b11011011010100: color_data = 12'b101000000000;
		14'b11011011010101: color_data = 12'b101000000000;
		14'b11011011010110: color_data = 12'b101000000000;
		14'b11011011010111: color_data = 12'b010100000000;
		14'b11011011011000: color_data = 12'b010100000000;
		default: color_data = 12'b000000000000;
	endcase
endmodule